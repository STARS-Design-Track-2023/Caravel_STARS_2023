* NGSPICE file created from synth.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

.subckt synth clk en keypad_i[0] keypad_i[10] keypad_i[11] keypad_i[12] keypad_i[13]
+ keypad_i[14] keypad_i[1] keypad_i[2] keypad_i[3] keypad_i[4] keypad_i[5] keypad_i[6]
+ keypad_i[7] keypad_i[8] keypad_i[9] n_rst pwm_o sound_series[0] sound_series[1]
+ sound_series[2] sound_series[3] vccd1 vssd1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1270_ _0583_ _0584_ _0585_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1606_ _0147_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__clkbuf_1
X_0985_ kp_encoder.sync_out\[4\] kp_encoder.sync_out\[5\] kp_encoder.sync_out\[6\]
+ kp_encoder.sync_out\[7\] vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__or4b_1
X_1468_ net114 _0632_ _0634_ seq_div.R\[21\] vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1537_ _0106_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__clkbuf_1
X_1399_ _0709_ seq_div.R\[8\] _0707_ vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1253_ clk8.count\[19\] clk8.count\[18\] _0567_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__and3_1
X_1322_ _0633_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__clkbuf_8
X_1184_ clk8.count\[3\] clk8.count\[2\] clk8.count\[4\] clk8.count\[5\] vssd1 vssd1
+ vccd1 vccd1 _0523_ sky130_fd_sc_hd__or4b_1
XFILLER_0_46_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_12_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0968_ kp_encoder.sync_out\[4\] kp_encoder.sync_out\[5\] kp_encoder.sync_out\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__or3b_1
XFILLER_0_24_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0899_ _0260_ _0272_ _0238_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0822_ _0154_ _0184_ _0196_ SS_FSM.count\[2\] vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1236_ clk8.count\[12\] clk8.count\[13\] _0553_ clk8.count\[14\] vssd1 vssd1 vccd1
+ vccd1 _0561_ sky130_fd_sc_hd__a31o_1
X_1305_ pwm.count\[5\] _0597_ _0593_ pwm.count\[6\] _0620_ vssd1 vssd1 vccd1 vccd1
+ _0621_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1167_ _0510_ _0511_ _0331_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__and3b_1
X_1098_ _0463_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1021_ _0375_ _0391_ _0382_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1785_ clknet_4_3_0_clk net55 net30 vssd1 vssd1 vccd1 vccd1 kp_encoder.last_sk sky130_fd_sc_hd__dfrtp_1
X_0805_ SS_FSM.count\[6\] SS_FSM.count\[7\] vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1219_ clk8.count\[9\] _0546_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold63 clk8.count\[13\] vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 seq_div.Q\[2\] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 clk8.count\[3\] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 SS_FSM.count\[7\] vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold30 seq_div.dividend\[0\] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold85 seq_div.dividend\[0\] vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ _0237_ _0214_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__nor2_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1004_ _0348_ _0349_ _0350_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_4_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1768_ clknet_4_10_0_clk net8 net34 vssd1 vssd1 vccd1 vccd1 kp_encoder.q\[1\] sky130_fd_sc_hd__dfrtp_1
X_1699_ clknet_4_1_0_clk _0055_ net29 vssd1 vssd1 vccd1 vccd1 SS_FSM.count\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 sound_series[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1622_ clknet_4_3_0_clk SS_FSM.next_sound\[1\] net30 vssd1 vssd1 vccd1 vccd1 SS_FSM.sound\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_1484_ _0778_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__clkbuf_1
X_1553_ _0179_ _0117_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__nand2_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0984_ kp_encoder.sync_out\[2\] kp_encoder.sync_out\[3\] vssd1 vssd1 vccd1 vccd1
+ _0355_ sky130_fd_sc_hd__nor2_1
X_1605_ net130 osc.count\[14\] _0132_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__mux2_1
X_1536_ seq_div.D\[11\] _0105_ _0631_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__mux2_1
X_1467_ _0765_ seq_div.R\[20\] _0707_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1398_ seq_div.D\[0\] _0695_ vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1252_ _0572_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[18\] sky130_fd_sc_hd__clkbuf_1
X_1321_ _0626_ _0631_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__nor2_1
X_1183_ net61 _0519_ _0522_ vssd1 vssd1 vccd1 vccd1 pwm.next_count\[7\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0967_ kp_encoder.sync_out\[10\] vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1519_ _0435_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__inv_2
X_0898_ _0232_ _0268_ _0271_ _0175_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0821_ SS_FSM.count\[3\] vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1235_ clk8.count\[13\] clk8.count\[14\] _0556_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__and3_1
X_1304_ pwm.count\[4\] _0601_ _0597_ pwm.count\[5\] _0619_ vssd1 vssd1 vccd1 vccd1
+ _0620_ sky130_fd_sc_hd__o221a_1
X_1166_ pwm.count\[0\] pwm.count\[1\] pwm.count\[2\] vssd1 vssd1 vccd1 vccd1 _0511_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1097_ _0461_ _0417_ _0448_ _0462_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__and4b_1
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1020_ _0361_ _0377_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_4_11_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1784_ clknet_4_7_0_clk net50 net31 vssd1 vssd1 vccd1 vccd1 kp_encoder.last_mk sky130_fd_sc_hd__dfrtp_1
X_0804_ SS_FSM.count\[0\] vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1218_ _0548_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_1149_ net93 _0497_ _0499_ vssd1 vssd1 vccd1 vccd1 clk_div.next_count\[4\] sky130_fd_sc_hd__o21a_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold64 clk8.next_count\[13\] vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 _0029_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 pwm.count\[0\] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 seq_div.dividend\[10\] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 _0003_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 seq_div.dividend\[1\] vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 seq_div.dividend\[4\] vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1003_ _0351_ _0361_ _0370_ _0373_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_16_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1698_ clknet_4_1_0_clk _0054_ net28 vssd1 vssd1 vccd1 vccd1 SS_FSM.count\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1767_ clknet_4_10_0_clk net2 net34 vssd1 vssd1 vccd1 vccd1 kp_encoder.q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 sound_series[2] sky130_fd_sc_hd__clkbuf_4
X_1621_ clknet_4_3_0_clk SS_FSM.next_sound\[0\] net30 vssd1 vssd1 vccd1 vccd1 SS_FSM.sound\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_1552_ _0172_ _0173_ _0269_ _0116_ _0236_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__a41o_1
XFILLER_0_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1483_ seq_div.Q\[1\] seq_div.q_out\[1\] _0776_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__mux2_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0983_ kp_encoder.sync_out\[9\] vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__inv_2
X_1604_ _0146_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__clkbuf_1
X_1535_ _0395_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__inv_2
X_1466_ _0671_ _0764_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__xnor2_1
X_1397_ net68 _0632_ _0634_ seq_div.R\[8\] _0708_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1320_ _0631_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__buf_6
X_1182_ net61 _0519_ _0331_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__o21ai_1
X_1251_ _0570_ _0531_ _0571_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__and3b_1
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0897_ _0167_ _0269_ _0270_ _0264_ _0214_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__a2111o_1
X_0966_ kp_encoder.sync_out\[8\] _0334_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1449_ _0749_ _0750_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1518_ _0094_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0820_ _0179_ _0162_ _0165_ _0183_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__or4_4
XFILLER_0_24_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1303_ pwm.count\[3\] _0605_ _0601_ pwm.count\[4\] _0618_ vssd1 vssd1 vccd1 vccd1
+ _0619_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1234_ net101 _0556_ _0559_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[13\] sky130_fd_sc_hd__o21a_1
X_1165_ pwm.count\[2\] pwm.count\[0\] pwm.count\[1\] vssd1 vssd1 vccd1 vccd1 _0510_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_35_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1096_ osc.count\[5\] _0458_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0949_ _0159_ _0314_ _0316_ _0320_ _0214_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__o311a_1
X_1783_ clknet_4_15_0_clk net7 net38 vssd1 vssd1 vccd1 vccd1 kp_encoder.q\[14\] sky130_fd_sc_hd__dfrtp_1
X_0803_ _0177_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1217_ _0546_ _0531_ _0547_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__and3b_1
X_1148_ net93 _0497_ _0350_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__a21oi_1
X_1079_ osc.count\[0\] osc.count\[1\] vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold21 seq_div.Q\[7\] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 seq_div.Q\[0\] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 seq_div.dividend\[13\] vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 clk_div.count\[3\] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 clk8.count\[4\] vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 seq_div.dividend\[11\] vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 _0013_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 kp_encoder.q\[2\] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1002_ net1 _0372_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__and2_2
XFILLER_0_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1766_ clknet_4_15_0_clk net46 net38 vssd1 vssd1 vccd1 vccd1 kp_encoder.sync_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1697_ clknet_4_1_0_clk _0053_ net29 vssd1 vssd1 vccd1 vccd1 SS_FSM.count\[2\] sky130_fd_sc_hd__dfstp_4
XFILLER_0_12_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 sound_series[3] sky130_fd_sc_hd__buf_2
X_1620_ clknet_4_13_0_clk _0002_ net37 vssd1 vssd1 vccd1 vccd1 seq_div.count_div\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1482_ _0777_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__clkbuf_1
X_1551_ _0196_ _0193_ _0222_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__or3_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1749_ clknet_4_5_0_clk clk8.next_count\[18\] net32 vssd1 vssd1 vccd1 vccd1 clk8.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0982_ net20 _0344_ _0346_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__or3_1
X_1603_ net129 osc.count\[13\] _0132_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__mux2_1
X_1465_ _0701_ _0760_ _0676_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__o21ai_2
X_1534_ _0104_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1396_ _0707_ _0628_ seq_div.D\[0\] vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__and3b_1
XFILLER_0_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1250_ clk8.count\[18\] _0567_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__or2_1
X_1181_ _0521_ vssd1 vssd1 vccd1 vccd1 pwm.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0965_ _0335_ kp_encoder.sync_out\[11\] kp_encoder.sync_out\[12\] vssd1 vssd1 vccd1
+ vccd1 _0336_ sky130_fd_sc_hd__or3b_1
X_0896_ _0154_ SS_FSM.count\[5\] vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__nor2_1
X_1448_ _0691_ _0742_ _0661_ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1517_ seq_div.D\[4\] _0093_ _0632_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__mux2_1
X_1379_ _0640_ _0659_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1233_ clk8.count\[13\] _0556_ _0531_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__a21boi_1
X_1302_ pwm.count\[2\] _0609_ _0605_ pwm.count\[3\] _0617_ vssd1 vssd1 vccd1 vccd1
+ _0618_ sky130_fd_sc_hd__o221a_1
X_1164_ net58 net71 _0509_ vssd1 vssd1 vccd1 vccd1 pwm.next_count\[1\] sky130_fd_sc_hd__a21oi_1
X_1095_ osc.count\[5\] osc.count\[4\] _0455_ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0948_ _0317_ _0318_ _0319_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0879_ SS_FSM.count\[3\] _0162_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0802_ _0157_ _0158_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1782_ clknet_4_7_0_clk net6 net31 vssd1 vssd1 vccd1 vccd1 kp_encoder.q\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1216_ clk8.count\[7\] clk8.count\[6\] _0540_ clk8.count\[8\] vssd1 vssd1 vccd1 vccd1
+ _0547_ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1147_ net70 _0494_ _0498_ vssd1 vssd1 vccd1 vccd1 clk_div.next_count\[3\] sky130_fd_sc_hd__o21a_1
X_1078_ _0331_ net97 _0417_ _0448_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[0\] sky130_fd_sc_hd__nand4_1
Xhold22 _0034_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 kp_encoder.q\[0\] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 _0028_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 pwm.count\[1\] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 clk_div.count\[4\] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 seq_div.D\[12\] vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 seq_div.dividend\[1\] vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 seq_div.D\[0\] vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1001_ _0334_ _0344_ _0346_ _0371_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__a31o_1
X_1765_ clknet_4_7_0_clk net43 net31 vssd1 vssd1 vccd1 vccd1 kp_encoder.sync_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1696_ clknet_4_0_0_clk _0052_ net28 vssd1 vssd1 vccd1 vccd1 SS_FSM.count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1481_ net120 seq_div.q_out\[0\] _0776_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__mux2_1
X_1550_ _0240_ _0114_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__nor2_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1748_ clknet_4_5_0_clk clk8.next_count\[17\] net32 vssd1 vssd1 vccd1 vccd1 clk8.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1679_ clknet_4_9_0_clk _0035_ net33 vssd1 vssd1 vccd1 vccd1 seq_div.D\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0981_ _0344_ _0346_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__nand2_2
X_1602_ _0145_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1464_ _0628_ _0762_ _0763_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1533_ net119 _0103_ _0631_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1395_ _0706_ vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__buf_6
XFILLER_0_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1180_ _0519_ _0331_ _0520_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__and3b_1
XFILLER_0_46_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0964_ kp_encoder.sync_out\[8\] kp_encoder.sync_out\[9\] kp_encoder.sync_out\[10\]
+ _0334_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__or4_1
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1516_ _0381_ _0392_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__nand2_1
X_0895_ SS_FSM.count\[3\] _0190_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__or2_2
X_1447_ _0689_ _0658_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__nor2_1
X_1378_ _0664_ _0689_ _0658_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1232_ _0558_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[12\] sky130_fd_sc_hd__clkbuf_1
X_1301_ pwm.count\[1\] _0615_ _0609_ pwm.count\[2\] _0616_ vssd1 vssd1 vccd1 vccd1
+ _0617_ sky130_fd_sc_hd__a221o_1
X_1163_ pwm.count\[0\] net71 _0331_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__o21ai_1
X_1094_ _0460_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0947_ _0167_ _0195_ _0213_ _0159_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0878_ _0228_ _0248_ _0251_ _0178_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1781_ clknet_4_5_0_clk net5 net31 vssd1 vssd1 vccd1 vccd1 kp_encoder.q\[12\] sky130_fd_sc_hd__dfrtp_1
X_0801_ _0169_ net25 vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_21_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1215_ clk8.count\[7\] clk8.count\[8\] _0543_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1146_ _0350_ _0497_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1077_ _0443_ _0445_ _0405_ _0413_ _0447_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__a2111o_4
XFILLER_0_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold12 kp_encoder.sync_out\[13\] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 pwm.count\[7\] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 pwm.next_count\[1\] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 clk_div.count\[1\] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 seq_div.dividend\[4\] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 clk8.count\[16\] vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 SS_FSM.count\[8\] vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 seq_div.dividend\[5\] vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1000_ _0327_ _0329_ _0344_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1764_ clknet_4_6_0_clk net51 net30 vssd1 vssd1 vccd1 vccd1 kp_encoder.sync_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1695_ clknet_4_0_0_clk _0051_ net28 vssd1 vssd1 vccd1 vccd1 SS_FSM.count\[0\] sky130_fd_sc_hd__dfrtp_4
X_1129_ _0485_ _0417_ _0448_ _0486_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__and4b_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1480_ seq_div.state\[1\] seq_div.state\[0\] vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__nand2_4
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1678_ clknet_4_13_0_clk net60 net37 vssd1 vssd1 vccd1 vccd1 seq_div.Q\[7\] sky130_fd_sc_hd__dfrtp_1
X_1747_ clknet_4_5_0_clk clk8.next_count\[16\] net32 vssd1 vssd1 vccd1 vccd1 clk8.count\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0980_ _0348_ _0349_ _0350_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__a21o_1
X_1601_ seq_div.dividend\[12\] osc.count\[12\] _0132_ vssd1 vssd1 vccd1 vccd1 _0145_
+ sky130_fd_sc_hd__mux2_1
X_1532_ _0411_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1463_ seq_div.dividend\[12\] _0632_ _0634_ seq_div.R\[20\] vssd1 vssd1 vccd1 vccd1
+ _0763_ sky130_fd_sc_hd__a22o_1
X_1394_ _0705_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0894_ _0178_ _0265_ _0267_ _0176_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__a211o_1
X_0963_ _0332_ _0333_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__or2_1
X_1515_ _0092_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__clkbuf_1
X_1377_ _0636_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__inv_2
X_1446_ net88 _0712_ _0717_ seq_div.R\[17\] _0748_ vssd1 vssd1 vccd1 vccd1 _0012_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1231_ _0556_ _0331_ _0557_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__and3b_1
X_1300_ pwm.count\[0\] _0592_ _0610_ _0614_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__o31a_1
X_1162_ _0350_ net58 vssd1 vssd1 vccd1 vccd1 pwm.next_count\[0\] sky130_fd_sc_hd__nor2_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1093_ _0458_ _0417_ _0448_ _0459_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__and4b_1
XFILLER_0_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0877_ _0249_ _0250_ _0228_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__o21ai_1
X_0946_ _0205_ _0288_ _0228_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1429_ _0628_ _0733_ _0734_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0800_ SS_FSM.count\[8\] _0171_ _0174_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__a21o_4
X_1780_ clknet_4_1_0_clk net4 net29 vssd1 vssd1 vccd1 vccd1 kp_encoder.q\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1214_ net106 _0543_ _0545_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[7\] sky130_fd_sc_hd__o21ba_1
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1145_ clk_div.count\[3\] _0494_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1076_ _0409_ _0446_ _0412_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__or3b_1
X_0929_ _0178_ _0300_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__or2_1
Xhold24 seq_div.Q\[5\] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold68 clk8.count\[7\] vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 seq_div.count_div\[1\] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 kp_encoder.q\[12\] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 seq_div.state\[1\] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 clk_div.next_count\[1\] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 seq_div.dividend\[11\] vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1694_ clknet_4_12_0_clk _0050_ net35 vssd1 vssd1 vccd1 vccd1 seq_div.D\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1763_ clknet_4_3_0_clk net47 net30 vssd1 vssd1 vccd1 vccd1 kp_encoder.sync_out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1128_ osc.count\[13\] _0482_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1059_ _0383_ _0378_ _0429_ _0382_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__o22ai_2
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1746_ clknet_4_5_0_clk clk8.next_count\[15\] net32 vssd1 vssd1 vccd1 vccd1 clk8.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1677_ clknet_4_13_0_clk net63 net36 vssd1 vssd1 vccd1 vccd1 seq_div.Q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1462_ _0761_ seq_div.R\[19\] _0707_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__mux2_1
X_1600_ _0144_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__clkbuf_1
X_1531_ _0102_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1393_ seq_div.R\[23\] _0681_ _0682_ _0704_ vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__and4b_1
XFILLER_0_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1729_ clknet_4_7_0_clk pwm.next_count\[6\] net31 vssd1 vssd1 vccd1 vccd1 pwm.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0962_ kp_encoder.sync_out\[4\] kp_encoder.sync_out\[5\] kp_encoder.sync_out\[6\]
+ kp_encoder.sync_out\[7\] vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__or4_1
X_0893_ _0228_ _0261_ _0253_ _0266_ _0178_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__a311oi_1
X_1445_ seq_div.R\[16\] _0707_ _0747_ _0625_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__a211o_1
X_1514_ seq_div.D\[3\] _0091_ _0632_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1376_ _0684_ _0686_ _0687_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1230_ clk8.count\[12\] _0553_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__or2_1
X_1161_ _0508_ vssd1 vssd1 vccd1 vccd1 clk_div.next_count\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1092_ osc.count\[4\] _0455_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0945_ _0189_ _0186_ _0205_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__o21a_1
X_0876_ _0154_ _0155_ _0196_ SS_FSM.count\[2\] vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__and4_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1428_ net78 _0632_ _0634_ seq_div.R\[14\] vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__a22o_1
X_1359_ _0668_ _0670_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1213_ clk8.count\[7\] clk8.count\[6\] _0540_ _0350_ vssd1 vssd1 vccd1 vccd1 _0545_
+ sky130_fd_sc_hd__a31o_1
X_1144_ _0496_ vssd1 vssd1 vccd1 vccd1 clk_div.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1075_ _0393_ _0407_ osc.count\[8\] vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0859_ _0180_ _0206_ _0178_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__or3_2
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0928_ _0185_ _0270_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__nand2_1
Xhold25 _0033_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 _0629_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 _0076_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 kp_encoder.q\[8\] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 seq_div.dividend\[2\] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 seq_div.dividend\[5\] vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1693_ clknet_4_12_0_clk _0049_ net35 vssd1 vssd1 vccd1 vccd1 seq_div.D\[14\] sky130_fd_sc_hd__dfrtp_1
X_1762_ clknet_4_2_0_clk net42 net28 vssd1 vssd1 vccd1 vccd1 kp_encoder.sync_out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1127_ osc.count\[13\] _0482_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__and2_1
X_1058_ _0361_ _0377_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1745_ clknet_4_5_0_clk clk8.next_count\[14\] net32 vssd1 vssd1 vccd1 vccd1 clk8.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1676_ clknet_4_15_0_clk _0032_ net37 vssd1 vssd1 vccd1 vccd1 seq_div.Q\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1461_ _0701_ _0760_ vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__xor2_1
X_1530_ seq_div.D\[9\] _0101_ _0631_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1392_ _0683_ _0688_ _0693_ _0703_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1728_ clknet_4_7_0_clk pwm.next_count\[5\] net31 vssd1 vssd1 vccd1 vccd1 pwm.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1659_ clknet_4_1_0_clk clk_div.next_count\[4\] net30 vssd1 vssd1 vccd1 vccd1 clk_div.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0961_ kp_encoder.sync_out\[0\] kp_encoder.sync_out\[1\] kp_encoder.sync_out\[2\]
+ kp_encoder.sync_out\[3\] vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__or4_2
XFILLER_0_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0892_ _0184_ SS_FSM.count\[2\] _0166_ _0196_ _0154_ vssd1 vssd1 vccd1 vccd1 _0266_
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1444_ _0707_ _0746_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__nor2_1
X_1513_ _0420_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__inv_2
X_1375_ _0647_ _0651_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1160_ _0331_ _0506_ _0507_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__and3_1
X_1091_ osc.count\[4\] osc.count\[3\] _0452_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0944_ _0249_ _0315_ _0228_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0875_ _0209_ _0210_ _0165_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__a21oi_2
X_1358_ _0669_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__inv_2
X_1427_ _0732_ seq_div.R\[13\] _0707_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__mux2_1
X_1289_ seq_div.q_out\[3\] _0588_ _0604_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1212_ _0543_ _0544_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[6\] sky130_fd_sc_hd__nor2_1
XFILLER_0_47_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1143_ _0494_ _0331_ _0495_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__and3b_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1074_ _0418_ _0419_ _0441_ _0444_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0927_ _0179_ _0184_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0789_ SS_FSM.count\[0\] _0155_ SS_FSM.count\[2\] SS_FSM.count\[3\] vssd1 vssd1 vccd1
+ vccd1 _0164_ sky130_fd_sc_hd__o31a_2
XFILLER_0_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0858_ _0176_ _0227_ _0231_ _0159_ _0232_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__o221a_1
Xhold37 seq_div.Q\[3\] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 clk_div.count\[0\] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 seq_div.count_div\[0\] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 osc.count\[0\] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 kp_encoder.q\[1\] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1761_ clknet_4_3_0_clk net54 net30 vssd1 vssd1 vccd1 vccd1 kp_encoder.sync_out\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1692_ clknet_4_12_0_clk _0048_ net35 vssd1 vssd1 vccd1 vccd1 seq_div.D\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1126_ _0484_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1057_ osc.count\[1\] _0427_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1744_ clknet_4_5_0_clk net102 net29 vssd1 vssd1 vccd1 vccd1 clk8.count\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1675_ clknet_4_15_0_clk _0031_ net37 vssd1 vssd1 vccd1 vccd1 seq_div.Q\[4\] sky130_fd_sc_hd__dfrtp_1
X_1109_ _0470_ _0417_ _0448_ _0471_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__and4b_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1460_ _0693_ _0741_ _0758_ _0759_ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1391_ _0696_ _0700_ _0701_ _0702_ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__or4b_1
XFILLER_0_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1727_ clknet_4_7_0_clk pwm.next_count\[4\] net31 vssd1 vssd1 vccd1 vccd1 pwm.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_1658_ clknet_4_4_0_clk clk_div.next_count\[3\] net30 vssd1 vssd1 vccd1 vccd1 clk_div.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1589_ net78 osc.count\[6\] _0132_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0960_ net1 vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__buf_4
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1512_ _0090_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0891_ _0167_ _0195_ _0263_ _0264_ _0225_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__a32o_1
X_1443_ _0691_ _0745_ vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__xor2_1
X_1374_ _0643_ _0685_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1090_ _0457_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
X_0943_ _0210_ _0262_ _0189_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__a21oi_1
X_0874_ _0165_ _0244_ _0195_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1288_ _0582_ _0602_ _0603_ _0591_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__a31o_1
X_1357_ seq_div.D\[13\] seq_div.R\[20\] vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__and2b_1
X_1426_ _0699_ _0731_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1142_ clk_div.count\[1\] clk_div.count\[0\] clk_div.count\[2\] vssd1 vssd1 vccd1
+ vccd1 _0495_ sky130_fd_sc_hd__a21o_1
X_1211_ clk8.count\[6\] _0540_ _0531_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1073_ _0438_ _0436_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__nand2_1
X_0857_ _0171_ _0216_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__nand2_2
X_0926_ _0240_ _0236_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__nor2_2
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold38 _0030_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 kp_encoder.q\[9\] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 clk8.count\[1\] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ net96 _0712_ _0716_ _0625_ _0718_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__o221a_1
X_0788_ SS_FSM.count\[0\] _0155_ SS_FSM.count\[3\] SS_FSM.count\[2\] vssd1 vssd1 vccd1
+ vccd1 _0163_ sky130_fd_sc_hd__nor4_4
Xhold49 seq_div.D\[6\] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1691_ clknet_4_14_0_clk _0047_ net37 vssd1 vssd1 vccd1 vccd1 seq_div.D\[12\] sky130_fd_sc_hd__dfrtp_1
X_1760_ clknet_4_3_0_clk net52 net30 vssd1 vssd1 vccd1 vccd1 kp_encoder.sync_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1125_ _0482_ _0417_ _0448_ _0483_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__and4b_1
XFILLER_0_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1056_ _0375_ _0425_ _0426_ _0420_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__a31o_1
X_0909_ _0178_ _0279_ _0281_ _0214_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1743_ clknet_4_7_0_clk clk8.next_count\[12\] net31 vssd1 vssd1 vccd1 vccd1 clk8.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1674_ clknet_4_13_0_clk net76 net37 vssd1 vssd1 vccd1 vccd1 seq_div.Q\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1039_ _0375_ _0361_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__nand2_1
X_1108_ osc.count\[8\] _0467_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1390_ seq_div.D\[15\] seq_div.R\[22\] vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1726_ clknet_4_7_0_clk pwm.next_count\[3\] net31 vssd1 vssd1 vccd1 vccd1 pwm.count\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_1657_ clknet_4_4_0_clk clk_div.next_count\[2\] net30 vssd1 vssd1 vccd1 vccd1 clk_div.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1588_ _0138_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__clkbuf_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0890_ _0166_ _0249_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1442_ _0660_ _0742_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__nand2_1
X_1511_ seq_div.D\[2\] _0089_ _0632_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1373_ _0645_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1709_ clknet_4_9_0_clk _0065_ net33 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout30 net32 vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_6
XFILLER_0_36_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0942_ _0228_ _0248_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__nor2_1
X_0873_ _0241_ _0243_ _0245_ _0246_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1425_ _0654_ _0727_ _0650_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__a21o_1
X_1287_ _0585_ seq_div.q_out\[2\] vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__nand2_1
X_1356_ seq_div.R\[20\] seq_div.D\[13\] vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__or2b_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1210_ clk8.count\[6\] _0540_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__and2_1
X_1141_ clk_div.count\[1\] clk_div.count\[0\] clk_div.count\[2\] vssd1 vssd1 vccd1
+ vccd1 _0494_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1072_ _0418_ _0419_ _0424_ _0433_ _0442_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0925_ _0175_ _0296_ _0297_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0787_ _0160_ _0161_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__and2_2
X_0856_ _0169_ _0165_ _0228_ _0229_ _0230_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__o41a_1
Xhold39 seq_div.Q\[4\] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 kp_encoder.sync_out\[14\] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold28 clk8.next_count\[1\] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ seq_div.R\[10\] _0717_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__or2_1
X_1339_ seq_div.D\[4\] seq_div.R\[11\] vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__or2b_1
XFILLER_0_21_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1690_ clknet_4_12_0_clk _0046_ net37 vssd1 vssd1 vccd1 vccd1 seq_div.D\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1124_ osc.count\[12\] _0479_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__or2_1
X_1055_ _0361_ _0370_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput18 net18 vssd1 vssd1 vccd1 vccd1 pwm_o sky130_fd_sc_hd__clkbuf_4
X_0839_ SS_FSM.count\[6\] net24 vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__xnor2_4
X_0908_ _0167_ _0187_ _0192_ _0280_ _0159_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__a311o_1
XFILLER_0_11_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1673_ clknet_4_13_0_clk net80 net36 vssd1 vssd1 vccd1 vccd1 seq_div.Q\[2\] sky130_fd_sc_hd__dfrtp_1
X_1742_ clknet_4_7_0_clk clk8.next_count\[11\] net31 vssd1 vssd1 vccd1 vccd1 clk8.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1038_ osc.count\[8\] _0393_ _0407_ _0408_ osc.count\[9\] vssd1 vssd1 vccd1 vccd1
+ _0409_ sky130_fd_sc_hd__a32o_1
X_1107_ osc.count\[8\] _0467_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1725_ clknet_4_7_0_clk pwm.next_count\[2\] net31 vssd1 vssd1 vccd1 vccd1 pwm.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1656_ clknet_4_6_0_clk net95 net30 vssd1 vssd1 vccd1 vccd1 clk_div.count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1587_ net127 osc.count\[5\] _0132_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1510_ _0422_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__inv_2
X_1441_ net99 _0712_ _0717_ seq_div.R\[16\] _0744_ vssd1 vssd1 vccd1 vccd1 _0011_
+ sky130_fd_sc_hd__o221a_1
X_1372_ _0644_ _0648_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__or2b_1
X_1708_ clknet_4_9_0_clk _0064_ net33 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1639_ clknet_4_3_0_clk osc.next_count\[0\] net30 vssd1 vssd1 vccd1 vccd1 osc.count\[0\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout31 net32 vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_4
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0941_ _0310_ _0312_ _0175_ _0232_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__a211o_1
X_0872_ _0167_ _0195_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__nor2_1
X_1355_ _0635_ _0665_ _0666_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__and3_1
X_1424_ _0628_ _0729_ _0730_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__a21o_1
X_1286_ _0585_ seq_div.q_out\[2\] vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1140_ net94 net64 _0493_ vssd1 vssd1 vccd1 vccd1 clk_div.next_count\[1\] sky130_fd_sc_hd__o21a_1
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1071_ _0434_ _0436_ _0438_ _0441_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__or4bb_1
X_0924_ SS_FSM.count\[3\] SS_FSM.count\[2\] _0234_ _0175_ vssd1 vssd1 vccd1 vccd1
+ _0297_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_11_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0786_ SS_FSM.count\[0\] _0155_ SS_FSM.count\[2\] vssd1 vssd1 vccd1 vccd1 _0161_
+ sky130_fd_sc_hd__o21ai_2
X_0855_ _0209_ _0210_ _0167_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__a21o_1
Xhold29 pwm.count\[7\] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 clk8.count\[20\] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1407_ _0625_ _0712_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__nand2_2
X_1338_ seq_div.D\[5\] seq_div.R\[12\] vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__and2b_1
X_1269_ seq_div.q_out\[7\] vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1123_ osc.count\[12\] osc.count\[11\] _0476_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__and3_1
X_1054_ _0361_ _0370_ _0382_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__o21ai_1
X_0907_ _0189_ _0229_ _0228_ _0209_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__o211a_1
Xoutput19 net19 vssd1 vssd1 vccd1 vccd1 sound_series[0] sky130_fd_sc_hd__clkbuf_4
X_0838_ _0166_ _0212_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__or2_1
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1741_ clknet_4_5_0_clk clk8.next_count\[10\] net29 vssd1 vssd1 vccd1 vccd1 clk8.count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_1672_ clknet_4_13_0_clk net82 net36 vssd1 vssd1 vccd1 vccd1 seq_div.Q\[1\] sky130_fd_sc_hd__dfrtp_1
X_1106_ _0469_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1037_ _0374_ _0394_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1724_ clknet_4_6_0_clk net72 net31 vssd1 vssd1 vccd1 vccd1 pwm.count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1655_ clknet_4_7_0_clk clk_div.next_count\[0\] net30 vssd1 vssd1 vccd1 vccd1 clk_div.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1586_ _0137_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__clkbuf_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1371_ _0650_ _0654_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__or2b_1
X_1440_ seq_div.R\[15\] _0707_ _0742_ _0743_ _0625_ vssd1 vssd1 vccd1 vccd1 _0744_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1638_ clknet_4_12_0_clk _0018_ net37 vssd1 vssd1 vccd1 vccd1 seq_div.R\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1707_ clknet_4_8_0_clk _0063_ net33 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1569_ SS_FSM.count\[5\] _0123_ _0127_ _0128_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__o22a_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout32 net17 vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_4
XFILLER_0_44_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0940_ _0201_ _0257_ _0311_ _0187_ _0176_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0871_ _0205_ _0165_ _0159_ _0244_ _0214_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__a41o_1
XFILLER_0_23_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1285_ seq_div.q_out\[4\] _0588_ _0600_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__o21ai_1
X_1354_ seq_div.R\[19\] seq_div.D\[12\] vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__or2b_1
X_1423_ net107 _0632_ _0634_ seq_div.R\[13\] vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1070_ _0418_ _0419_ _0440_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0923_ _0282_ _0287_ _0295_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0854_ _0179_ _0162_ _0183_ _0190_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__o31a_1
XFILLER_0_11_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0785_ SS_FSM.count\[0\] _0155_ SS_FSM.count\[2\] vssd1 vssd1 vccd1 vccd1 _0160_
+ sky130_fd_sc_hd__or3_2
XFILLER_0_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1268_ mode_FSM.mode\[1\] seq_div.q_out\[6\] mode_FSM.mode\[0\] vssd1 vssd1 vccd1
+ vccd1 _0584_ sky130_fd_sc_hd__o21a_1
Xhold19 seq_div.count_div\[2\] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__dlygate4sd3_1
X_1406_ _0715_ seq_div.R\[9\] _0707_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__mux2_1
X_1337_ _0646_ _0647_ _0648_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1199_ _0534_ _0331_ _0535_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__and3b_1
XFILLER_0_46_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1122_ _0481_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
X_1053_ osc.count\[3\] _0420_ _0423_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0837_ _0196_ _0160_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0906_ _0167_ _0276_ _0277_ _0278_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1740_ clknet_4_4_0_clk clk8.next_count\[9\] net29 vssd1 vssd1 vccd1 vccd1 clk8.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1671_ clknet_4_13_0_clk _0027_ net35 vssd1 vssd1 vccd1 vccd1 seq_div.Q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1105_ _0467_ _0417_ _0448_ _0468_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__and4b_1
X_1036_ _0379_ _0406_ _0382_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1723_ clknet_4_6_0_clk pwm.next_count\[0\] net36 vssd1 vssd1 vccd1 vccd1 pwm.count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_1654_ clknet_4_6_0_clk osc.next_count\[15\] net35 vssd1 vssd1 vccd1 vccd1 osc.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1585_ net124 osc.count\[4\] _0132_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1019_ _0375_ _0370_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1370_ _0678_ seq_div.R\[22\] vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1637_ clknet_4_15_0_clk _0017_ net37 vssd1 vssd1 vccd1 vccd1 seq_div.R\[22\] sky130_fd_sc_hd__dfrtp_2
X_1706_ clknet_4_8_0_clk _0062_ net33 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1499_ seq_div.Q\[1\] _0628_ _0634_ net79 vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__a22o_1
X_1568_ _0237_ _0159_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__nor2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout33 net38 vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_6
XFILLER_0_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0870_ _0219_ _0222_ _0223_ _0185_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__a31o_1
X_1422_ _0728_ seq_div.R\[12\] _0707_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__mux2_1
X_1284_ _0582_ _0598_ _0599_ _0591_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__a31o_1
X_1353_ _0636_ _0662_ _0664_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0999_ _0352_ _0362_ _0369_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0922_ _0176_ _0290_ _0291_ _0294_ _0217_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__o311a_1
X_0853_ _0205_ net26 vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__xnor2_4
X_0784_ _0157_ _0158_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__nor2_8
X_1405_ _0686_ _0714_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1267_ seq_div.q_out\[6\] _0582_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__nand2_1
Xinput1 en vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_4
X_1198_ clk8.count\[1\] clk8.count\[0\] clk8.count\[2\] vssd1 vssd1 vccd1 vccd1 _0535_
+ sky130_fd_sc_hd__a21o_1
X_1336_ seq_div.R\[10\] seq_div.D\[3\] vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__or2b_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1121_ _0479_ _0417_ _0448_ _0480_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__and4b_1
X_1052_ osc.count\[3\] _0420_ _0422_ osc.count\[2\] vssd1 vssd1 vccd1 vccd1 _0423_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0836_ SS_FSM.count\[4\] net27 _0164_ _0210_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__or4_2
X_0905_ SS_FSM.count\[4\] _0156_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__nor2_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1319_ _0630_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1670_ clknet_4_13_0_clk _0026_ net36 vssd1 vssd1 vccd1 vccd1 seq_div.q_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1104_ osc.count\[7\] _0464_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__or2_1
X_1035_ _0351_ _0361_ _0377_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__nand3_2
XFILLER_0_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0819_ _0154_ SS_FSM.count\[3\] _0193_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1722_ clknet_4_13_0_clk pwm.pwm net36 vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__dfrtp_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1653_ clknet_4_6_0_clk osc.next_count\[14\] net35 vssd1 vssd1 vccd1 vccd1 osc.count\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1584_ _0136_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__clkbuf_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1018_ osc.count\[12\] _0385_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1705_ clknet_4_8_0_clk _0061_ net33 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1636_ clknet_4_15_0_clk _0016_ net37 vssd1 vssd1 vccd1 vccd1 seq_div.R\[21\] sky130_fd_sc_hd__dfrtp_1
X_1567_ SS_FSM.count\[4\] _0123_ _0126_ _0127_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__o22a_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1498_ net81 _0628_ _0634_ seq_div.Q\[1\] vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__a22o_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout34 net38 vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_6
XFILLER_0_32_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1421_ _0683_ _0727_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__xnor2_1
X_1283_ _0585_ seq_div.q_out\[3\] vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__nand2_1
X_1352_ _0635_ _0663_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0998_ _0344_ _0346_ _0368_ _0350_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__a31o_1
X_1619_ clknet_4_15_0_clk _0001_ net37 vssd1 vssd1 vccd1 vccd1 seq_div.count_div\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0921_ _0178_ _0207_ _0245_ _0293_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__a211o_1
X_0783_ SS_FSM.count\[4\] _0156_ SS_FSM.count\[5\] vssd1 vssd1 vccd1 vccd1 _0158_
+ sky130_fd_sc_hd__o21a_2
X_0852_ _0167_ _0226_ _0211_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1404_ _0713_ _0694_ _0642_ vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1335_ seq_div.R\[11\] seq_div.D\[4\] vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__or2b_1
X_1266_ _0581_ mode_FSM.mode\[0\] vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__and2_2
X_1197_ clk8.count\[1\] clk8.count\[0\] clk8.count\[2\] vssd1 vssd1 vccd1 vccd1 _0534_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_36_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 keypad_i[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1120_ osc.count\[11\] _0476_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__or2_1
X_1051_ _0375_ _0391_ _0421_ _0377_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_22_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0904_ _0206_ _0191_ _0156_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0835_ _0179_ _0155_ _0193_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__or3_2
X_1318_ _0623_ seq_div.state\[0\] vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1249_ clk8.count\[18\] _0567_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__and2_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1034_ _0388_ _0389_ _0396_ _0404_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__or4b_2
X_1103_ osc.count\[7\] osc.count\[6\] _0461_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0818_ SS_FSM.count\[2\] vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1721_ clknet_4_12_0_clk _0077_ net37 vssd1 vssd1 vccd1 vccd1 seq_div.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1652_ clknet_4_3_0_clk osc.next_count\[13\] net35 vssd1 vssd1 vccd1 vccd1 osc.count\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1583_ seq_div.dividend\[3\] osc.count\[3\] _0132_ vssd1 vssd1 vccd1 vccd1 _0136_
+ sky130_fd_sc_hd__mux2_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1017_ osc.count\[12\] _0385_ _0387_ osc.count\[13\] vssd1 vssd1 vccd1 vccd1 _0388_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1704_ clknet_4_8_0_clk _0060_ net33 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1497_ _0625_ _0707_ _0634_ net81 vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__a2bb2o_1
X_1635_ clknet_4_14_0_clk _0015_ net37 vssd1 vssd1 vccd1 vccd1 seq_div.R\[20\] sky130_fd_sc_hd__dfrtp_1
X_1566_ _0174_ _0299_ _0115_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__a21o_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout35 net38 vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_6
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1351_ seq_div.D\[11\] seq_div.R\[18\] vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__or2b_1
X_1420_ _0687_ _0723_ _0651_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__o21ai_1
X_1282_ _0585_ seq_div.q_out\[3\] vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1618_ clknet_4_15_0_clk _0000_ net37 vssd1 vssd1 vccd1 vccd1 seq_div.count_div\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0997_ kp_encoder.sync_out\[9\] _0337_ _0343_ _0367_ vssd1 vssd1 vccd1 vccd1 _0368_
+ sky130_fd_sc_hd__a211o_1
X_1549_ _0350_ _0529_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0920_ _0195_ _0292_ _0167_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__a21oi_1
X_0782_ SS_FSM.count\[4\] SS_FSM.count\[5\] _0156_ vssd1 vssd1 vccd1 vccd1 _0157_
+ sky130_fd_sc_hd__nor3_4
XFILLER_0_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0851_ _0179_ _0221_ _0225_ _0159_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__o22a_1
X_1265_ mode_FSM.mode\[1\] vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__inv_2
X_1334_ _0642_ _0643_ _0644_ _0645_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__a211o_1
X_1403_ seq_div.D\[0\] vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__inv_2
X_1196_ net65 clk8.count\[0\] _0533_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[1\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput3 keypad_i[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1050_ _0375_ _0361_ _0382_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0903_ _0179_ _0165_ _0186_ _0275_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__o31a_1
X_0834_ _0156_ _0180_ _0181_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__or3_2
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1248_ _0569_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[17\] sky130_fd_sc_hd__clkbuf_1
X_1317_ net57 _0627_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1179_ pwm.count\[6\] _0516_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__or2_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1102_ _0466_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
X_1033_ _0399_ _0400_ _0401_ _0403_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__and4b_1
XFILLER_0_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0817_ _0189_ _0191_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1720_ clknet_4_13_0_clk net74 net38 vssd1 vssd1 vccd1 vccd1 seq_div.state\[0\] sky130_fd_sc_hd__dfrtp_4
X_1651_ clknet_4_3_0_clk osc.next_count\[12\] net35 vssd1 vssd1 vccd1 vccd1 osc.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1582_ _0135_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1016_ _0375_ _0379_ _0386_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1703_ clknet_4_1_0_clk _0059_ net29 vssd1 vssd1 vccd1 vccd1 SS_FSM.count\[8\] sky130_fd_sc_hd__dfstp_1
X_1634_ clknet_4_14_0_clk _0014_ net37 vssd1 vssd1 vccd1 vccd1 seq_div.R\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1496_ _0085_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1565_ _0237_ _0167_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__nor2_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout36 net38 vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_4
XFILLER_0_32_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1281_ seq_div.q_out\[5\] _0588_ _0596_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__o21ai_1
X_1350_ _0641_ _0657_ _0658_ _0661_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0996_ _0332_ _0356_ _0366_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__o21ai_1
X_1617_ _0153_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1479_ _0628_ _0774_ net109 vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__a21o_1
X_1548_ _0113_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0850_ _0189_ _0224_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__or2_1
X_1402_ _0623_ seq_div.state\[0\] vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__nand2_4
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0781_ SS_FSM.count\[0\] _0155_ SS_FSM.count\[3\] SS_FSM.count\[2\] vssd1 vssd1 vccd1
+ vccd1 _0156_ sky130_fd_sc_hd__or4_4
XFILLER_0_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1264_ _0274_ _0577_ _0578_ SS_FSM.sound\[1\] vssd1 vssd1 vccd1 vccd1 SS_FSM.next_sound\[1\]
+ sky130_fd_sc_hd__a22o_1
Xinput4 keypad_i[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_1333_ seq_div.D\[2\] seq_div.R\[9\] vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__and2b_1
X_1195_ net65 clk8.count\[0\] _0331_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0979_ net1 vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__clkinv_8
XFILLER_0_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0833_ _0178_ _0207_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__nor2_1
X_0902_ _0179_ _0184_ SS_FSM.count\[3\] vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1247_ _0567_ _0531_ _0568_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__and3b_1
X_1178_ pwm.count\[6\] _0516_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__and2_1
X_1316_ _0627_ net85 vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1032_ osc.count\[14\] _0402_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1101_ _0464_ _0417_ _0448_ _0465_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__and4b_1
XFILLER_0_56_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0816_ _0162_ _0183_ _0190_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1650_ clknet_4_3_0_clk osc.next_count\[11\] net30 vssd1 vssd1 vccd1 vccd1 osc.count\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_1581_ net128 osc.count\[2\] _0132_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__mux2_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1015_ _0373_ _0361_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__nand2_2
XFILLER_0_60_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1779_ clknet_4_0_0_clk net3 net28 vssd1 vssd1 vccd1 vccd1 kp_encoder.q\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1702_ clknet_4_4_0_clk _0058_ net29 vssd1 vssd1 vccd1 vccd1 SS_FSM.count\[7\] sky130_fd_sc_hd__dfrtp_1
X_1633_ clknet_4_14_0_clk net92 net37 vssd1 vssd1 vccd1 vccd1 seq_div.R\[18\] sky130_fd_sc_hd__dfrtp_1
X_1564_ SS_FSM.count\[3\] _0115_ _0119_ _0125_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__a22o_1
X_1495_ net59 _0585_ _0776_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout37 net38 vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1280_ _0582_ _0594_ _0595_ _0591_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0995_ kp_encoder.sync_out\[4\] _0363_ _0332_ _0365_ kp_encoder.sync_out\[0\] vssd1
+ vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__o32a_1
X_1616_ mode_FSM.mode\[0\] _0581_ _0151_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__mux2_1
X_1547_ seq_div.D\[15\] _0112_ _0631_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__mux2_1
X_1478_ seq_div.dividend\[15\] _0632_ _0633_ net108 vssd1 vssd1 vccd1 vccd1 _0775_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0780_ SS_FSM.count\[1\] vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__buf_4
X_1401_ _0628_ _0710_ _0711_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__a21o_1
Xinput5 keypad_i[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_1194_ _0532_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[0\] sky130_fd_sc_hd__clkbuf_1
X_1263_ _0580_ vssd1 vssd1 vccd1 vccd1 SS_FSM.next_sound\[0\] sky130_fd_sc_hd__clkbuf_1
X_1332_ seq_div.D\[3\] seq_div.R\[10\] vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__and2b_1
XFILLER_0_52_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0978_ net21 _0344_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0901_ _0240_ SS_FSM.sound\[1\] vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__nor2_1
X_0832_ _0206_ _0191_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__nor2_1
X_1315_ seq_div.count_div\[0\] _0628_ net84 vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1246_ clk8.count\[15\] clk8.count\[16\] _0560_ clk8.count\[17\] vssd1 vssd1 vccd1
+ vccd1 _0568_ sky130_fd_sc_hd__a31o_1
X_1177_ _0518_ vssd1 vssd1 vccd1 vccd1 pwm.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap23 _0120_ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_9_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1100_ osc.count\[6\] _0461_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__or2_1
X_1031_ _0375_ _0386_ _0381_ _0383_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_33_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0815_ _0154_ _0155_ SS_FSM.count\[2\] vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__or3_2
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1229_ clk8.count\[12\] _0553_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1580_ _0134_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1014_ _0374_ _0376_ _0384_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1778_ clknet_4_15_0_clk net16 net38 vssd1 vssd1 vccd1 vccd1 kp_encoder.q\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1701_ clknet_4_1_0_clk _0057_ net30 vssd1 vssd1 vccd1 vccd1 SS_FSM.count\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1494_ _0084_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1632_ clknet_4_14_0_clk net89 net34 vssd1 vssd1 vccd1 vccd1 seq_div.R\[17\] sky130_fd_sc_hd__dfrtp_1
X_1563_ _0165_ _0117_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__nand2_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout38 net17 vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_6
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0994_ _0364_ kp_encoder.sync_out\[3\] kp_encoder.sync_out\[1\] vssd1 vssd1 vccd1
+ vccd1 _0365_ sky130_fd_sc_hd__a21oi_1
X_1615_ _0152_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1477_ _0773_ seq_div.R\[22\] _0707_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__mux2_1
X_1546_ _0382_ _0397_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1400_ net113 _0632_ _0634_ seq_div.R\[9\] vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__a22o_1
X_1331_ seq_div.R\[9\] seq_div.D\[2\] vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__or2b_1
Xinput6 keypad_i[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
X_1193_ clk8.count\[0\] _0531_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__and2b_1
X_1262_ _0578_ _0579_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__and2_1
X_0977_ _0336_ _0344_ _0346_ _0347_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__nand4_2
XFILLER_0_6_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1529_ _0408_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0900_ _0155_ _0159_ _0168_ _0273_ _0240_ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__a311o_2
X_0831_ _0205_ _0165_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__nand2_2
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1314_ _0626_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1245_ clk8.count\[16\] clk8.count\[17\] _0563_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__and3_1
X_1176_ _0516_ _0331_ _0517_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__and3b_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap24 net25 vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1030_ osc.count\[13\] _0387_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0814_ _0188_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1228_ _0555_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1159_ clk_div.count\[7\] _0503_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1013_ _0378_ _0379_ _0381_ _0383_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_60_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1777_ clknet_4_14_0_clk net15 net37 vssd1 vssd1 vccd1 vccd1 kp_encoder.q\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1700_ clknet_4_1_0_clk _0056_ net29 vssd1 vssd1 vccd1 vccd1 SS_FSM.count\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1631_ clknet_4_11_0_clk net100 net34 vssd1 vssd1 vccd1 vccd1 seq_div.R\[16\] sky130_fd_sc_hd__dfrtp_1
X_1493_ seq_div.Q\[6\] seq_div.q_out\[6\] _0776_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__mux2_1
X_1562_ _0124_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__clkbuf_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout28 net17 vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_6
XFILLER_0_4_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0993_ kp_encoder.sync_out\[2\] vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__inv_2
X_1614_ mode_FSM.mode\[1\] mode_FSM.mode\[0\] _0151_ vssd1 vssd1 vccd1 vccd1 _0152_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1545_ _0111_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__clkbuf_1
X_1476_ _0702_ _0772_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1261_ SS_FSM.sound\[0\] _0577_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__or2_1
X_1330_ seq_div.D\[1\] seq_div.R\[8\] vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__and2b_1
Xinput7 keypad_i[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
X_1192_ _0530_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__buf_2
XFILLER_0_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0976_ _0332_ _0333_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1459_ _0664_ _0689_ _0658_ _0661_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__or4b_1
X_1528_ _0100_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0830_ SS_FSM.count\[4\] vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1244_ net105 _0563_ _0566_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[16\] sky130_fd_sc_hd__o21ba_1
X_1313_ seq_div.count_div\[0\] seq_div.count_div\[1\] _0626_ vssd1 vssd1 vccd1 vccd1
+ _0627_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1175_ pwm.count\[4\] pwm.count\[3\] _0510_ pwm.count\[5\] vssd1 vssd1 vccd1 vccd1
+ _0517_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0959_ _0330_ vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
Xmax_cap25 _0157_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput10 keypad_i[3] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_1
X_0813_ _0163_ _0164_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1227_ _0553_ _0331_ _0554_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__and3b_1
X_1158_ clk_div.count\[7\] _0503_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__or2_1
X_1089_ _0455_ _0417_ _0448_ _0456_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__and4b_1
XFILLER_0_15_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1012_ _0382_ _0375_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__nand2_2
XFILLER_0_60_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1776_ clknet_4_2_0_clk net14 net17 vssd1 vssd1 vccd1 vccd1 kp_encoder.q\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1630_ clknet_4_11_0_clk _0010_ net34 vssd1 vssd1 vccd1 vccd1 seq_div.R\[15\] sky130_fd_sc_hd__dfrtp_1
X_1492_ _0083_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1561_ SS_FSM.count\[2\] _0121_ _0123_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__mux2_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout29 net32 vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_6
X_1759_ clknet_4_2_0_clk net44 net28 vssd1 vssd1 vccd1 vccd1 kp_encoder.sync_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0992_ kp_encoder.sync_out\[5\] vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__inv_2
X_1613_ kp_encoder.last_mk kp_encoder.sync_out\[13\] vssd1 vssd1 vccd1 vccd1 _0151_
+ sky130_fd_sc_hd__and2b_1
X_1544_ seq_div.D\[14\] _0402_ _0631_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_1475_ _0672_ _0768_ _0679_ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1191_ _0331_ _0529_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__and2_1
X_1260_ SS_FSM.sound\[0\] _0577_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__nand2_1
Xinput8 keypad_i[1] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0975_ SS_FSM.sound\[1\] _0298_ _0345_ SS_FSM.sound\[0\] vssd1 vssd1 vccd1 vccd1
+ _0346_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1527_ seq_div.D\[8\] _0099_ _0632_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__mux2_1
X_1389_ _0666_ _0676_ vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__nand2_1
X_1458_ _0635_ _0658_ _0663_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1243_ clk8.count\[15\] clk8.count\[16\] _0560_ _0350_ vssd1 vssd1 vccd1 vccd1 _0566_
+ sky130_fd_sc_hd__a31o_1
X_1174_ pwm.count\[5\] pwm.count\[4\] _0513_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1312_ _0623_ seq_div.state\[0\] vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0958_ _0327_ _0329_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0889_ _0219_ _0261_ _0262_ _0210_ _0189_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap26 net27 vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput11 keypad_i[4] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0812_ _0179_ _0165_ _0186_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1226_ clk8.count\[9\] clk8.count\[10\] _0546_ clk8.count\[11\] vssd1 vssd1 vccd1
+ vccd1 _0554_ sky130_fd_sc_hd__a31o_1
X_1157_ _0505_ vssd1 vssd1 vccd1 vccd1 clk_div.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
X_1088_ osc.count\[3\] _0452_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1011_ net1 _0372_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__nand2_4
XFILLER_0_56_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1775_ clknet_4_2_0_clk net13 net28 vssd1 vssd1 vccd1 vccd1 kp_encoder.q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1209_ _0542_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1560_ _0122_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1491_ net62 seq_div.q_out\[5\] _0776_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__mux2_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1689_ clknet_4_14_0_clk _0045_ net38 vssd1 vssd1 vccd1 vccd1 seq_div.D\[10\] sky130_fd_sc_hd__dfrtp_1
X_1758_ clknet_4_2_0_clk net45 net28 vssd1 vssd1 vccd1 vccd1 kp_encoder.sync_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0991_ net19 _0344_ _0346_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__or3_2
X_1474_ _0628_ _0770_ _0771_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__a21o_1
X_1612_ _0623_ _0132_ _0634_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__o21ai_1
X_1543_ _0110_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1190_ clk8.count\[1\] clk8.count\[0\] _0523_ _0528_ vssd1 vssd1 vccd1 vccd1 _0529_
+ sky130_fd_sc_hd__or4b_1
Xinput9 keypad_i[2] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0974_ _0297_ _0313_ _0326_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__nand3_1
XFILLER_0_6_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1457_ _0628_ _0756_ _0757_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__a21o_1
X_1526_ _0393_ _0407_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__nand2_1
X_1388_ _0697_ _0655_ _0699_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1311_ net86 _0625_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__xnor2_1
X_1242_ _0565_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[15\] sky130_fd_sc_hd__clkbuf_1
X_1173_ pwm.count\[4\] _0513_ _0515_ vssd1 vssd1 vccd1 vccd1 pwm.next_count\[4\] sky130_fd_sc_hd__o21ba_1
X_0957_ _0206_ _0328_ _0299_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0888_ _0162_ _0183_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1509_ _0088_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__clkbuf_1
Xmax_cap27 _0163_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0811_ _0162_ _0183_ _0185_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__o21ba_2
Xinput12 keypad_i[5] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1225_ clk8.count\[11\] clk8.count\[10\] _0549_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__and3_1
X_1156_ _0503_ _0331_ _0504_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__and3b_1
X_1087_ osc.count\[3\] _0452_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1010_ _0380_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__buf_2
XFILLER_0_29_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1774_ clknet_4_0_0_clk net12 net28 vssd1 vssd1 vccd1 vccd1 kp_encoder.q\[5\] sky130_fd_sc_hd__dfrtp_1
X_1208_ _0540_ _0541_ _0531_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__and3b_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1139_ net94 clk_div.count\[0\] _0350_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1490_ _0082_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1 kp_encoder.q\[4\] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1688_ clknet_4_11_0_clk _0044_ net38 vssd1 vssd1 vccd1 vccd1 seq_div.D\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1757_ clknet_4_0_0_clk net41 net28 vssd1 vssd1 vccd1 vccd1 kp_encoder.sync_out\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1611_ net73 _0149_ _0150_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0990_ _0360_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__buf_4
X_1473_ net111 _0632_ _0634_ seq_div.R\[22\] vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__a22o_1
X_1542_ seq_div.D\[13\] _0109_ _0631_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0973_ kp_encoder.sync_out\[9\] _0337_ _0341_ _0343_ vssd1 vssd1 vccd1 vccd1 _0344_
+ sky130_fd_sc_hd__a211o_2
X_1456_ net117 _0632_ _0634_ seq_div.R\[19\] vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__a22o_1
X_1387_ _0653_ _0698_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__nand2_1
X_1525_ _0098_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1241_ _0563_ _0531_ _0564_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__and3b_1
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1310_ _0624_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__clkbuf_4
X_1172_ pwm.count\[4\] pwm.count\[3\] _0510_ _0350_ vssd1 vssd1 vccd1 vccd1 _0515_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0956_ SS_FSM.count\[5\] _0302_ _0219_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0887_ _0179_ _0183_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__nor2_1
X_1508_ seq_div.D\[1\] _0087_ _0632_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__mux2_1
X_1439_ _0692_ _0741_ _0706_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput13 keypad_i[6] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_1
X_0810_ _0184_ _0160_ _0161_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1224_ net110 _0549_ _0552_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[10\] sky130_fd_sc_hd__o21ba_1
X_1155_ clk_div.count\[6\] _0500_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__or2_1
X_1086_ _0454_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0939_ _0189_ _0186_ _0178_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1773_ clknet_4_7_0_clk _0079_ net36 vssd1 vssd1 vccd1 vccd1 mode_FSM.mode\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1207_ clk8.count\[3\] clk8.count\[4\] _0534_ clk8.count\[5\] vssd1 vssd1 vccd1 vccd1
+ _0541_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1138_ _0350_ net64 vssd1 vssd1 vccd1 vccd1 clk_div.next_count\[0\] sky130_fd_sc_hd__nor2_1
XFILLER_0_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1069_ _0382_ _0375_ _0391_ _0439_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2 kp_encoder.q\[3\] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1756_ clknet_4_2_0_clk net39 net28 vssd1 vssd1 vccd1 vccd1 kp_encoder.sync_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1687_ clknet_4_9_0_clk _0043_ net34 vssd1 vssd1 vccd1 vccd1 seq_div.D\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1610_ seq_div.count_div\[0\] seq_div.count_div\[1\] net57 _0625_ vssd1 vssd1 vccd1
+ vccd1 _0150_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1472_ _0769_ seq_div.R\[21\] _0707_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__mux2_1
X_1541_ _0387_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1739_ clknet_4_4_0_clk clk8.next_count\[8\] net29 vssd1 vssd1 vccd1 vccd1 clk8.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0972_ _0342_ _0335_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1524_ seq_div.D\[7\] _0419_ _0632_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__mux2_1
X_1455_ _0755_ seq_div.R\[18\] _0707_ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__mux2_1
X_1386_ seq_div.D\[6\] seq_div.R\[13\] vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__or2b_1
XFILLER_0_60_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1240_ clk8.count\[15\] _0560_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__or2_1
X_1171_ _0513_ _0514_ vssd1 vssd1 vccd1 vccd1 pwm.next_count\[3\] sky130_fd_sc_hd__nor2_1
XFILLER_0_47_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0955_ _0297_ _0313_ _0326_ _0237_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0886_ _0247_ _0259_ _0217_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1507_ _0427_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1369_ _0677_ _0680_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1438_ _0692_ _0741_ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 keypad_i[7] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
X_1223_ clk8.count\[9\] clk8.count\[10\] _0546_ _0350_ vssd1 vssd1 vccd1 vccd1 _0552_
+ sky130_fd_sc_hd__a31o_1
X_1154_ clk_div.count\[6\] _0500_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1085_ _0452_ _0417_ _0448_ _0453_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__and4b_1
XFILLER_0_23_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0869_ _0154_ _0242_ _0159_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__a21o_1
X_0938_ _0305_ _0309_ _0214_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1772_ clknet_4_7_0_clk _0078_ net36 vssd1 vssd1 vccd1 vccd1 mode_FSM.mode\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1206_ clk8.count\[4\] clk8.count\[5\] _0537_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__and3_1
X_1137_ _0492_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[15\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1068_ osc.count\[6\] vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 kp_encoder.q\[5\] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1755_ clknet_4_2_0_clk net40 net28 vssd1 vssd1 vccd1 vccd1 kp_encoder.sync_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1686_ clknet_4_11_0_clk _0042_ net34 vssd1 vssd1 vccd1 vccd1 seq_div.D\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1540_ _0108_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1471_ _0674_ _0768_ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1669_ clknet_4_13_0_clk _0025_ net36 vssd1 vssd1 vccd1 vccd1 seq_div.q_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1738_ clknet_4_5_0_clk clk8.next_count\[7\] net29 vssd1 vssd1 vccd1 vccd1 clk8.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0971_ kp_encoder.sync_out\[11\] vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1454_ _0664_ _0754_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__xnor2_1
X_1523_ net87 _0632_ _0097_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1385_ seq_div.R\[14\] seq_div.D\[7\] vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1170_ pwm.count\[3\] _0510_ _0331_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0954_ _0321_ _0325_ _0232_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0885_ _0252_ _0258_ _0214_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1506_ _0430_ _0712_ _0086_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__o21ai_1
X_1437_ _0638_ _0736_ _0655_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__a21oi_1
X_1299_ pwm.count\[0\] _0592_ _0610_ _0614_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__or4_1
X_1368_ _0678_ seq_div.R\[22\] _0668_ _0679_ _0672_ vssd1 vssd1 vccd1 vccd1 _0680_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput15 keypad_i[8] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1222_ _0551_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[9\] sky130_fd_sc_hd__clkbuf_1
X_1153_ _0502_ vssd1 vssd1 vccd1 vccd1 clk_div.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
X_1084_ osc.count\[0\] osc.count\[1\] osc.count\[2\] vssd1 vssd1 vccd1 vccd1 _0453_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0799_ net27 _0172_ _0173_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__and3_1
X_0868_ _0206_ _0186_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__nor2_1
X_0937_ _0167_ _0306_ _0308_ _0178_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1771_ clknet_4_0_0_clk net11 net28 vssd1 vssd1 vccd1 vccd1 kp_encoder.q\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1205_ net103 _0537_ _0539_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[4\] sky130_fd_sc_hd__o21a_1
X_1136_ _0331_ _0417_ _0448_ _0491_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__and4_1
X_1067_ osc.count\[6\] _0373_ _0437_ _0435_ osc.count\[5\] vssd1 vssd1 vccd1 vccd1
+ _0438_ sky130_fd_sc_hd__o32a_1
XFILLER_0_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4 kp_encoder.q\[10\] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1754_ clknet_4_8_0_clk net48 net33 vssd1 vssd1 vccd1 vccd1 kp_encoder.sync_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1685_ clknet_4_11_0_clk _0041_ net34 vssd1 vssd1 vccd1 vccd1 seq_div.D\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1119_ osc.count\[11\] osc.count\[10\] _0473_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1470_ _0668_ _0764_ _0669_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1668_ clknet_4_13_0_clk _0024_ net36 vssd1 vssd1 vccd1 vccd1 seq_div.q_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1737_ clknet_4_4_0_clk clk8.next_count\[6\] net29 vssd1 vssd1 vccd1 vccd1 clk8.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1599_ net125 osc.count\[11\] _0132_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0970_ _0340_ _0336_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__nand2_1
X_1453_ _0749_ _0750_ _0658_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__a21o_1
X_1522_ _0382_ _0375_ _0391_ _0712_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1384_ seq_div.D\[0\] _0675_ _0695_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__or3b_1
XFILLER_0_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0953_ _0284_ _0324_ _0176_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0884_ _0167_ _0254_ _0255_ _0257_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__o31a_1
X_1367_ seq_div.D\[14\] seq_div.R\[21\] vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__and2b_1
X_1505_ net104 _0712_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__nand2_1
X_1436_ net98 _0712_ _0739_ _0625_ _0740_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__o221a_1
X_1298_ seq_div.q_out\[1\] _0588_ _0613_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput16 keypad_i[9] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1221_ _0549_ _0531_ _0550_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__and3b_1
X_1152_ _0500_ _0331_ _0501_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__and3b_1
X_1083_ osc.count\[0\] osc.count\[2\] osc.count\[1\] vssd1 vssd1 vccd1 vccd1 _0452_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0936_ _0165_ _0229_ _0212_ _0307_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0798_ SS_FSM.count\[4\] SS_FSM.count\[5\] SS_FSM.count\[8\] vssd1 vssd1 vccd1 vccd1
+ _0173_ sky130_fd_sc_hd__nor3_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0867_ _0159_ _0213_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1419_ net83 _0712_ _0725_ _0625_ _0726_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__o221a_1
XFILLER_0_21_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1770_ clknet_4_2_0_clk net10 net28 vssd1 vssd1 vccd1 vccd1 kp_encoder.q\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1204_ clk8.count\[4\] _0537_ _0350_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1135_ osc.count\[15\] _0488_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__xnor2_1
X_1066_ _0375_ _0391_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0919_ _0179_ SS_FSM.count\[2\] _0196_ _0155_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5 kp_encoder.q\[13\] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1753_ clknet_4_2_0_clk net53 net28 vssd1 vssd1 vccd1 vccd1 kp_encoder.sync_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1684_ clknet_4_10_0_clk _0040_ net34 vssd1 vssd1 vccd1 vccd1 seq_div.D\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1118_ _0478_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[10\] sky130_fd_sc_hd__clkbuf_1
X_1049_ _0382_ _0361_ _0370_ _0351_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__o31a_2
XFILLER_0_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1736_ clknet_4_4_0_clk clk8.next_count\[5\] net29 vssd1 vssd1 vccd1 vccd1 clk8.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1667_ clknet_4_15_0_clk _0023_ net37 vssd1 vssd1 vccd1 vccd1 seq_div.q_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1598_ _0143_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1452_ net91 _0712_ _0717_ seq_div.R\[18\] _0753_ vssd1 vssd1 vccd1 vccd1 _0013_
+ sky130_fd_sc_hd__o221a_1
X_1383_ _0642_ _0694_ vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1521_ _0096_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1719_ clknet_4_12_0_clk _0075_ net35 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0952_ _0230_ _0323_ _0159_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__a21oi_1
X_1504_ seq_div.Q\[6\] _0628_ _0634_ net59 vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0883_ _0228_ _0256_ _0159_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__o21a_1
X_1366_ seq_div.D\[15\] vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__inv_2
X_1435_ seq_div.R\[15\] _0717_ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1297_ _0582_ _0611_ _0612_ _0591_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
Xinput17 n_rst vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_2
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1220_ clk8.count\[9\] _0546_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__or2_1
X_1151_ clk_div.count\[3\] clk_div.count\[4\] _0494_ clk_div.count\[5\] vssd1 vssd1
+ vccd1 vccd1 _0501_ sky130_fd_sc_hd__a31o_1
X_1082_ _0451_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
X_0935_ _0179_ _0162_ _0228_ _0183_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0866_ _0154_ _0159_ _0168_ _0239_ _0240_ vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__a311o_1
X_0797_ SS_FSM.count\[6\] SS_FSM.count\[7\] vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1349_ _0659_ _0660_ _0640_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1418_ seq_div.R\[12\] _0717_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1134_ _0490_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
X_1203_ net90 _0534_ _0538_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[3\] sky130_fd_sc_hd__o21a_1
XFILLER_0_47_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1065_ osc.count\[4\] _0381_ _0392_ _0435_ osc.count\[5\] vssd1 vssd1 vccd1 vccd1
+ _0436_ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0849_ _0219_ _0222_ _0223_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__nand3_1
X_0918_ _0249_ _0250_ SS_FSM.count\[5\] _0167_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6 kp_encoder.q\[7\] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1752_ clknet_4_8_0_clk net49 net28 vssd1 vssd1 vccd1 vccd1 kp_encoder.sync_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1683_ clknet_4_10_0_clk _0039_ net34 vssd1 vssd1 vccd1 vccd1 seq_div.D\[4\] sky130_fd_sc_hd__dfrtp_1
X_1117_ _0476_ _0417_ _0448_ _0477_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__and4b_1
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1048_ _0383_ _0381_ _0386_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__nand3_2
XFILLER_0_31_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1666_ clknet_4_13_0_clk _0022_ net36 vssd1 vssd1 vccd1 vccd1 seq_div.q_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1735_ clknet_4_4_0_clk clk8.next_count\[4\] net29 vssd1 vssd1 vccd1 vccd1 clk8.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1597_ net91 osc.count\[10\] _0132_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1520_ net118 _0095_ _0632_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__mux2_1
X_1451_ seq_div.R\[17\] _0707_ _0751_ _0752_ _0625_ vssd1 vssd1 vccd1 vccd1 _0753_
+ sky130_fd_sc_hd__a221o_1
X_1382_ seq_div.R\[8\] seq_div.D\[1\] vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__or2b_1
XFILLER_0_10_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1718_ clknet_4_6_0_clk _0074_ net35 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1649_ clknet_4_12_0_clk osc.next_count\[10\] net35 vssd1 vssd1 vccd1 vccd1 osc.count\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0882_ _0155_ _0196_ SS_FSM.count\[2\] _0179_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__a211o_1
X_0951_ _0322_ _0250_ _0167_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__o21ai_1
X_1503_ net62 _0628_ _0634_ seq_div.Q\[6\] vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1296_ _0585_ seq_div.q_out\[0\] vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1365_ _0667_ _0675_ _0676_ vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__or3b_1
X_1434_ seq_div.R\[14\] _0707_ _0737_ _0738_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__a22o_1
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1150_ clk_div.count\[5\] clk_div.count\[4\] _0497_ vssd1 vssd1 vccd1 vccd1 _0500_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1081_ _0417_ _0448_ _0449_ _0450_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__and4_1
X_0865_ SS_FSM.sound\[0\] vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0934_ _0165_ _0229_ _0212_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__o21ai_1
X_0796_ SS_FSM.count\[7\] _0170_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1417_ _0724_ seq_div.R\[11\] _0707_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1279_ _0585_ seq_div.q_out\[4\] vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__nand2_1
X_1348_ seq_div.D\[8\] seq_div.R\[15\] vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__or2b_1
XFILLER_0_56_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1133_ _0417_ _0448_ _0488_ _0489_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__and4_1
X_1202_ _0350_ _0537_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__nor2_1
Xclkbuf_4_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_1064_ _0373_ _0429_ _0379_ _0378_ _0406_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_47_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0917_ _0202_ _0289_ _0178_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__a21oi_1
X_0779_ SS_FSM.count\[0\] vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__inv_2
X_0848_ net27 _0172_ _0173_ _0179_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7 kp_encoder.q\[6\] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1751_ clknet_4_5_0_clk clk8.next_count\[20\] net32 vssd1 vssd1 vccd1 vccd1 clk8.count\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_1682_ clknet_4_8_0_clk _0038_ net33 vssd1 vssd1 vccd1 vccd1 seq_div.D\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1116_ osc.count\[10\] _0473_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__or2_1
X_1047_ osc.count\[7\] vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1665_ clknet_4_13_0_clk _0021_ net35 vssd1 vssd1 vccd1 vccd1 seq_div.q_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1734_ clknet_4_4_0_clk clk8.next_count\[3\] net29 vssd1 vssd1 vccd1 vccd1 clk8.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1596_ _0142_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1450_ _0749_ _0750_ _0706_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__a21oi_1
X_1381_ _0690_ _0691_ _0692_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1717_ clknet_4_6_0_clk _0073_ net35 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1648_ clknet_4_9_0_clk osc.next_count\[9\] net33 vssd1 vssd1 vccd1 vccd1 osc.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1579_ net126 osc.count\[1\] _0132_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0881_ _0224_ _0198_ _0165_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__a21oi_1
X_0950_ _0190_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1502_ net77 _0628_ _0634_ net62 vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__a22o_1
X_1433_ _0735_ _0736_ _0706_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__a21oi_1
X_1295_ _0585_ seq_div.q_out\[0\] vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1364_ seq_div.D\[12\] seq_div.R\[19\] vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1080_ osc.count\[0\] osc.count\[1\] vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0795_ _0169_ net25 vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0933_ _0242_ _0246_ _0178_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__o21ai_1
X_0864_ _0175_ _0218_ _0233_ _0238_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__o31a_1
X_1347_ seq_div.D\[9\] _0639_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__or2_1
X_1416_ _0687_ _0723_ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__xor2_1
X_1278_ _0585_ seq_div.q_out\[4\] vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1201_ clk8.count\[3\] _0534_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1132_ osc.count\[14\] _0485_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1063_ _0381_ _0392_ osc.count\[4\] vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0916_ _0195_ _0197_ _0288_ _0167_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0847_ _0179_ _0155_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold8 kp_encoder.q\[14\] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dlygate4sd3_1
X_1750_ clknet_4_5_0_clk clk8.next_count\[19\] net32 vssd1 vssd1 vccd1 vccd1 clk8.count\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1681_ clknet_4_8_0_clk _0037_ net33 vssd1 vssd1 vccd1 vccd1 seq_div.D\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1046_ _0405_ _0414_ _0415_ _0416_ _0400_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__o2111a_4
X_1115_ osc.count\[10\] _0473_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1733_ clknet_4_4_0_clk clk8.next_count\[2\] net29 vssd1 vssd1 vccd1 vccd1 clk8.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1664_ clknet_4_13_0_clk _0020_ net35 vssd1 vssd1 vccd1 vccd1 seq_div.q_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1595_ net88 osc.count\[9\] _0132_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1029_ osc.count\[15\] _0398_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1380_ _0637_ _0660_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__nand2_1
X_1716_ clknet_4_12_0_clk _0072_ net35 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1578_ _0133_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1647_ clknet_4_9_0_clk osc.next_count\[8\] net33 vssd1 vssd1 vccd1 vccd1 osc.count\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0880_ _0184_ SS_FSM.count\[5\] _0253_ _0198_ _0224_ vssd1 vssd1 vccd1 vccd1 _0254_
+ sky130_fd_sc_hd__o311a_1
X_1501_ net75 _0628_ _0634_ net77 vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__a22o_1
X_1363_ _0671_ _0674_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__or2_1
X_1432_ _0735_ _0736_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__or2_1
X_1294_ mode_FSM.mode\[1\] seq_div.q_out\[0\] vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0932_ _0274_ _0298_ _0299_ _0304_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__a22oi_4
XFILLER_0_23_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0794_ SS_FSM.count\[6\] vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__inv_2
X_0863_ _0175_ _0235_ _0237_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1346_ seq_div.D\[10\] seq_div.R\[17\] vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__and2b_1
X_1415_ _0648_ _0719_ _0644_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__a21oi_1
X_1277_ seq_div.q_out\[6\] _0588_ _0590_ _0592_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1200_ _0536_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
X_1131_ osc.count\[14\] _0485_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__nand2_1
X_1062_ _0428_ _0431_ _0432_ _0423_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0915_ _0189_ _0198_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__or2_1
X_0846_ _0159_ _0220_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1329_ _0637_ _0638_ _0640_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold9 kp_encoder.q\[11\] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1680_ clknet_4_10_0_clk _0036_ net34 vssd1 vssd1 vccd1 vccd1 seq_div.D\[1\] sky130_fd_sc_hd__dfrtp_1
X_1114_ _0475_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[9\] sky130_fd_sc_hd__clkbuf_1
X_1045_ _0399_ _0402_ osc.count\[14\] vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__or3b_1
XFILLER_0_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0829_ _0178_ _0187_ _0192_ _0203_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1663_ clknet_4_6_0_clk _0019_ net35 vssd1 vssd1 vccd1 vccd1 seq_div.q_out\[0\] sky130_fd_sc_hd__dfrtp_1
X_1732_ clknet_4_4_0_clk net66 net29 vssd1 vssd1 vccd1 vccd1 clk8.count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1594_ _0141_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__clkbuf_1
X_1028_ osc.count\[15\] _0398_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1715_ clknet_4_12_0_clk _0071_ net35 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1646_ clknet_4_9_0_clk osc.next_count\[7\] net33 vssd1 vssd1 vccd1 vccd1 osc.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1577_ net123 osc.count\[0\] _0132_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1500_ seq_div.Q\[2\] _0628_ _0634_ net75 vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__a22o_1
X_1293_ seq_div.q_out\[2\] _0588_ _0608_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__o21ai_1
X_1362_ _0672_ _0673_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__nand2_1
X_1431_ _0653_ _0731_ _0656_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1629_ clknet_4_10_0_clk _0009_ net34 vssd1 vssd1 vccd1 vccd1 seq_div.R\[14\] sky130_fd_sc_hd__dfrtp_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0862_ SS_FSM.sound\[0\] _0236_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0931_ _0189_ _0300_ _0301_ _0303_ _0228_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0793_ _0162_ _0165_ _0167_ SS_FSM.sound\[1\] vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__o211a_1
X_1276_ _0591_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1414_ _0628_ _0721_ _0722_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__a21o_1
X_1345_ _0652_ _0653_ _0654_ _0655_ _0656_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__a311o_1
XFILLER_0_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1130_ _0487_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[13\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1061_ osc.count\[3\] _0420_ _0422_ osc.count\[2\] vssd1 vssd1 vccd1 vccd1 _0432_
+ sky130_fd_sc_hd__o22ai_1
XFILLER_0_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0845_ _0219_ _0165_ _0174_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__a21o_1
X_0914_ _0214_ _0284_ _0286_ _0232_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__o31a_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1259_ kp_encoder.last_sk kp_encoder.sync_out\[14\] vssd1 vssd1 vccd1 vccd1 _0577_
+ sky130_fd_sc_hd__and2b_1
X_1328_ seq_div.D\[9\] _0639_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1044_ _0388_ _0404_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__nand2_1
X_1113_ _0473_ _0417_ _0448_ _0474_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__and4b_1
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0828_ _0194_ _0201_ _0202_ _0159_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1731_ clknet_4_4_0_clk clk8.next_count\[0\] net29 vssd1 vssd1 vccd1 vccd1 clk8.count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_1662_ clknet_4_6_0_clk clk_div.next_count\[7\] net30 vssd1 vssd1 vccd1 vccd1 clk_div.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1593_ net99 osc.count\[8\] _0132_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__mux2_1
X_1027_ _0382_ _0397_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold90 seq_div.dividend\[2\] vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1576_ _0350_ _0507_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__nor2_8
X_1714_ clknet_4_9_0_clk _0070_ net35 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1645_ clknet_4_2_0_clk osc.next_count\[6\] net28 vssd1 vssd1 vccd1 vccd1 osc.count\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1430_ _0697_ _0655_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__nor2_1
X_1292_ _0582_ _0606_ _0607_ _0591_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__a31o_1
X_1361_ seq_div.D\[14\] seq_div.R\[21\] vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__or2b_1
XFILLER_0_37_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1559_ _0240_ _0114_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__or2_1
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1628_ clknet_4_10_0_clk _0008_ net34 vssd1 vssd1 vccd1 vccd1 seq_div.R\[13\] sky130_fd_sc_hd__dfrtp_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0861_ SS_FSM.sound\[1\] vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__inv_2
X_0792_ _0166_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__buf_4
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0930_ SS_FSM.count\[5\] _0162_ _0302_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__or3b_1
XFILLER_0_2_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1413_ seq_div.dividend\[3\] _0632_ _0634_ seq_div.R\[11\] vssd1 vssd1 vccd1 vccd1
+ _0722_ sky130_fd_sc_hd__a22o_1
X_1275_ _0581_ _0585_ mode_FSM.mode\[0\] vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__o21ba_2
X_1344_ seq_div.D\[6\] seq_div.R\[13\] vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1060_ osc.count\[1\] _0427_ _0430_ osc.count\[0\] vssd1 vssd1 vccd1 vccd1 _0431_
+ sky130_fd_sc_hd__o22ai_1
XFILLER_0_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0844_ _0160_ _0161_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__nand2_2
X_0913_ _0159_ _0285_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1258_ net56 _0573_ _0576_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[20\] sky130_fd_sc_hd__a21oi_1
X_1189_ _0524_ _0525_ _0526_ _0527_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__and4b_1
X_1327_ seq_div.R\[16\] vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1043_ _0409_ _0412_ _0413_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__a21oi_1
X_1112_ osc.count\[9\] _0470_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0827_ _0167_ _0194_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1730_ clknet_4_7_0_clk pwm.next_count\[7\] net31 vssd1 vssd1 vccd1 vccd1 pwm.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1661_ clknet_4_6_0_clk clk_div.next_count\[6\] net30 vssd1 vssd1 vccd1 vccd1 clk_div.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1592_ _0140_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1026_ _0351_ _0361_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold91 seq_div.dividend\[13\] vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 seq_div.D\[5\] vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dlygate4sd3_1
X_1713_ clknet_4_9_0_clk _0069_ net38 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1575_ net116 _0123_ _0131_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__o21a_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1644_ clknet_4_8_0_clk osc.next_count\[5\] net33 vssd1 vssd1 vccd1 vccd1 osc.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1009_ _0373_ _0361_ _0377_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__or3_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1360_ seq_div.R\[21\] seq_div.D\[14\] vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__or2b_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1291_ _0585_ seq_div.q_out\[1\] vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1489_ net121 seq_div.q_out\[4\] _0776_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__mux2_1
X_1558_ _0219_ net23 _0117_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__or3b_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1627_ clknet_4_10_0_clk _0007_ net34 vssd1 vssd1 vccd1 vccd1 seq_div.R\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0860_ _0219_ _0234_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__or2_1
X_0791_ SS_FSM.count\[4\] net27 vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1412_ _0720_ seq_div.R\[10\] _0707_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__mux2_1
X_1343_ seq_div.D\[7\] seq_div.R\[14\] vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__and2b_1
X_1274_ _0585_ seq_div.q_out\[5\] _0589_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0989_ _0352_ _0353_ _0359_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0912_ _0179_ _0193_ _0228_ _0269_ _0209_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__o311a_1
XFILLER_0_59_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0843_ _0176_ _0204_ _0208_ _0215_ _0217_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__o221a_1
X_1326_ seq_div.R\[14\] seq_div.D\[7\] vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__or2b_1
X_1257_ net56 _0573_ _0531_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__o21ai_1
X_1188_ clk8.count\[19\] clk8.count\[18\] clk8.count\[17\] vssd1 vssd1 vccd1 vccd1
+ _0527_ sky130_fd_sc_hd__and3b_1
XFILLER_0_19_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1042_ osc.count\[11\] _0395_ _0411_ osc.count\[10\] vssd1 vssd1 vccd1 vccd1 _0413_
+ sky130_fd_sc_hd__a22o_1
X_1111_ osc.count\[9\] osc.count\[8\] _0467_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0826_ _0195_ _0197_ _0200_ _0167_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__a31o_1
X_1309_ _0623_ seq_div.state\[0\] vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_15_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1660_ clknet_4_6_0_clk clk_div.next_count\[5\] net30 vssd1 vssd1 vccd1 vccd1 clk_div.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1591_ net98 osc.count\[7\] _0132_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__mux2_1
X_1025_ osc.count\[11\] _0395_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0809_ _0155_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold92 seq_div.dividend\[14\] vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 seq_div.R\[23\] vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 seq_div.D\[10\] vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1643_ clknet_4_8_0_clk osc.next_count\[4\] net33 vssd1 vssd1 vccd1 vccd1 osc.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_1712_ clknet_4_9_0_clk _0068_ net38 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1574_ _0236_ _0175_ _0120_ _0127_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__a211o_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1008_ _0361_ _0377_ _0351_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1290_ _0585_ seq_div.q_out\[1\] vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1626_ clknet_4_10_0_clk _0006_ net34 vssd1 vssd1 vccd1 vccd1 seq_div.R\[11\] sky130_fd_sc_hd__dfrtp_1
X_1488_ _0081_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__clkbuf_1
X_1557_ SS_FSM.sound\[1\] _0180_ _0181_ _0269_ SS_FSM.sound\[0\] vssd1 vssd1 vccd1
+ vccd1 _0120_ sky130_fd_sc_hd__o41ai_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0790_ _0163_ _0164_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__nor2_8
XFILLER_0_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1273_ _0585_ seq_div.q_out\[5\] _0582_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__o21ai_1
X_1411_ _0684_ _0719_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__xnor2_1
X_1342_ seq_div.R\[12\] seq_div.D\[5\] vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0988_ _0344_ _0346_ _0358_ _0350_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__a31o_1
X_1609_ seq_div.state\[0\] _0132_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0842_ _0171_ _0216_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__and2_1
X_0911_ _0211_ _0283_ _0178_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1256_ _0575_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[19\] sky130_fd_sc_hd__clkbuf_1
X_1325_ seq_div.R\[15\] seq_div.D\[8\] vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__or2b_1
X_1187_ clk8.count\[16\] clk8.count\[20\] clk8.count\[14\] clk8.count\[15\] vssd1
+ vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__and4b_1
XFILLER_0_19_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1110_ _0472_ vssd1 vssd1 vccd1 vccd1 osc.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1041_ osc.count\[9\] _0408_ _0411_ osc.count\[10\] vssd1 vssd1 vccd1 vccd1 _0412_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0825_ _0198_ _0199_ _0189_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1239_ clk8.count\[15\] _0560_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__and2_1
X_1308_ seq_div.state\[1\] vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1590_ _0139_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1024_ _0390_ _0392_ _0393_ _0394_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0808_ _0156_ _0180_ _0181_ _0182_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__o31a_2
XFILLER_0_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold82 seq_div.Q\[0\] vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 _0775_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 seq_div.dividend\[7\] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_14_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1642_ clknet_4_8_0_clk osc.next_count\[3\] net33 vssd1 vssd1 vccd1 vccd1 osc.count\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_1711_ clknet_4_9_0_clk _0067_ net38 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ net112 _0123_ _0127_ _0130_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__o22a_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1007_ _0361_ _0377_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__nor2_2
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1625_ clknet_4_10_0_clk _0005_ net34 vssd1 vssd1 vccd1 vccd1 seq_div.R\[10\] sky130_fd_sc_hd__dfrtp_1
X_1556_ _0182_ _0117_ _0119_ _0115_ _0155_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__a32o_1
X_1487_ net122 seq_div.q_out\[3\] _0776_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__mux2_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1410_ _0643_ _0714_ _0645_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1272_ _0587_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1341_ seq_div.R\[13\] seq_div.D\[6\] vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0987_ _0354_ kp_encoder.sync_out\[10\] _0337_ _0343_ _0357_ vssd1 vssd1 vccd1 vccd1
+ _0358_ sky130_fd_sc_hd__a311o_1
X_1608_ _0148_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__clkbuf_1
X_1539_ net115 _0107_ _0631_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0841_ SS_FSM.count\[7\] _0170_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__nand2_1
X_0910_ _0179_ _0165_ _0166_ _0186_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1255_ _0573_ _0331_ _0574_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__and3b_1
X_1186_ clk8.count\[7\] clk8.count\[6\] clk8.count\[9\] clk8.count\[8\] vssd1 vssd1
+ vccd1 vccd1 _0525_ sky130_fd_sc_hd__and4b_1
X_1324_ seq_div.R\[17\] seq_div.D\[10\] vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__or2b_1
XFILLER_0_46_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1040_ _0382_ _0375_ _0410_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0824_ _0160_ _0161_ _0155_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1307_ net61 _0586_ _0622_ _0350_ vssd1 vssd1 vccd1 vccd1 pwm.pwm sky130_fd_sc_hd__a211oi_1
X_1238_ _0562_ vssd1 vssd1 vccd1 vccd1 clk8.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
X_1169_ pwm.count\[3\] _0510_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1023_ _0370_ _0383_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0807_ SS_FSM.count\[0\] _0155_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold83 seq_div.Q\[4\] vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 clk8.count\[10\] vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 seq_div.dividend\[9\] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 seq_div.dividend\[8\] vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1572_ _0237_ _0217_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1641_ clknet_4_8_0_clk osc.next_count\[2\] net33 vssd1 vssd1 vccd1 vccd1 osc.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1710_ clknet_4_11_0_clk _0066_ net38 vssd1 vssd1 vccd1 vccd1 seq_div.dividend\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1006_ _0352_ _0362_ _0369_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__a21o_2
XFILLER_0_32_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1555_ _0179_ _0115_ _0118_ _0119_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__a22o_1
X_1624_ clknet_4_10_0_clk _0004_ net34 vssd1 vssd1 vccd1 vccd1 seq_div.R\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1486_ _0080_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__clkbuf_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_13_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1340_ _0649_ _0650_ _0651_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__or3b_1
X_1271_ mode_FSM.mode\[1\] mode_FSM.mode\[0\] vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0986_ _0355_ _0339_ _0356_ kp_encoder.sync_out\[1\] kp_encoder.sync_out\[0\] vssd1
+ vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_14_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1469_ _0628_ _0766_ _0767_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__a21o_1
X_1607_ seq_div.dividend\[15\] osc.count\[15\] _0132_ vssd1 vssd1 vccd1 vccd1 _0148_
+ sky130_fd_sc_hd__mux2_1
X_1538_ _0385_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0840_ _0209_ _0178_ _0211_ _0213_ _0214_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__a41o_1
X_1323_ seq_div.R\[18\] seq_div.D\[11\] vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__or2b_1
X_1254_ clk8.count\[19\] _0570_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__or2_1
X_1185_ clk8.count\[11\] clk8.count\[10\] clk8.count\[12\] clk8.count\[13\] vssd1
+ vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__or4b_1
XFILLER_0_46_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0969_ kp_encoder.sync_out\[9\] _0338_ _0332_ _0339_ _0337_ vssd1 vssd1 vccd1 vccd1
+ _0340_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0823_ SS_FSM.count\[0\] _0184_ SS_FSM.count\[2\] vssd1 vssd1 vccd1 vccd1 _0198_
+ sky130_fd_sc_hd__or3_2
X_1306_ pwm.count\[6\] _0593_ _0586_ net67 _0621_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__o221a_1
X_1237_ _0560_ _0531_ _0561_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__and3b_1
X_1168_ _0512_ vssd1 vssd1 vccd1 vccd1 pwm.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
X_1099_ osc.count\[6\] _0461_ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1022_ _0375_ _0381_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0806_ SS_FSM.count\[4\] SS_FSM.count\[5\] SS_FSM.count\[8\] vssd1 vssd1 vccd1 vccd1
+ _0181_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold40 seq_div.dividend\[6\] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 seq_div.Q\[3\] vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 seq_div.dividend\[14\] vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 _0012_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 _0011_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1571_ SS_FSM.count\[6\] _0123_ _0127_ _0129_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__o22a_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1640_ clknet_4_8_0_clk osc.next_count\[1\] net33 vssd1 vssd1 vccd1 vccd1 osc.count\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1005_ _0375_ _0361_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1769_ clknet_4_8_0_clk net9 net28 vssd1 vssd1 vccd1 vccd1 kp_encoder.q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1485_ seq_div.Q\[2\] seq_div.q_out\[2\] _0776_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1554_ SS_FSM.sound\[0\] _0114_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__and2_1
X_1623_ clknet_4_8_0_clk net69 net34 vssd1 vssd1 vccd1 vccd1 seq_div.R\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

