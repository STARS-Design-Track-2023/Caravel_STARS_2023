magic
tech sky130A
magscale 1 2
timestamp 1693932206
<< viali >>
rect 6745 30345 6779 30379
rect 10241 30277 10275 30311
rect 22293 30277 22327 30311
rect 25697 30277 25731 30311
rect 1593 30209 1627 30243
rect 2789 30209 2823 30243
rect 6653 30209 6687 30243
rect 9873 30209 9907 30243
rect 14197 30209 14231 30243
rect 17601 30209 17635 30243
rect 21925 30209 21959 30243
rect 25329 30209 25363 30243
rect 28365 30209 28399 30243
rect 28733 30209 28767 30243
rect 29009 30141 29043 30175
rect 2973 30073 3007 30107
rect 14381 30073 14415 30107
rect 17785 30073 17819 30107
rect 1409 30005 1443 30039
rect 28549 30005 28583 30039
rect 23673 29801 23707 29835
rect 5641 29665 5675 29699
rect 16773 29665 16807 29699
rect 5089 29597 5123 29631
rect 5457 29597 5491 29631
rect 5549 29597 5583 29631
rect 5733 29597 5767 29631
rect 9045 29597 9079 29631
rect 11253 29597 11287 29631
rect 14749 29597 14783 29631
rect 16865 29597 16899 29631
rect 17509 29597 17543 29631
rect 20821 29597 20855 29631
rect 23857 29597 23891 29631
rect 7389 29529 7423 29563
rect 7573 29529 7607 29563
rect 9413 29529 9447 29563
rect 15117 29529 15151 29563
rect 4905 29461 4939 29495
rect 5273 29461 5307 29495
rect 7757 29461 7791 29495
rect 11805 29461 11839 29495
rect 17233 29461 17267 29495
rect 17325 29461 17359 29495
rect 20637 29461 20671 29495
rect 13277 29257 13311 29291
rect 16497 29257 16531 29291
rect 19165 29257 19199 29291
rect 1685 29189 1719 29223
rect 8769 29189 8803 29223
rect 16957 29189 16991 29223
rect 20177 29189 20211 29223
rect 24041 29189 24075 29223
rect 1409 29121 1443 29155
rect 3249 29121 3283 29155
rect 6837 29121 6871 29155
rect 8953 29121 8987 29155
rect 9045 29121 9079 29155
rect 10701 29121 10735 29155
rect 11345 29121 11379 29155
rect 16221 29121 16255 29155
rect 16313 29121 16347 29155
rect 19901 29121 19935 29155
rect 22661 29121 22695 29155
rect 23121 29121 23155 29155
rect 23305 29121 23339 29155
rect 24409 29121 24443 29155
rect 3525 29053 3559 29087
rect 5089 29053 5123 29087
rect 6929 29053 6963 29087
rect 7205 29053 7239 29087
rect 8677 29053 8711 29087
rect 10793 29053 10827 29087
rect 11529 29053 11563 29087
rect 13461 29053 13495 29087
rect 13737 29053 13771 29087
rect 15301 29053 15335 29087
rect 16681 29053 16715 29087
rect 18521 29053 18555 29087
rect 22569 29053 22603 29087
rect 23397 29053 23431 29087
rect 24685 29053 24719 29087
rect 3157 28985 3191 29019
rect 4997 28985 5031 29019
rect 5733 28985 5767 29019
rect 6653 28985 6687 29019
rect 11069 28985 11103 29019
rect 8769 28917 8803 28951
rect 11161 28917 11195 28951
rect 11786 28917 11820 28951
rect 15209 28917 15243 28951
rect 15945 28917 15979 28951
rect 18429 28917 18463 28951
rect 21649 28917 21683 28951
rect 23029 28917 23063 28951
rect 23121 28917 23155 28951
rect 6101 28713 6135 28747
rect 7389 28713 7423 28747
rect 7849 28713 7883 28747
rect 9781 28713 9815 28747
rect 10333 28713 10367 28747
rect 12449 28713 12483 28747
rect 12633 28713 12667 28747
rect 13461 28713 13495 28747
rect 14933 28713 14967 28747
rect 16129 28713 16163 28747
rect 16681 28713 16715 28747
rect 20361 28713 20395 28747
rect 20545 28713 20579 28747
rect 21833 28713 21867 28747
rect 15853 28645 15887 28679
rect 22201 28645 22235 28679
rect 24225 28645 24259 28679
rect 3341 28577 3375 28611
rect 4353 28577 4387 28611
rect 8217 28577 8251 28611
rect 9137 28577 9171 28611
rect 10701 28577 10735 28611
rect 13645 28577 13679 28611
rect 15393 28577 15427 28611
rect 17049 28577 17083 28611
rect 19533 28577 19567 28611
rect 22477 28577 22511 28611
rect 22753 28577 22787 28611
rect 24777 28577 24811 28611
rect 25237 28577 25271 28611
rect 3249 28509 3283 28543
rect 4077 28509 4111 28543
rect 6469 28509 6503 28543
rect 6929 28509 6963 28543
rect 7113 28509 7147 28543
rect 10425 28509 10459 28543
rect 13185 28509 13219 28543
rect 13369 28509 13403 28543
rect 13737 28509 13771 28543
rect 14197 28509 14231 28543
rect 15117 28509 15151 28543
rect 15301 28509 15335 28543
rect 15577 28509 15611 28543
rect 15669 28509 15703 28543
rect 16037 28509 16071 28543
rect 16221 28509 16255 28543
rect 16497 28509 16531 28543
rect 16773 28509 16807 28543
rect 19257 28509 19291 28543
rect 19349 28509 19383 28543
rect 20821 28509 20855 28543
rect 20913 28509 20947 28543
rect 21006 28509 21040 28543
rect 21097 28509 21131 28543
rect 21373 28509 21407 28543
rect 21465 28509 21499 28543
rect 21823 28509 21857 28543
rect 22293 28509 22327 28543
rect 22385 28509 22419 28543
rect 24501 28509 24535 28543
rect 3893 28441 3927 28475
rect 4629 28441 4663 28475
rect 6193 28441 6227 28475
rect 6377 28441 6411 28475
rect 7205 28441 7239 28475
rect 7665 28441 7699 28475
rect 7865 28441 7899 28475
rect 8769 28441 8803 28475
rect 9965 28441 9999 28475
rect 10149 28441 10183 28475
rect 12265 28441 12299 28475
rect 12465 28441 12499 28475
rect 13461 28441 13495 28475
rect 16313 28441 16347 28475
rect 20177 28441 20211 28475
rect 20393 28441 20427 28475
rect 22109 28441 22143 28475
rect 3617 28373 3651 28407
rect 4261 28373 4295 28407
rect 6561 28373 6595 28407
rect 6745 28373 6779 28407
rect 7021 28373 7055 28407
rect 7405 28373 7439 28407
rect 7573 28373 7607 28407
rect 8033 28373 8067 28407
rect 12173 28373 12207 28407
rect 13277 28373 13311 28407
rect 13921 28373 13955 28407
rect 14749 28373 14783 28407
rect 18521 28373 18555 28407
rect 19533 28373 19567 28407
rect 20637 28373 20671 28407
rect 22017 28373 22051 28407
rect 25881 28373 25915 28407
rect 3433 28169 3467 28203
rect 5457 28169 5491 28203
rect 6009 28169 6043 28203
rect 7297 28169 7331 28203
rect 9413 28169 9447 28203
rect 9873 28169 9907 28203
rect 11253 28169 11287 28203
rect 11713 28169 11747 28203
rect 13369 28169 13403 28203
rect 17049 28169 17083 28203
rect 20729 28169 20763 28203
rect 24685 28169 24719 28203
rect 3985 28101 4019 28135
rect 7941 28101 7975 28135
rect 11897 28101 11931 28135
rect 13001 28101 13035 28135
rect 13201 28101 13235 28135
rect 16681 28101 16715 28135
rect 23213 28101 23247 28135
rect 3617 28033 3651 28067
rect 6377 28033 6411 28067
rect 6837 28033 6871 28067
rect 7113 28033 7147 28067
rect 7297 28033 7331 28067
rect 9689 28033 9723 28067
rect 10425 28033 10459 28067
rect 10793 28033 10827 28067
rect 11069 28033 11103 28067
rect 11253 28033 11287 28067
rect 11529 28033 11563 28067
rect 11805 28033 11839 28067
rect 13461 28033 13495 28067
rect 15945 28033 15979 28067
rect 16037 28033 16071 28067
rect 16221 28033 16255 28067
rect 16865 28033 16899 28067
rect 16957 28033 16991 28067
rect 17325 28033 17359 28067
rect 17785 28033 17819 28067
rect 18521 28033 18555 28067
rect 20821 28033 20855 28067
rect 22569 28033 22603 28067
rect 22845 28033 22879 28067
rect 3709 27965 3743 27999
rect 5549 27965 5583 27999
rect 6653 27965 6687 27999
rect 7665 27965 7699 27999
rect 9505 27965 9539 27999
rect 10333 27965 10367 27999
rect 13737 27965 13771 27999
rect 15393 27965 15427 27999
rect 17601 27965 17635 27999
rect 18245 27965 18279 27999
rect 18337 27965 18371 27999
rect 18429 27965 18463 27999
rect 18981 27965 19015 27999
rect 19257 27965 19291 27999
rect 21833 27965 21867 27999
rect 22937 27965 22971 27999
rect 5825 27897 5859 27931
rect 16037 27897 16071 27931
rect 21465 27897 21499 27931
rect 22661 27897 22695 27931
rect 6469 27829 6503 27863
rect 7021 27829 7055 27863
rect 10793 27829 10827 27863
rect 10977 27829 11011 27863
rect 12081 27829 12115 27863
rect 13185 27829 13219 27863
rect 15209 27829 15243 27863
rect 17233 27829 17267 27863
rect 17785 27829 17819 27863
rect 17969 27829 18003 27863
rect 18061 27829 18095 27863
rect 22477 27829 22511 27863
rect 22569 27829 22603 27863
rect 9321 27625 9355 27659
rect 14565 27625 14599 27659
rect 18245 27625 18279 27659
rect 19257 27625 19291 27659
rect 20164 27625 20198 27659
rect 4629 27557 4663 27591
rect 8125 27557 8159 27591
rect 12173 27557 12207 27591
rect 13921 27557 13955 27591
rect 14841 27557 14875 27591
rect 21741 27557 21775 27591
rect 2697 27489 2731 27523
rect 4261 27489 4295 27523
rect 4813 27489 4847 27523
rect 9413 27489 9447 27523
rect 10241 27489 10275 27523
rect 11529 27489 11563 27523
rect 11713 27489 11747 27523
rect 12541 27489 12575 27523
rect 13001 27489 13035 27523
rect 13277 27489 13311 27523
rect 14197 27489 14231 27523
rect 16497 27489 16531 27523
rect 22569 27489 22603 27523
rect 22753 27489 22787 27523
rect 4445 27421 4479 27455
rect 4721 27421 4755 27455
rect 4905 27421 4939 27455
rect 7757 27421 7791 27455
rect 8493 27421 8527 27455
rect 9137 27421 9171 27455
rect 9689 27421 9723 27455
rect 10333 27421 10367 27455
rect 10517 27421 10551 27455
rect 11621 27421 11655 27455
rect 11805 27421 11839 27455
rect 11989 27421 12023 27455
rect 12633 27421 12667 27455
rect 14289 27421 14323 27455
rect 14657 27421 14691 27455
rect 16405 27421 16439 27455
rect 19257 27421 19291 27455
rect 19533 27421 19567 27455
rect 19901 27421 19935 27455
rect 21925 27421 21959 27455
rect 22017 27421 22051 27455
rect 22293 27421 22327 27455
rect 22385 27421 22419 27455
rect 22661 27421 22695 27455
rect 22845 27421 22879 27455
rect 1501 27353 1535 27387
rect 7941 27353 7975 27387
rect 10425 27353 10459 27387
rect 16773 27353 16807 27387
rect 21741 27353 21775 27387
rect 1593 27285 1627 27319
rect 3341 27285 3375 27319
rect 8585 27285 8619 27319
rect 8953 27285 8987 27319
rect 11345 27285 11379 27319
rect 16221 27285 16255 27319
rect 19441 27285 19475 27319
rect 21649 27285 21683 27319
rect 9689 27081 9723 27115
rect 14289 27081 14323 27115
rect 14565 27081 14599 27115
rect 17601 27081 17635 27115
rect 21189 27081 21223 27115
rect 8217 27013 8251 27047
rect 12817 27013 12851 27047
rect 14381 27013 14415 27047
rect 17141 27013 17175 27047
rect 20821 27013 20855 27047
rect 21051 26979 21085 27013
rect 11805 26945 11839 26979
rect 12541 26945 12575 26979
rect 14657 26945 14691 26979
rect 28825 26945 28859 26979
rect 7941 26877 7975 26911
rect 11720 26877 11754 26911
rect 11897 26877 11931 26911
rect 14381 26809 14415 26843
rect 17509 26809 17543 26843
rect 11529 26741 11563 26775
rect 21005 26741 21039 26775
rect 29009 26741 29043 26775
rect 2237 26537 2271 26571
rect 11056 26537 11090 26571
rect 12541 26537 12575 26571
rect 10793 26401 10827 26435
rect 2421 26333 2455 26367
rect 5733 26333 5767 26367
rect 5917 26333 5951 26367
rect 6285 26333 6319 26367
rect 19625 26333 19659 26367
rect 6837 26265 6871 26299
rect 19257 26265 19291 26299
rect 19441 26265 19475 26299
rect 5825 26197 5859 26231
rect 6193 25993 6227 26027
rect 19073 25925 19107 25959
rect 4997 25857 5031 25891
rect 5181 25857 5215 25891
rect 5273 25857 5307 25891
rect 5457 25857 5491 25891
rect 5733 25857 5767 25891
rect 6009 25857 6043 25891
rect 7113 25857 7147 25891
rect 7297 25857 7331 25891
rect 7389 25857 7423 25891
rect 8125 25857 8159 25891
rect 8217 25857 8251 25891
rect 8401 25857 8435 25891
rect 5917 25789 5951 25823
rect 6469 25789 6503 25823
rect 7573 25789 7607 25823
rect 18797 25789 18831 25823
rect 7113 25721 7147 25755
rect 8217 25721 8251 25755
rect 4997 25653 5031 25687
rect 5641 25653 5675 25687
rect 5733 25653 5767 25687
rect 7021 25653 7055 25687
rect 20545 25653 20579 25687
rect 4984 25449 5018 25483
rect 6469 25449 6503 25483
rect 6745 25449 6779 25483
rect 6929 25449 6963 25483
rect 7284 25449 7318 25483
rect 8769 25449 8803 25483
rect 1869 25313 1903 25347
rect 4721 25313 4755 25347
rect 7021 25313 7055 25347
rect 20637 25313 20671 25347
rect 20913 25313 20947 25347
rect 4445 25245 4479 25279
rect 4629 25245 4663 25279
rect 12081 25245 12115 25279
rect 15025 25245 15059 25279
rect 18153 25245 18187 25279
rect 18613 25245 18647 25279
rect 18705 25245 18739 25279
rect 18915 25245 18949 25279
rect 19073 25245 19107 25279
rect 19349 25245 19383 25279
rect 19533 25245 19567 25279
rect 2145 25177 2179 25211
rect 6561 25177 6595 25211
rect 15301 25177 15335 25211
rect 16957 25177 16991 25211
rect 17417 25177 17451 25211
rect 18797 25177 18831 25211
rect 19625 25177 19659 25211
rect 20361 25177 20395 25211
rect 22661 25177 22695 25211
rect 3617 25109 3651 25143
rect 4629 25109 4663 25143
rect 6761 25109 6795 25143
rect 11897 25109 11931 25143
rect 16773 25109 16807 25143
rect 17049 25109 17083 25143
rect 18429 25109 18463 25143
rect 19441 25109 19475 25143
rect 5365 24905 5399 24939
rect 7389 24905 7423 24939
rect 7481 24905 7515 24939
rect 14933 24905 14967 24939
rect 7297 24837 7331 24871
rect 11805 24837 11839 24871
rect 14197 24837 14231 24871
rect 18061 24837 18095 24871
rect 18705 24837 18739 24871
rect 21097 24837 21131 24871
rect 3157 24769 3191 24803
rect 5181 24769 5215 24803
rect 6377 24769 6411 24803
rect 7849 24769 7883 24803
rect 9689 24769 9723 24803
rect 11529 24769 11563 24803
rect 14381 24769 14415 24803
rect 15117 24769 15151 24803
rect 15209 24769 15243 24803
rect 15301 24769 15335 24803
rect 15439 24769 15473 24803
rect 15669 24769 15703 24803
rect 15853 24769 15887 24803
rect 16129 24769 16163 24803
rect 16313 24769 16347 24803
rect 16865 24769 16899 24803
rect 17877 24769 17911 24803
rect 17969 24769 18003 24803
rect 18179 24769 18213 24803
rect 20361 24769 20395 24803
rect 20821 24769 20855 24803
rect 3433 24701 3467 24735
rect 4905 24701 4939 24735
rect 4997 24701 5031 24735
rect 5549 24701 5583 24735
rect 8125 24701 8159 24735
rect 13553 24701 13587 24735
rect 14473 24701 14507 24735
rect 14565 24701 14599 24735
rect 15577 24701 15611 24735
rect 18337 24701 18371 24735
rect 18429 24701 18463 24735
rect 20177 24701 20211 24735
rect 6193 24633 6227 24667
rect 7113 24633 7147 24667
rect 16037 24633 16071 24667
rect 17693 24633 17727 24667
rect 7021 24565 7055 24599
rect 7665 24565 7699 24599
rect 9597 24565 9631 24599
rect 9781 24565 9815 24599
rect 10149 24565 10183 24599
rect 16221 24565 16255 24599
rect 16957 24565 16991 24599
rect 20453 24565 20487 24599
rect 4077 24361 4111 24395
rect 19257 24361 19291 24395
rect 19901 24361 19935 24395
rect 7021 24293 7055 24327
rect 5273 24225 5307 24259
rect 11621 24225 11655 24259
rect 15301 24225 15335 24259
rect 16405 24225 16439 24259
rect 4261 24157 4295 24191
rect 7113 24157 7147 24191
rect 7297 24157 7331 24191
rect 10057 24157 10091 24191
rect 15853 24157 15887 24191
rect 16313 24157 16347 24191
rect 19441 24157 19475 24191
rect 19625 24157 19659 24191
rect 19717 24157 19751 24191
rect 20085 24157 20119 24191
rect 5549 24089 5583 24123
rect 11897 24089 11931 24123
rect 13645 24089 13679 24123
rect 14565 24089 14599 24123
rect 15945 24089 15979 24123
rect 16037 24089 16071 24123
rect 16175 24089 16209 24123
rect 16681 24089 16715 24123
rect 18429 24089 18463 24123
rect 19809 24089 19843 24123
rect 19993 24089 20027 24123
rect 7205 24021 7239 24055
rect 10609 24021 10643 24055
rect 15669 24021 15703 24055
rect 13001 23817 13035 23851
rect 14749 23817 14783 23851
rect 17601 23817 17635 23851
rect 13369 23749 13403 23783
rect 15669 23749 15703 23783
rect 17233 23749 17267 23783
rect 1501 23681 1535 23715
rect 13461 23681 13495 23715
rect 14565 23681 14599 23715
rect 14841 23681 14875 23715
rect 15025 23681 15059 23715
rect 15301 23681 15335 23715
rect 15485 23681 15519 23715
rect 15577 23681 15611 23715
rect 16957 23681 16991 23715
rect 17141 23681 17175 23715
rect 17325 23681 17359 23715
rect 17785 23681 17819 23715
rect 9229 23613 9263 23647
rect 9505 23613 9539 23647
rect 11529 23613 11563 23647
rect 13553 23613 13587 23647
rect 14105 23613 14139 23647
rect 14473 23613 14507 23647
rect 15117 23613 15151 23647
rect 17509 23613 17543 23647
rect 17877 23613 17911 23647
rect 17969 23613 18003 23647
rect 18061 23613 18095 23647
rect 15945 23545 15979 23579
rect 1593 23477 1627 23511
rect 10977 23477 11011 23511
rect 12173 23477 12207 23511
rect 14841 23477 14875 23511
rect 16129 23477 16163 23511
rect 10793 23273 10827 23307
rect 14657 23273 14691 23307
rect 14933 23273 14967 23307
rect 25237 23273 25271 23307
rect 15209 23205 15243 23239
rect 15577 23205 15611 23239
rect 17601 23205 17635 23239
rect 6837 23137 6871 23171
rect 9045 23137 9079 23171
rect 11621 23137 11655 23171
rect 14841 23137 14875 23171
rect 16037 23137 16071 23171
rect 21005 23137 21039 23171
rect 4537 23069 4571 23103
rect 10885 23069 10919 23103
rect 14381 23069 14415 23103
rect 14749 23069 14783 23103
rect 15025 23069 15059 23103
rect 15301 23069 15335 23103
rect 15575 23047 15609 23081
rect 15669 23069 15703 23103
rect 15853 23069 15887 23103
rect 17601 23069 17635 23103
rect 17785 23069 17819 23103
rect 20729 23069 20763 23103
rect 20821 23069 20855 23103
rect 21097 23069 21131 23103
rect 24501 23069 24535 23103
rect 24593 23069 24627 23103
rect 24777 23069 24811 23103
rect 24869 23069 24903 23103
rect 6009 23001 6043 23035
rect 9321 23001 9355 23035
rect 14105 23001 14139 23035
rect 15485 23001 15519 23035
rect 21189 23001 21223 23035
rect 25053 23001 25087 23035
rect 5089 22933 5123 22967
rect 14289 22933 14323 22967
rect 14473 22933 14507 22967
rect 21005 22933 21039 22967
rect 12817 22729 12851 22763
rect 20913 22729 20947 22763
rect 24409 22729 24443 22763
rect 5273 22661 5307 22695
rect 8217 22661 8251 22695
rect 8953 22661 8987 22695
rect 12449 22661 12483 22695
rect 12541 22661 12575 22695
rect 15393 22661 15427 22695
rect 23213 22661 23247 22695
rect 24225 22661 24259 22695
rect 25421 22661 25455 22695
rect 6745 22593 6779 22627
rect 6929 22593 6963 22627
rect 7021 22593 7055 22627
rect 7113 22593 7147 22627
rect 8677 22593 8711 22627
rect 8861 22593 8895 22627
rect 9045 22593 9079 22627
rect 9321 22593 9355 22627
rect 12265 22593 12299 22627
rect 12633 22593 12667 22627
rect 15025 22593 15059 22627
rect 15301 22593 15335 22627
rect 17325 22593 17359 22627
rect 20729 22593 20763 22627
rect 21281 22593 21315 22627
rect 21465 22593 21499 22627
rect 21557 22593 21591 22627
rect 21833 22593 21867 22627
rect 22011 22593 22045 22627
rect 22753 22593 22787 22627
rect 22937 22593 22971 22627
rect 23121 22593 23155 22627
rect 23305 22593 23339 22627
rect 23673 22593 23707 22627
rect 23765 22593 23799 22627
rect 23949 22593 23983 22627
rect 24041 22593 24075 22627
rect 24133 22593 24167 22627
rect 24317 22593 24351 22627
rect 24593 22593 24627 22627
rect 24777 22593 24811 22627
rect 24869 22593 24903 22627
rect 25053 22593 25087 22627
rect 25237 22593 25271 22627
rect 28825 22593 28859 22627
rect 4537 22525 4571 22559
rect 6009 22525 6043 22559
rect 7665 22525 7699 22559
rect 9597 22525 9631 22559
rect 11069 22525 11103 22559
rect 11529 22525 11563 22559
rect 15209 22525 15243 22559
rect 16221 22525 16255 22559
rect 16681 22525 16715 22559
rect 20545 22525 20579 22559
rect 21373 22525 21407 22559
rect 24685 22525 24719 22559
rect 9229 22457 9263 22491
rect 29009 22457 29043 22491
rect 5089 22389 5123 22423
rect 7297 22389 7331 22423
rect 12173 22389 12207 22423
rect 14841 22389 14875 22423
rect 21097 22389 21131 22423
rect 21833 22389 21867 22423
rect 22753 22389 22787 22423
rect 23489 22389 23523 22423
rect 6272 22185 6306 22219
rect 7757 22185 7791 22219
rect 14736 22185 14770 22219
rect 21649 22185 21683 22219
rect 22109 22185 22143 22219
rect 23765 22185 23799 22219
rect 24777 22185 24811 22219
rect 20361 22117 20395 22151
rect 22477 22117 22511 22151
rect 23949 22117 23983 22151
rect 6009 22049 6043 22083
rect 14473 22049 14507 22083
rect 20177 22049 20211 22083
rect 22569 22049 22603 22083
rect 23009 22049 23043 22083
rect 23397 22049 23431 22083
rect 24869 22049 24903 22083
rect 4261 21981 4295 22015
rect 4537 21981 4571 22015
rect 5365 21981 5399 22015
rect 5917 21981 5951 22015
rect 7849 21981 7883 22015
rect 9045 21981 9079 22015
rect 9321 21981 9355 22015
rect 9413 21981 9447 22015
rect 9689 21981 9723 22015
rect 10333 21981 10367 22015
rect 10425 21981 10459 22015
rect 10518 21981 10552 22015
rect 10793 21981 10827 22015
rect 10931 21981 10965 22015
rect 17325 21981 17359 22015
rect 20085 21981 20119 22015
rect 20269 21981 20303 22015
rect 20545 21981 20579 22015
rect 20821 21981 20855 22015
rect 21097 21981 21131 22015
rect 21373 21981 21407 22015
rect 21465 21981 21499 22015
rect 21741 21981 21775 22015
rect 21925 21981 21959 22015
rect 22385 21981 22419 22015
rect 22661 21981 22695 22015
rect 22845 21981 22879 22015
rect 23222 21981 23256 22015
rect 23489 21981 23523 22015
rect 23939 21981 23973 22015
rect 24225 21981 24259 22015
rect 24593 21981 24627 22015
rect 25145 21981 25179 22015
rect 25421 21981 25455 22015
rect 25697 21981 25731 22015
rect 25973 21981 26007 22015
rect 9229 21913 9263 21947
rect 10701 21913 10735 21947
rect 21281 21913 21315 21947
rect 22937 21913 22971 21947
rect 23857 21913 23891 21947
rect 25329 21913 25363 21947
rect 4077 21845 4111 21879
rect 8493 21845 8527 21879
rect 9597 21845 9631 21879
rect 11069 21845 11103 21879
rect 16221 21845 16255 21879
rect 17877 21845 17911 21879
rect 20729 21845 20763 21879
rect 22201 21845 22235 21879
rect 23121 21845 23155 21879
rect 24133 21845 24167 21879
rect 24409 21845 24443 21879
rect 24961 21845 24995 21879
rect 25513 21845 25547 21879
rect 25881 21845 25915 21879
rect 5549 21641 5583 21675
rect 6193 21641 6227 21675
rect 18429 21641 18463 21675
rect 18521 21641 18555 21675
rect 20821 21641 20855 21675
rect 21557 21641 21591 21675
rect 23397 21641 23431 21675
rect 23673 21641 23707 21675
rect 3341 21573 3375 21607
rect 8401 21573 8435 21607
rect 8493 21573 8527 21607
rect 12449 21573 12483 21607
rect 20177 21573 20211 21607
rect 22845 21539 22879 21573
rect 3157 21505 3191 21539
rect 3433 21505 3467 21539
rect 3525 21505 3559 21539
rect 5641 21505 5675 21539
rect 5825 21505 5859 21539
rect 5917 21505 5951 21539
rect 6009 21505 6043 21539
rect 6377 21505 6411 21539
rect 8217 21505 8251 21539
rect 8585 21505 8619 21539
rect 9045 21505 9079 21539
rect 12081 21505 12115 21539
rect 12174 21505 12208 21539
rect 12357 21505 12391 21539
rect 12587 21505 12621 21539
rect 12909 21505 12943 21539
rect 18797 21505 18831 21539
rect 18889 21505 18923 21539
rect 19165 21505 19199 21539
rect 19349 21505 19383 21539
rect 21097 21505 21131 21539
rect 21465 21505 21499 21539
rect 21833 21505 21867 21539
rect 22017 21505 22051 21539
rect 22109 21505 22143 21539
rect 22385 21505 22419 21539
rect 22477 21505 22511 21539
rect 23857 21505 23891 21539
rect 24317 21505 24351 21539
rect 24685 21505 24719 21539
rect 24961 21505 24995 21539
rect 25329 21505 25363 21539
rect 25513 21505 25547 21539
rect 26985 21505 27019 21539
rect 27169 21505 27203 21539
rect 27537 21505 27571 21539
rect 27721 21505 27755 21539
rect 3801 21437 3835 21471
rect 4077 21437 4111 21471
rect 6653 21437 6687 21471
rect 9321 21437 9355 21471
rect 13185 21437 13219 21471
rect 16681 21437 16715 21471
rect 16957 21437 16991 21471
rect 18705 21437 18739 21471
rect 18981 21437 19015 21471
rect 20545 21437 20579 21471
rect 20637 21437 20671 21471
rect 21281 21437 21315 21471
rect 21373 21437 21407 21471
rect 22201 21437 22235 21471
rect 22569 21437 22603 21471
rect 22661 21437 22695 21471
rect 22937 21437 22971 21471
rect 23489 21437 23523 21471
rect 8769 21369 8803 21403
rect 20913 21369 20947 21403
rect 21833 21369 21867 21403
rect 23213 21369 23247 21403
rect 24409 21369 24443 21403
rect 27077 21369 27111 21403
rect 3709 21301 3743 21335
rect 8125 21301 8159 21335
rect 10793 21301 10827 21335
rect 12725 21301 12759 21335
rect 14657 21301 14691 21335
rect 19533 21301 19567 21335
rect 23857 21301 23891 21335
rect 25329 21301 25363 21335
rect 27629 21301 27663 21335
rect 4058 21097 4092 21131
rect 5549 21097 5583 21131
rect 14749 21097 14783 21131
rect 16497 21097 16531 21131
rect 23489 21097 23523 21131
rect 25881 21097 25915 21131
rect 27077 21097 27111 21131
rect 27813 21097 27847 21131
rect 23305 21029 23339 21063
rect 3801 20961 3835 20995
rect 9597 20961 9631 20995
rect 12173 20961 12207 20995
rect 12449 20961 12483 20995
rect 18337 20961 18371 20995
rect 18521 20961 18555 20995
rect 20361 20961 20395 20995
rect 21189 20961 21223 20995
rect 25237 20961 25271 20995
rect 26709 20961 26743 20995
rect 27629 20961 27663 20995
rect 6009 20893 6043 20927
rect 6102 20893 6136 20927
rect 6285 20893 6319 20927
rect 6515 20893 6549 20927
rect 7297 20893 7331 20927
rect 7390 20893 7424 20927
rect 7665 20893 7699 20927
rect 7762 20893 7796 20927
rect 10425 20893 10459 20927
rect 11437 20893 11471 20927
rect 11530 20893 11564 20927
rect 11713 20893 11747 20927
rect 11902 20893 11936 20927
rect 14105 20893 14139 20927
rect 14198 20893 14232 20927
rect 14570 20893 14604 20927
rect 14841 20893 14875 20927
rect 15945 20893 15979 20927
rect 16221 20893 16255 20927
rect 16313 20893 16347 20927
rect 16589 20893 16623 20927
rect 19533 20893 19567 20927
rect 19625 20893 19659 20927
rect 19993 20893 20027 20927
rect 20637 20893 20671 20927
rect 20913 20893 20947 20927
rect 21097 20893 21131 20927
rect 21281 20893 21315 20927
rect 21465 20893 21499 20927
rect 21649 20893 21683 20927
rect 22109 20893 22143 20927
rect 22385 20893 22419 20927
rect 22661 20893 22695 20927
rect 23213 20893 23247 20927
rect 23673 20893 23707 20927
rect 23857 20893 23891 20927
rect 23949 20893 23983 20927
rect 24961 20893 24995 20927
rect 26157 20893 26191 20927
rect 26801 20893 26835 20927
rect 27353 20893 27387 20927
rect 27445 20893 27479 20927
rect 27721 20893 27755 20927
rect 28457 20893 28491 20927
rect 6377 20825 6411 20859
rect 7573 20825 7607 20859
rect 11161 20825 11195 20859
rect 11805 20825 11839 20859
rect 14381 20825 14415 20859
rect 14473 20825 14507 20859
rect 16129 20825 16163 20859
rect 16865 20825 16899 20859
rect 25881 20825 25915 20859
rect 28273 20825 28307 20859
rect 6653 20757 6687 20791
rect 7941 20757 7975 20791
rect 10149 20757 10183 20791
rect 12081 20757 12115 20791
rect 13921 20757 13955 20791
rect 15485 20757 15519 20791
rect 19073 20757 19107 20791
rect 25789 20757 25823 20791
rect 26065 20757 26099 20791
rect 28181 20757 28215 20791
rect 28641 20757 28675 20791
rect 14933 20553 14967 20587
rect 16957 20553 16991 20587
rect 17049 20553 17083 20587
rect 21373 20553 21407 20587
rect 22033 20553 22067 20587
rect 22201 20553 22235 20587
rect 23121 20553 23155 20587
rect 23489 20553 23523 20587
rect 3617 20485 3651 20519
rect 9965 20485 9999 20519
rect 10517 20485 10551 20519
rect 10609 20485 10643 20519
rect 17969 20485 18003 20519
rect 21005 20485 21039 20519
rect 21833 20485 21867 20519
rect 24317 20485 24351 20519
rect 3341 20417 3375 20451
rect 3525 20417 3559 20451
rect 3709 20417 3743 20451
rect 4169 20417 4203 20451
rect 4537 20417 4571 20451
rect 9689 20417 9723 20451
rect 9873 20417 9907 20451
rect 10057 20417 10091 20451
rect 10333 20417 10367 20451
rect 10701 20417 10735 20451
rect 11805 20417 11839 20451
rect 13737 20417 13771 20451
rect 14381 20417 14415 20451
rect 14565 20417 14599 20451
rect 14657 20417 14691 20451
rect 14749 20417 14783 20451
rect 16865 20417 16899 20451
rect 17233 20417 17267 20451
rect 17325 20417 17359 20451
rect 17509 20417 17543 20451
rect 17601 20417 17635 20451
rect 17693 20417 17727 20451
rect 18153 20417 18187 20451
rect 18337 20417 18371 20451
rect 18797 20417 18831 20451
rect 19165 20417 19199 20451
rect 19441 20417 19475 20451
rect 21189 20417 21223 20451
rect 21465 20417 21499 20451
rect 21649 20417 21683 20451
rect 22937 20417 22971 20451
rect 23673 20417 23707 20451
rect 23857 20417 23891 20451
rect 23949 20417 23983 20451
rect 24041 20417 24075 20451
rect 24133 20417 24167 20451
rect 26617 20417 26651 20451
rect 27077 20417 27111 20451
rect 27445 20417 27479 20451
rect 27905 20417 27939 20451
rect 27997 20417 28031 20451
rect 28181 20417 28215 20451
rect 28273 20417 28307 20451
rect 28552 20439 28586 20473
rect 28641 20417 28675 20451
rect 28825 20417 28859 20451
rect 28917 20417 28951 20451
rect 4721 20349 4755 20383
rect 6377 20349 6411 20383
rect 6653 20349 6687 20383
rect 8217 20349 8251 20383
rect 12081 20349 12115 20383
rect 13553 20349 13587 20383
rect 18429 20349 18463 20383
rect 22753 20349 22787 20383
rect 24317 20349 24351 20383
rect 26709 20349 26743 20383
rect 10241 20281 10275 20315
rect 10885 20281 10919 20315
rect 16681 20281 16715 20315
rect 18889 20281 18923 20315
rect 3893 20213 3927 20247
rect 8125 20213 8159 20247
rect 8861 20213 8895 20247
rect 14289 20213 14323 20247
rect 17877 20213 17911 20247
rect 21557 20213 21591 20247
rect 22017 20213 22051 20247
rect 27353 20213 27387 20247
rect 27629 20213 27663 20247
rect 27721 20213 27755 20247
rect 28365 20213 28399 20247
rect 4445 20009 4479 20043
rect 6929 20009 6963 20043
rect 8769 20009 8803 20043
rect 12633 20009 12667 20043
rect 16129 20009 16163 20043
rect 27629 20009 27663 20043
rect 2145 19873 2179 19907
rect 1869 19805 1903 19839
rect 3893 19805 3927 19839
rect 6377 19805 6411 19839
rect 6653 19805 6687 19839
rect 6745 19805 6779 19839
rect 7021 19805 7055 19839
rect 7169 19805 7203 19839
rect 7527 19805 7561 19839
rect 8217 19805 8251 19839
rect 8953 19805 8987 19839
rect 10057 19805 10091 19839
rect 10609 19805 10643 19839
rect 10793 19805 10827 19839
rect 11023 19805 11057 19839
rect 12081 19805 12115 19839
rect 12265 19805 12299 19839
rect 12357 19805 12391 19839
rect 12495 19805 12529 19839
rect 13001 19805 13035 19839
rect 15945 19805 15979 19839
rect 27261 19805 27295 19839
rect 27537 19805 27571 19839
rect 27629 19805 27663 19839
rect 27813 19805 27847 19839
rect 28089 19805 28123 19839
rect 28365 19805 28399 19839
rect 6561 19737 6595 19771
rect 7297 19737 7331 19771
rect 7389 19737 7423 19771
rect 10885 19737 10919 19771
rect 15761 19737 15795 19771
rect 28273 19737 28307 19771
rect 3617 19669 3651 19703
rect 7665 19669 7699 19703
rect 9597 19669 9631 19703
rect 10149 19669 10183 19703
rect 11161 19669 11195 19703
rect 13553 19669 13587 19703
rect 27077 19669 27111 19703
rect 27445 19669 27479 19703
rect 27905 19669 27939 19703
rect 1593 19465 1627 19499
rect 12173 19465 12207 19499
rect 13369 19465 13403 19499
rect 17233 19465 17267 19499
rect 18981 19465 19015 19499
rect 19073 19465 19107 19499
rect 19901 19465 19935 19499
rect 20545 19465 20579 19499
rect 7573 19397 7607 19431
rect 8217 19397 8251 19431
rect 16405 19397 16439 19431
rect 16957 19397 16991 19431
rect 19257 19397 19291 19431
rect 19625 19397 19659 19431
rect 20269 19397 20303 19431
rect 1501 19329 1535 19363
rect 7297 19329 7331 19363
rect 7481 19329 7515 19363
rect 7665 19329 7699 19363
rect 7941 19329 7975 19363
rect 12817 19329 12851 19363
rect 13001 19329 13035 19363
rect 13093 19329 13127 19363
rect 13185 19329 13219 19363
rect 14933 19329 14967 19363
rect 15117 19329 15151 19363
rect 15209 19329 15243 19363
rect 15301 19329 15335 19363
rect 16681 19329 16715 19363
rect 16865 19329 16899 19363
rect 17049 19329 17083 19363
rect 18889 19329 18923 19363
rect 19349 19329 19383 19363
rect 19533 19329 19567 19363
rect 19717 19329 19751 19363
rect 19993 19329 20027 19363
rect 20177 19329 20211 19363
rect 20361 19329 20395 19363
rect 27537 19329 27571 19363
rect 27629 19329 27663 19363
rect 9689 19261 9723 19295
rect 11621 19261 11655 19295
rect 15853 19261 15887 19295
rect 27813 19261 27847 19295
rect 18705 19193 18739 19227
rect 7849 19125 7883 19159
rect 15485 19125 15519 19159
rect 8769 18921 8803 18955
rect 9597 18921 9631 18955
rect 11897 18921 11931 18955
rect 15945 18921 15979 18955
rect 19809 18921 19843 18955
rect 20269 18921 20303 18955
rect 29009 18921 29043 18955
rect 7021 18785 7055 18819
rect 7297 18785 7331 18819
rect 10149 18785 10183 18819
rect 10425 18785 10459 18819
rect 14473 18785 14507 18819
rect 19073 18785 19107 18819
rect 4077 18717 4111 18751
rect 6193 18717 6227 18751
rect 6469 18717 6503 18751
rect 6561 18717 6595 18751
rect 8953 18717 8987 18751
rect 9046 18717 9080 18751
rect 9321 18717 9355 18751
rect 9418 18717 9452 18751
rect 12265 18717 12299 18751
rect 12633 18717 12667 18751
rect 14197 18717 14231 18751
rect 16313 18717 16347 18751
rect 16589 18717 16623 18751
rect 17417 18717 17451 18751
rect 17785 18717 17819 18751
rect 18521 18717 18555 18751
rect 19257 18717 19291 18751
rect 19625 18717 19659 18751
rect 19901 18717 19935 18751
rect 20085 18717 20119 18751
rect 28825 18717 28859 18751
rect 6377 18649 6411 18683
rect 9229 18649 9263 18683
rect 12449 18649 12483 18683
rect 12541 18649 12575 18683
rect 17601 18649 17635 18683
rect 17693 18649 17727 18683
rect 19441 18649 19475 18683
rect 19533 18649 19567 18683
rect 4721 18581 4755 18615
rect 6745 18581 6779 18615
rect 12817 18581 12851 18615
rect 16129 18581 16163 18615
rect 17969 18581 18003 18615
rect 8217 18377 8251 18411
rect 11345 18377 11379 18411
rect 14013 18377 14047 18411
rect 18797 18377 18831 18411
rect 21005 18377 21039 18411
rect 5917 18309 5951 18343
rect 10333 18309 10367 18343
rect 13001 18309 13035 18343
rect 17325 18309 17359 18343
rect 1869 18241 1903 18275
rect 3709 18241 3743 18275
rect 5641 18241 5675 18275
rect 5825 18241 5859 18275
rect 6009 18241 6043 18275
rect 6837 18241 6871 18275
rect 7205 18241 7239 18275
rect 9413 18241 9447 18275
rect 9597 18241 9631 18275
rect 9689 18241 9723 18275
rect 9781 18241 9815 18275
rect 10057 18241 10091 18275
rect 10241 18241 10275 18275
rect 10425 18241 10459 18275
rect 12633 18241 12667 18275
rect 12781 18241 12815 18275
rect 12909 18241 12943 18275
rect 13139 18241 13173 18275
rect 14749 18241 14783 18275
rect 17049 18241 17083 18275
rect 19349 18241 19383 18275
rect 19441 18241 19475 18275
rect 19809 18241 19843 18275
rect 20361 18241 20395 18275
rect 20454 18241 20488 18275
rect 20637 18241 20671 18275
rect 20729 18241 20763 18275
rect 20826 18241 20860 18275
rect 22937 18241 22971 18275
rect 2145 18173 2179 18207
rect 3617 18173 3651 18207
rect 3985 18173 4019 18207
rect 7297 18173 7331 18207
rect 7573 18173 7607 18207
rect 10793 18173 10827 18207
rect 11529 18173 11563 18207
rect 13461 18173 13495 18207
rect 15025 18173 15059 18207
rect 19257 18173 19291 18207
rect 23213 18173 23247 18207
rect 24961 18173 24995 18207
rect 25053 18173 25087 18207
rect 26985 18173 27019 18207
rect 27261 18173 27295 18207
rect 29009 18173 29043 18207
rect 12173 18105 12207 18139
rect 20269 18105 20303 18139
rect 5457 18037 5491 18071
rect 6193 18037 6227 18071
rect 9965 18037 9999 18071
rect 10609 18037 10643 18071
rect 13277 18037 13311 18071
rect 16497 18037 16531 18071
rect 25697 18037 25731 18071
rect 11345 17833 11379 17867
rect 12081 17833 12115 17867
rect 13921 17833 13955 17867
rect 19809 17833 19843 17867
rect 21833 17833 21867 17867
rect 23305 17833 23339 17867
rect 27169 17833 27203 17867
rect 5273 17697 5307 17731
rect 7021 17697 7055 17731
rect 9597 17697 9631 17731
rect 12173 17697 12207 17731
rect 17325 17697 17359 17731
rect 20085 17697 20119 17731
rect 22385 17697 22419 17731
rect 22937 17697 22971 17731
rect 23949 17697 23983 17731
rect 25053 17697 25087 17731
rect 25789 17697 25823 17731
rect 26157 17697 26191 17731
rect 26433 17697 26467 17731
rect 26525 17697 26559 17731
rect 4445 17629 4479 17663
rect 7297 17629 7331 17663
rect 7389 17629 7423 17663
rect 7573 17629 7607 17663
rect 7665 17629 7699 17663
rect 11437 17629 11471 17663
rect 11530 17629 11564 17663
rect 11805 17629 11839 17663
rect 11943 17629 11977 17663
rect 16129 17629 16163 17663
rect 19257 17629 19291 17663
rect 19441 17629 19475 17663
rect 19625 17629 19659 17663
rect 22293 17629 22327 17663
rect 22753 17629 22787 17663
rect 23029 17629 23063 17663
rect 23489 17629 23523 17663
rect 24409 17629 24443 17663
rect 25145 17629 25179 17663
rect 25329 17629 25363 17663
rect 25513 17629 25547 17663
rect 26065 17629 26099 17663
rect 26617 17629 26651 17663
rect 26985 17629 27019 17663
rect 27905 17629 27939 17663
rect 28181 17629 28215 17663
rect 28365 17629 28399 17663
rect 5549 17561 5583 17595
rect 7113 17561 7147 17595
rect 9873 17561 9907 17595
rect 11713 17561 11747 17595
rect 12449 17561 12483 17595
rect 14197 17561 14231 17595
rect 15945 17561 15979 17595
rect 17601 17561 17635 17595
rect 19533 17561 19567 17595
rect 20361 17561 20395 17595
rect 23581 17561 23615 17595
rect 23673 17561 23707 17595
rect 23811 17561 23845 17595
rect 25421 17561 25455 17595
rect 25651 17561 25685 17595
rect 26801 17561 26835 17595
rect 26893 17561 26927 17595
rect 27445 17561 27479 17595
rect 27629 17561 27663 17595
rect 4997 17493 5031 17527
rect 16681 17493 16715 17527
rect 19073 17493 19107 17527
rect 22569 17493 22603 17527
rect 25881 17493 25915 17527
rect 26249 17493 26283 17527
rect 27813 17493 27847 17527
rect 27997 17493 28031 17527
rect 28273 17493 28307 17527
rect 4537 17289 4571 17323
rect 5181 17289 5215 17323
rect 13921 17289 13955 17323
rect 18797 17289 18831 17323
rect 19257 17289 19291 17323
rect 20821 17289 20855 17323
rect 21833 17289 21867 17323
rect 23397 17289 23431 17323
rect 25881 17289 25915 17323
rect 26985 17289 27019 17323
rect 3525 17221 3559 17255
rect 4813 17221 4847 17255
rect 5457 17221 5491 17255
rect 12449 17221 12483 17255
rect 15209 17221 15243 17255
rect 18889 17221 18923 17255
rect 23765 17221 23799 17255
rect 25605 17221 25639 17255
rect 28457 17221 28491 17255
rect 3341 17153 3375 17187
rect 3617 17153 3651 17187
rect 3709 17153 3743 17187
rect 3985 17153 4019 17187
rect 4169 17153 4203 17187
rect 4261 17153 4295 17187
rect 4377 17153 4411 17187
rect 4629 17153 4663 17187
rect 4905 17153 4939 17187
rect 4997 17153 5031 17187
rect 5273 17153 5307 17187
rect 5549 17153 5583 17187
rect 5641 17153 5675 17187
rect 9597 17153 9631 17187
rect 12173 17153 12207 17187
rect 14013 17153 14047 17187
rect 15025 17153 15059 17187
rect 15301 17153 15335 17187
rect 15393 17153 15427 17187
rect 16957 17153 16991 17187
rect 17049 17153 17083 17187
rect 17141 17153 17175 17187
rect 17325 17153 17359 17187
rect 17601 17153 17635 17187
rect 18153 17153 18187 17187
rect 18245 17153 18279 17187
rect 18429 17153 18463 17187
rect 18521 17153 18555 17187
rect 18613 17153 18647 17187
rect 19073 17153 19107 17187
rect 21005 17153 21039 17187
rect 21281 17153 21315 17187
rect 22201 17153 22235 17187
rect 22293 17153 22327 17187
rect 22845 17153 22879 17187
rect 23489 17153 23523 17187
rect 25421 17153 25455 17187
rect 26065 17153 26099 17187
rect 26249 17153 26283 17187
rect 26341 17153 26375 17187
rect 26433 17153 26467 17187
rect 27169 17153 27203 17187
rect 27445 17153 27479 17187
rect 27629 17153 27663 17187
rect 27905 17153 27939 17187
rect 28273 17153 28307 17187
rect 9873 17085 9907 17119
rect 16681 17085 16715 17119
rect 21373 17085 21407 17119
rect 22477 17085 22511 17119
rect 23121 17085 23155 17119
rect 26525 17085 26559 17119
rect 27353 17085 27387 17119
rect 28089 17085 28123 17119
rect 28181 17085 28215 17119
rect 11345 17017 11379 17051
rect 15577 17017 15611 17051
rect 21649 17017 21683 17051
rect 25237 17017 25271 17051
rect 26801 17017 26835 17051
rect 27261 17017 27295 17051
rect 27721 17017 27755 17051
rect 3893 16949 3927 16983
rect 5825 16949 5859 16983
rect 14657 16949 14691 16983
rect 23121 16949 23155 16983
rect 25789 16949 25823 16983
rect 26525 16949 26559 16983
rect 28641 16949 28675 16983
rect 6285 16745 6319 16779
rect 14657 16745 14691 16779
rect 22017 16745 22051 16779
rect 22385 16745 22419 16779
rect 22753 16745 22787 16779
rect 23121 16745 23155 16779
rect 23765 16745 23799 16779
rect 24409 16745 24443 16779
rect 26157 16745 26191 16779
rect 27077 16745 27111 16779
rect 27813 16745 27847 16779
rect 28273 16745 28307 16779
rect 23305 16677 23339 16711
rect 23673 16677 23707 16711
rect 3157 16609 3191 16643
rect 3801 16609 3835 16643
rect 10701 16609 10735 16643
rect 22845 16609 22879 16643
rect 23857 16609 23891 16643
rect 1409 16541 1443 16575
rect 4997 16541 5031 16575
rect 5181 16541 5215 16575
rect 5273 16541 5307 16575
rect 5365 16541 5399 16575
rect 5733 16541 5767 16575
rect 9873 16541 9907 16575
rect 10241 16541 10275 16575
rect 14105 16541 14139 16575
rect 14473 16541 14507 16575
rect 15117 16541 15151 16575
rect 15209 16541 15243 16575
rect 15301 16541 15335 16575
rect 15485 16541 15519 16575
rect 22201 16541 22235 16575
rect 22477 16541 22511 16575
rect 22753 16541 22787 16575
rect 23213 16541 23247 16575
rect 23489 16541 23523 16575
rect 23581 16541 23615 16575
rect 24593 16541 24627 16575
rect 24869 16541 24903 16575
rect 24961 16541 24995 16575
rect 25513 16541 25547 16575
rect 25697 16541 25731 16575
rect 26341 16541 26375 16575
rect 26617 16541 26651 16575
rect 27445 16541 27479 16575
rect 27629 16541 27663 16575
rect 27721 16541 27755 16575
rect 28085 16535 28119 16569
rect 28181 16551 28215 16585
rect 28373 16541 28407 16575
rect 1685 16473 1719 16507
rect 10057 16473 10091 16507
rect 10149 16473 10183 16507
rect 11253 16473 11287 16507
rect 14289 16473 14323 16507
rect 14381 16473 14415 16507
rect 25053 16473 25087 16507
rect 25605 16473 25639 16507
rect 26709 16473 26743 16507
rect 26893 16473 26927 16507
rect 27813 16473 27847 16507
rect 4445 16405 4479 16439
rect 5549 16405 5583 16439
rect 10425 16405 10459 16439
rect 14841 16405 14875 16439
rect 23213 16405 23247 16439
rect 24777 16405 24811 16439
rect 26525 16405 26559 16439
rect 27261 16405 27295 16439
rect 27997 16405 28031 16439
rect 1409 16201 1443 16235
rect 4997 16201 5031 16235
rect 6193 16201 6227 16235
rect 7665 16201 7699 16235
rect 2789 16133 2823 16167
rect 6653 16133 6687 16167
rect 7297 16133 7331 16167
rect 7389 16133 7423 16167
rect 9321 16133 9355 16167
rect 12173 16133 12207 16167
rect 13277 16133 13311 16167
rect 16037 16133 16071 16167
rect 23305 16133 23339 16167
rect 1593 16065 1627 16099
rect 5549 16065 5583 16099
rect 6377 16065 6411 16099
rect 6470 16065 6504 16099
rect 6745 16065 6779 16099
rect 6842 16065 6876 16099
rect 7113 16065 7147 16099
rect 7481 16065 7515 16099
rect 7941 16065 7975 16099
rect 9873 16065 9907 16099
rect 10057 16065 10091 16099
rect 10149 16065 10183 16099
rect 10241 16065 10275 16099
rect 13001 16065 13035 16099
rect 13185 16065 13219 16099
rect 13369 16065 13403 16099
rect 15669 16065 15703 16099
rect 15761 16065 15795 16099
rect 15945 16065 15979 16099
rect 16129 16065 16163 16099
rect 23489 16065 23523 16099
rect 25697 16065 25731 16099
rect 25881 16065 25915 16099
rect 2513 15997 2547 16031
rect 4445 15997 4479 16031
rect 8217 15997 8251 16031
rect 8677 15997 8711 16031
rect 10517 15997 10551 16031
rect 11529 15997 11563 16031
rect 15117 15997 15151 16031
rect 7021 15929 7055 15963
rect 23673 15929 23707 15963
rect 4261 15861 4295 15895
rect 10425 15861 10459 15895
rect 11161 15861 11195 15895
rect 13553 15861 13587 15895
rect 16313 15861 16347 15895
rect 25789 15861 25823 15895
rect 3617 15657 3651 15691
rect 6009 15657 6043 15691
rect 8401 15657 8435 15691
rect 9492 15657 9526 15691
rect 10977 15657 11011 15691
rect 16129 15657 16163 15691
rect 23581 15657 23615 15691
rect 26249 15657 26283 15691
rect 26985 15657 27019 15691
rect 13921 15589 13955 15623
rect 18797 15589 18831 15623
rect 23213 15589 23247 15623
rect 26433 15589 26467 15623
rect 26525 15589 26559 15623
rect 1869 15521 1903 15555
rect 2145 15521 2179 15555
rect 6929 15521 6963 15555
rect 12633 15521 12667 15555
rect 14657 15521 14691 15555
rect 16497 15521 16531 15555
rect 18705 15521 18739 15555
rect 23765 15521 23799 15555
rect 24041 15521 24075 15555
rect 27169 15521 27203 15555
rect 4261 15453 4295 15487
rect 6653 15453 6687 15487
rect 9229 15453 9263 15487
rect 11897 15453 11931 15487
rect 12173 15453 12207 15487
rect 12265 15453 12299 15487
rect 13369 15453 13403 15487
rect 14381 15453 14415 15487
rect 18429 15453 18463 15487
rect 19625 15453 19659 15487
rect 19717 15453 19751 15487
rect 19901 15453 19935 15487
rect 19993 15453 20027 15487
rect 20177 15453 20211 15487
rect 23213 15453 23247 15487
rect 23397 15453 23431 15487
rect 23857 15453 23891 15487
rect 23949 15453 23983 15487
rect 26525 15453 26559 15487
rect 26801 15453 26835 15487
rect 26893 15453 26927 15487
rect 27261 15453 27295 15487
rect 27445 15453 27479 15487
rect 4537 15385 4571 15419
rect 12081 15385 12115 15419
rect 16773 15385 16807 15419
rect 19257 15385 19291 15419
rect 19441 15385 19475 15419
rect 26065 15385 26099 15419
rect 12449 15317 12483 15351
rect 13185 15317 13219 15351
rect 18245 15317 18279 15351
rect 19809 15317 19843 15351
rect 20085 15317 20119 15351
rect 26265 15317 26299 15351
rect 26709 15317 26743 15351
rect 27169 15317 27203 15351
rect 27353 15317 27387 15351
rect 5825 15113 5859 15147
rect 10977 15113 11011 15147
rect 13921 15113 13955 15147
rect 8769 15045 8803 15079
rect 9505 15045 9539 15079
rect 11713 15045 11747 15079
rect 11805 15045 11839 15079
rect 12449 15045 12483 15079
rect 16681 15045 16715 15079
rect 18245 15045 18279 15079
rect 19073 15045 19107 15079
rect 24041 15045 24075 15079
rect 25007 15045 25041 15079
rect 26525 15045 26559 15079
rect 27261 15045 27295 15079
rect 27721 15045 27755 15079
rect 6561 14977 6595 15011
rect 8401 14977 8435 15011
rect 8494 14977 8528 15011
rect 8677 14977 8711 15011
rect 8907 14977 8941 15011
rect 11529 14977 11563 15011
rect 11921 14977 11955 15011
rect 16313 14977 16347 15011
rect 17693 14977 17727 15011
rect 19441 14977 19475 15011
rect 19625 14977 19659 15011
rect 19717 14977 19751 15011
rect 19901 14977 19935 15011
rect 22109 14977 22143 15011
rect 22937 14977 22971 15011
rect 23305 14977 23339 15011
rect 23765 14977 23799 15011
rect 24685 14977 24719 15011
rect 24777 14977 24811 15011
rect 24869 14977 24903 15011
rect 25145 14977 25179 15011
rect 26065 14977 26099 15011
rect 26157 14977 26191 15011
rect 26433 14977 26467 15011
rect 27169 14977 27203 15011
rect 27353 14977 27387 15011
rect 27471 14977 27505 15011
rect 27905 14977 27939 15011
rect 27997 14977 28031 15011
rect 4077 14909 4111 14943
rect 4353 14909 4387 14943
rect 6837 14909 6871 14943
rect 9229 14909 9263 14943
rect 12173 14909 12207 14943
rect 14473 14909 14507 14943
rect 14749 14909 14783 14943
rect 17417 14909 17451 14943
rect 20177 14909 20211 14943
rect 21649 14909 21683 14943
rect 22293 14909 22327 14943
rect 25513 14909 25547 14943
rect 27629 14909 27663 14943
rect 9045 14841 9079 14875
rect 12081 14841 12115 14875
rect 17969 14841 18003 14875
rect 27721 14841 27755 14875
rect 8309 14773 8343 14807
rect 16221 14773 16255 14807
rect 16405 14773 16439 14807
rect 18153 14773 18187 14807
rect 19257 14773 19291 14807
rect 24501 14773 24535 14807
rect 26985 14773 27019 14807
rect 7665 14569 7699 14603
rect 13369 14569 13403 14603
rect 16037 14569 16071 14603
rect 16221 14569 16255 14603
rect 18797 14569 18831 14603
rect 20085 14569 20119 14603
rect 20729 14569 20763 14603
rect 23121 14569 23155 14603
rect 23581 14569 23615 14603
rect 24758 14569 24792 14603
rect 20637 14501 20671 14535
rect 22293 14501 22327 14535
rect 8125 14433 8159 14467
rect 11621 14433 11655 14467
rect 11897 14433 11931 14467
rect 14473 14433 14507 14467
rect 15117 14433 15151 14467
rect 16405 14433 16439 14467
rect 19901 14433 19935 14467
rect 22753 14433 22787 14467
rect 24501 14433 24535 14467
rect 26801 14433 26835 14467
rect 27077 14433 27111 14467
rect 28825 14433 28859 14467
rect 7113 14365 7147 14399
rect 7481 14365 7515 14399
rect 10425 14365 10459 14399
rect 10573 14365 10607 14399
rect 10793 14365 10827 14399
rect 10890 14365 10924 14399
rect 14197 14365 14231 14399
rect 15761 14365 15795 14399
rect 16589 14365 16623 14399
rect 18521 14365 18555 14399
rect 18613 14365 18647 14399
rect 18889 14365 18923 14399
rect 19441 14365 19475 14399
rect 19743 14365 19777 14399
rect 20361 14365 20395 14399
rect 20453 14365 20487 14399
rect 20913 14365 20947 14399
rect 21373 14365 21407 14399
rect 21557 14365 21591 14399
rect 21649 14365 21683 14399
rect 21742 14365 21776 14399
rect 22155 14365 22189 14399
rect 22385 14365 22419 14399
rect 22569 14365 22603 14399
rect 22661 14365 22695 14399
rect 22937 14365 22971 14399
rect 23489 14365 23523 14399
rect 7297 14297 7331 14331
rect 7389 14297 7423 14331
rect 10701 14297 10735 14331
rect 19533 14297 19567 14331
rect 19625 14297 19659 14331
rect 19993 14297 20027 14331
rect 21465 14297 21499 14331
rect 21925 14297 21959 14331
rect 22017 14297 22051 14331
rect 26525 14297 26559 14331
rect 8677 14229 8711 14263
rect 11069 14229 11103 14263
rect 15669 14229 15703 14263
rect 16773 14229 16807 14263
rect 18337 14229 18371 14263
rect 19257 14229 19291 14263
rect 23949 14229 23983 14263
rect 6377 14025 6411 14059
rect 20545 14025 20579 14059
rect 21557 14025 21591 14059
rect 23673 14025 23707 14059
rect 15209 13957 15243 13991
rect 20085 13957 20119 13991
rect 1593 13889 1627 13923
rect 3617 13889 3651 13923
rect 6561 13889 6595 13923
rect 6745 13889 6779 13923
rect 9873 13889 9907 13923
rect 10057 13889 10091 13923
rect 10149 13889 10183 13923
rect 10241 13889 10275 13923
rect 14105 13889 14139 13923
rect 14197 13889 14231 13923
rect 14473 13889 14507 13923
rect 14933 13889 14967 13923
rect 15117 13889 15151 13923
rect 15301 13889 15335 13923
rect 18613 13889 18647 13923
rect 18705 13889 18739 13923
rect 18889 13889 18923 13923
rect 18981 13889 19015 13923
rect 19073 13889 19107 13923
rect 19257 13889 19291 13923
rect 19349 13889 19383 13923
rect 19533 13889 19567 13923
rect 19625 13889 19659 13923
rect 19717 13889 19751 13923
rect 19901 13889 19935 13923
rect 20177 13889 20211 13923
rect 22661 13889 22695 13923
rect 23489 13889 23523 13923
rect 24501 13889 24535 13923
rect 28181 13889 28215 13923
rect 1869 13821 1903 13855
rect 6653 13821 6687 13855
rect 6837 13821 6871 13855
rect 10793 13821 10827 13855
rect 11345 13821 11379 13855
rect 13921 13821 13955 13855
rect 14381 13821 14415 13855
rect 20269 13821 20303 13855
rect 21097 13821 21131 13855
rect 24041 13821 24075 13855
rect 24133 13821 24167 13855
rect 24317 13821 24351 13855
rect 24777 13821 24811 13855
rect 28365 13821 28399 13855
rect 15485 13753 15519 13787
rect 21465 13753 21499 13787
rect 10425 13685 10459 13719
rect 18429 13685 18463 13719
rect 20177 13685 20211 13719
rect 26249 13685 26283 13719
rect 2237 13481 2271 13515
rect 6285 13481 6319 13515
rect 8493 13481 8527 13515
rect 18797 13481 18831 13515
rect 19533 13481 19567 13515
rect 23305 13481 23339 13515
rect 25789 13481 25823 13515
rect 29009 13481 29043 13515
rect 2605 13413 2639 13447
rect 12081 13413 12115 13447
rect 15301 13413 15335 13447
rect 15853 13413 15887 13447
rect 3249 13345 3283 13379
rect 17325 13345 17359 13379
rect 19349 13345 19383 13379
rect 25237 13345 25271 13379
rect 2421 13277 2455 13311
rect 2973 13277 3007 13311
rect 3433 13277 3467 13311
rect 3617 13277 3651 13311
rect 6193 13277 6227 13311
rect 6561 13277 6595 13311
rect 7389 13277 7423 13311
rect 7573 13277 7607 13311
rect 8125 13277 8159 13311
rect 8401 13277 8435 13311
rect 8953 13277 8987 13311
rect 9137 13277 9171 13311
rect 9689 13277 9723 13311
rect 10425 13277 10459 13311
rect 10518 13277 10552 13311
rect 10793 13277 10827 13311
rect 10890 13277 10924 13311
rect 11529 13277 11563 13311
rect 11897 13277 11931 13311
rect 15577 13277 15611 13311
rect 15761 13277 15795 13311
rect 16313 13277 16347 13311
rect 16957 13277 16991 13311
rect 17141 13277 17175 13311
rect 18797 13277 18831 13311
rect 18981 13277 19015 13311
rect 19257 13277 19291 13311
rect 19533 13277 19567 13311
rect 21741 13277 21775 13311
rect 21925 13277 21959 13311
rect 22937 13277 22971 13311
rect 23305 13277 23339 13311
rect 28825 13277 28859 13311
rect 7849 13209 7883 13243
rect 10701 13209 10735 13243
rect 11713 13209 11747 13243
rect 11805 13209 11839 13243
rect 16129 13209 16163 13243
rect 3065 13141 3099 13175
rect 3525 13141 3559 13175
rect 7113 13141 7147 13175
rect 9137 13141 9171 13175
rect 11069 13141 11103 13175
rect 16865 13141 16899 13175
rect 19717 13141 19751 13175
rect 21833 13141 21867 13175
rect 10977 12937 11011 12971
rect 12173 12937 12207 12971
rect 14657 12937 14691 12971
rect 17233 12937 17267 12971
rect 21189 12937 21223 12971
rect 5365 12869 5399 12903
rect 5917 12869 5951 12903
rect 9505 12869 9539 12903
rect 14013 12869 14047 12903
rect 14289 12869 14323 12903
rect 15025 12869 15059 12903
rect 18337 12869 18371 12903
rect 22017 12869 22051 12903
rect 1777 12801 1811 12835
rect 3893 12801 3927 12835
rect 4077 12801 4111 12835
rect 4629 12801 4663 12835
rect 5641 12801 5675 12835
rect 5825 12801 5859 12835
rect 6009 12801 6043 12835
rect 7021 12801 7055 12835
rect 7297 12801 7331 12835
rect 7573 12801 7607 12835
rect 12265 12801 12299 12835
rect 12449 12801 12483 12835
rect 12541 12801 12575 12835
rect 12633 12801 12667 12835
rect 13461 12801 13495 12835
rect 14105 12801 14139 12835
rect 14381 12801 14415 12835
rect 14473 12801 14507 12835
rect 16681 12801 16715 12835
rect 16865 12801 16899 12835
rect 16957 12801 16991 12835
rect 17049 12801 17083 12835
rect 21465 12801 21499 12835
rect 21557 12801 21591 12835
rect 23029 12801 23063 12835
rect 23213 12801 23247 12835
rect 2053 12733 2087 12767
rect 3801 12733 3835 12767
rect 7205 12733 7239 12767
rect 7849 12733 7883 12767
rect 9229 12733 9263 12767
rect 11529 12733 11563 12767
rect 14749 12733 14783 12767
rect 16497 12733 16531 12767
rect 18061 12733 18095 12767
rect 20085 12733 20119 12767
rect 21373 12733 21407 12767
rect 22753 12733 22787 12767
rect 4261 12597 4295 12631
rect 6193 12597 6227 12631
rect 12817 12597 12851 12631
rect 23029 12597 23063 12631
rect 23397 12597 23431 12631
rect 2697 12393 2731 12427
rect 6929 12393 6963 12427
rect 7941 12393 7975 12427
rect 10977 12393 11011 12427
rect 15393 12325 15427 12359
rect 4537 12257 4571 12291
rect 5181 12257 5215 12291
rect 5457 12257 5491 12291
rect 7389 12257 7423 12291
rect 7573 12257 7607 12291
rect 9229 12257 9263 12291
rect 11805 12257 11839 12291
rect 12173 12257 12207 12291
rect 12449 12257 12483 12291
rect 16773 12257 16807 12291
rect 23029 12257 23063 12291
rect 2881 12189 2915 12223
rect 2973 12189 3007 12223
rect 3065 12189 3099 12223
rect 3203 12189 3237 12223
rect 3341 12189 3375 12223
rect 3433 12189 3467 12223
rect 3617 12189 3651 12223
rect 4445 12189 4479 12223
rect 4629 12189 4663 12223
rect 4721 12189 4755 12223
rect 7205 12189 7239 12223
rect 7297 12189 7331 12223
rect 7757 12189 7791 12223
rect 14105 12189 14139 12223
rect 14749 12189 14783 12223
rect 14841 12189 14875 12223
rect 15025 12189 15059 12223
rect 15209 12189 15243 12223
rect 16129 12189 16163 12223
rect 16681 12189 16715 12223
rect 19993 12189 20027 12223
rect 22569 12189 22603 12223
rect 22937 12189 22971 12223
rect 24041 12189 24075 12223
rect 9505 12121 9539 12155
rect 11069 12121 11103 12155
rect 15117 12121 15151 12155
rect 23397 12121 23431 12155
rect 23765 12121 23799 12155
rect 3525 12053 3559 12087
rect 4261 12053 4295 12087
rect 7021 12053 7055 12087
rect 13921 12053 13955 12087
rect 16037 12053 16071 12087
rect 19809 12053 19843 12087
rect 23857 12053 23891 12087
rect 4077 11849 4111 11883
rect 7021 11849 7055 11883
rect 13829 11849 13863 11883
rect 19993 11849 20027 11883
rect 23765 11849 23799 11883
rect 4905 11781 4939 11815
rect 6469 11781 6503 11815
rect 10885 11781 10919 11815
rect 12357 11781 12391 11815
rect 13921 11781 13955 11815
rect 16221 11781 16255 11815
rect 1409 11713 1443 11747
rect 1777 11713 1811 11747
rect 2237 11713 2271 11747
rect 4261 11713 4295 11747
rect 6929 11713 6963 11747
rect 7573 11713 7607 11747
rect 10471 11713 10505 11747
rect 10609 11713 10643 11747
rect 12081 11713 12115 11747
rect 14105 11713 14139 11747
rect 15945 11713 15979 11747
rect 16129 11713 16163 11747
rect 16313 11713 16347 11747
rect 18521 11713 18555 11747
rect 19349 11713 19383 11747
rect 19809 11713 19843 11747
rect 20269 11713 20303 11747
rect 20545 11713 20579 11747
rect 21833 11713 21867 11747
rect 22569 11713 22603 11747
rect 22845 11713 22879 11747
rect 23489 11713 23523 11747
rect 23949 11713 23983 11747
rect 24225 11713 24259 11747
rect 25697 11713 25731 11747
rect 2329 11645 2363 11679
rect 2605 11645 2639 11679
rect 5641 11645 5675 11679
rect 8677 11645 8711 11679
rect 9045 11645 9079 11679
rect 17049 11645 17083 11679
rect 23029 11645 23063 11679
rect 23581 11645 23615 11679
rect 25605 11645 25639 11679
rect 6469 11577 6503 11611
rect 18429 11577 18463 11611
rect 4813 11509 4847 11543
rect 7205 11509 7239 11543
rect 8217 11509 8251 11543
rect 14289 11509 14323 11543
rect 16497 11509 16531 11543
rect 17601 11509 17635 11543
rect 24133 11509 24167 11543
rect 24409 11509 24443 11543
rect 26065 11509 26099 11543
rect 2132 11305 2166 11339
rect 4353 11305 4387 11339
rect 5720 11305 5754 11339
rect 7849 11305 7883 11339
rect 18061 11305 18095 11339
rect 20250 11305 20284 11339
rect 22109 11305 22143 11339
rect 26709 11305 26743 11339
rect 3617 11237 3651 11271
rect 7205 11237 7239 11271
rect 16221 11237 16255 11271
rect 22477 11237 22511 11271
rect 24685 11237 24719 11271
rect 1869 11169 1903 11203
rect 5457 11169 5491 11203
rect 16313 11169 16347 11203
rect 18889 11169 18923 11203
rect 19993 11169 20027 11203
rect 26893 11169 26927 11203
rect 3801 11101 3835 11135
rect 3985 11101 4019 11135
rect 4169 11101 4203 11135
rect 4537 11101 4571 11135
rect 7297 11101 7331 11135
rect 7481 11101 7515 11135
rect 7665 11101 7699 11135
rect 9965 11101 9999 11135
rect 15669 11101 15703 11135
rect 16037 11101 16071 11135
rect 18521 11101 18555 11135
rect 18705 11101 18739 11135
rect 19441 11101 19475 11135
rect 19717 11101 19751 11135
rect 22133 11101 22167 11135
rect 22293 11101 22327 11135
rect 22385 11101 22419 11135
rect 22661 11101 22695 11135
rect 23397 11101 23431 11135
rect 24961 11101 24995 11135
rect 28733 11101 28767 11135
rect 4077 11033 4111 11067
rect 7573 11033 7607 11067
rect 10701 11033 10735 11067
rect 15853 11033 15887 11067
rect 15945 11033 15979 11067
rect 16589 11033 16623 11067
rect 22017 11033 22051 11067
rect 23121 11033 23155 11067
rect 24041 11033 24075 11067
rect 24409 11033 24443 11067
rect 25237 11033 25271 11067
rect 29101 11033 29135 11067
rect 5089 10965 5123 10999
rect 24869 10965 24903 10999
rect 27537 10965 27571 10999
rect 5181 10761 5215 10795
rect 5917 10761 5951 10795
rect 6009 10761 6043 10795
rect 6837 10761 6871 10795
rect 9689 10761 9723 10795
rect 14473 10761 14507 10795
rect 14565 10761 14599 10795
rect 17877 10761 17911 10795
rect 19993 10761 20027 10795
rect 21465 10761 21499 10795
rect 22753 10761 22787 10795
rect 25421 10761 25455 10795
rect 26157 10761 26191 10795
rect 3985 10693 4019 10727
rect 4813 10693 4847 10727
rect 4905 10693 4939 10727
rect 5457 10693 5491 10727
rect 6377 10693 6411 10727
rect 10515 10693 10549 10727
rect 17141 10693 17175 10727
rect 17233 10693 17267 10727
rect 23121 10693 23155 10727
rect 26065 10693 26099 10727
rect 3801 10625 3835 10659
rect 4077 10625 4111 10659
rect 4169 10625 4203 10659
rect 4629 10625 4663 10659
rect 4997 10625 5031 10659
rect 6653 10625 6687 10659
rect 9873 10625 9907 10659
rect 9965 10625 9999 10659
rect 10149 10625 10183 10659
rect 10241 10625 10275 10659
rect 10351 10625 10385 10659
rect 13737 10625 13771 10659
rect 14381 10625 14415 10659
rect 16313 10625 16347 10659
rect 16497 10625 16531 10659
rect 16865 10625 16899 10659
rect 17013 10625 17047 10659
rect 17330 10625 17364 10659
rect 17874 10625 17908 10659
rect 18245 10625 18279 10659
rect 18337 10625 18371 10659
rect 18613 10625 18647 10659
rect 18805 10625 18839 10659
rect 19165 10625 19199 10659
rect 19257 10625 19291 10659
rect 20177 10625 20211 10659
rect 20637 10625 20671 10659
rect 20913 10625 20947 10659
rect 22109 10625 22143 10659
rect 22569 10625 22603 10659
rect 22845 10625 22879 10659
rect 25697 10625 25731 10659
rect 26341 10625 26375 10659
rect 26433 10625 26467 10659
rect 26525 10625 26559 10659
rect 26709 10625 26743 10659
rect 26801 10625 26835 10659
rect 6193 10557 6227 10591
rect 6469 10557 6503 10591
rect 13829 10557 13863 10591
rect 13921 10557 13955 10591
rect 14013 10557 14047 10591
rect 16129 10557 16163 10591
rect 19717 10557 19751 10591
rect 22385 10557 22419 10591
rect 24869 10557 24903 10591
rect 25605 10557 25639 10591
rect 25973 10557 26007 10591
rect 5457 10489 5491 10523
rect 14197 10489 14231 10523
rect 17693 10489 17727 10523
rect 4353 10421 4387 10455
rect 6561 10421 6595 10455
rect 10701 10421 10735 10455
rect 13553 10421 13587 10455
rect 14749 10421 14783 10455
rect 17509 10421 17543 10455
rect 18981 10421 19015 10455
rect 19625 10421 19659 10455
rect 22569 10421 22603 10455
rect 4721 10217 4755 10251
rect 10609 10217 10643 10251
rect 12173 10217 12207 10251
rect 13553 10217 13587 10251
rect 13737 10217 13771 10251
rect 20545 10217 20579 10251
rect 22845 10217 22879 10251
rect 23305 10217 23339 10251
rect 25881 10217 25915 10251
rect 20361 10149 20395 10183
rect 9505 10081 9539 10115
rect 9597 10081 9631 10115
rect 10241 10081 10275 10115
rect 11345 10081 11379 10115
rect 16589 10081 16623 10115
rect 19901 10081 19935 10115
rect 20453 10081 20487 10115
rect 23029 10081 23063 10115
rect 4077 10013 4111 10047
rect 9873 10013 9907 10047
rect 10057 10013 10091 10047
rect 10149 10013 10183 10047
rect 10425 10013 10459 10047
rect 10885 10013 10919 10047
rect 11161 10013 11195 10047
rect 11253 10013 11287 10047
rect 11437 10013 11471 10047
rect 11713 10013 11747 10047
rect 12541 10013 12575 10047
rect 12817 10013 12851 10047
rect 13277 10013 13311 10047
rect 14289 10013 14323 10047
rect 15393 10013 15427 10047
rect 15486 10013 15520 10047
rect 15669 10013 15703 10047
rect 15899 10013 15933 10047
rect 18429 10013 18463 10047
rect 19993 10013 20027 10047
rect 22293 10013 22327 10047
rect 22477 10013 22511 10047
rect 23121 10013 23155 10047
rect 26157 10013 26191 10047
rect 9413 9945 9447 9979
rect 13369 9945 13403 9979
rect 15761 9945 15795 9979
rect 16865 9945 16899 9979
rect 22845 9945 22879 9979
rect 25881 9945 25915 9979
rect 9045 9877 9079 9911
rect 10701 9877 10735 9911
rect 11069 9877 11103 9911
rect 12817 9877 12851 9911
rect 13569 9877 13603 9911
rect 14105 9877 14139 9911
rect 16037 9877 16071 9911
rect 18337 9877 18371 9911
rect 19073 9877 19107 9911
rect 22385 9877 22419 9911
rect 26065 9877 26099 9911
rect 3709 9673 3743 9707
rect 9689 9673 9723 9707
rect 10609 9673 10643 9707
rect 17233 9673 17267 9707
rect 17785 9673 17819 9707
rect 18521 9673 18555 9707
rect 5273 9605 5307 9639
rect 6469 9605 6503 9639
rect 7021 9605 7055 9639
rect 10149 9605 10183 9639
rect 10241 9605 10275 9639
rect 10379 9605 10413 9639
rect 10885 9605 10919 9639
rect 11161 9605 11195 9639
rect 13185 9605 13219 9639
rect 13553 9605 13587 9639
rect 27721 9605 27755 9639
rect 1961 9537 1995 9571
rect 4997 9537 5031 9571
rect 5089 9537 5123 9571
rect 5357 9537 5391 9571
rect 5457 9537 5491 9571
rect 6929 9537 6963 9571
rect 8769 9537 8803 9571
rect 9321 9537 9355 9571
rect 9551 9537 9585 9571
rect 10057 9537 10091 9571
rect 10517 9537 10551 9571
rect 10609 9537 10643 9571
rect 10977 9537 11011 9571
rect 11253 9537 11287 9571
rect 11897 9537 11931 9571
rect 12541 9537 12575 9571
rect 13277 9537 13311 9571
rect 16681 9537 16715 9571
rect 16865 9537 16899 9571
rect 16957 9537 16991 9571
rect 17049 9537 17083 9571
rect 17782 9537 17816 9571
rect 18153 9537 18187 9571
rect 18462 9537 18496 9571
rect 26249 9537 26283 9571
rect 26479 9537 26513 9571
rect 27905 9537 27939 9571
rect 27997 9537 28031 9571
rect 28181 9537 28215 9571
rect 28273 9537 28307 9571
rect 2237 9469 2271 9503
rect 4353 9469 4387 9503
rect 8677 9469 8711 9503
rect 8861 9469 8895 9503
rect 8953 9469 8987 9503
rect 9137 9469 9171 9503
rect 9413 9469 9447 9503
rect 9781 9469 9815 9503
rect 10701 9469 10735 9503
rect 15301 9469 15335 9503
rect 18245 9469 18279 9503
rect 18981 9469 19015 9503
rect 26985 9469 27019 9503
rect 6469 9401 6503 9435
rect 8493 9401 8527 9435
rect 9873 9401 9907 9435
rect 10977 9401 11011 9435
rect 27629 9401 27663 9435
rect 5641 9333 5675 9367
rect 7205 9333 7239 9367
rect 17601 9333 17635 9367
rect 18337 9333 18371 9367
rect 18889 9333 18923 9367
rect 26341 9333 26375 9367
rect 2132 9129 2166 9163
rect 13093 9129 13127 9163
rect 22569 9129 22603 9163
rect 23029 9129 23063 9163
rect 27997 9129 28031 9163
rect 4905 9061 4939 9095
rect 5365 9061 5399 9095
rect 1869 8993 1903 9027
rect 3617 8993 3651 9027
rect 5825 8993 5859 9027
rect 6193 8993 6227 9027
rect 9321 8993 9355 9027
rect 11161 8993 11195 9027
rect 11370 8993 11404 9027
rect 14657 8993 14691 9027
rect 22385 8993 22419 9027
rect 22661 8993 22695 9027
rect 26249 8993 26283 9027
rect 4261 8925 4295 8959
rect 5917 8925 5951 8959
rect 6561 8925 6595 8959
rect 8953 8925 8987 8959
rect 10885 8925 10919 8959
rect 11621 8925 11655 8959
rect 11897 8925 11931 8959
rect 13001 8925 13035 8959
rect 13829 8925 13863 8959
rect 17969 8925 18003 8959
rect 18153 8925 18187 8959
rect 18337 8925 18371 8959
rect 19349 8925 19383 8959
rect 22109 8925 22143 8959
rect 22201 8925 22235 8959
rect 22845 8925 22879 8959
rect 25697 8925 25731 8959
rect 26157 8925 26191 8959
rect 28365 8925 28399 8959
rect 5365 8857 5399 8891
rect 11253 8857 11287 8891
rect 13553 8857 13587 8891
rect 18241 8857 18275 8891
rect 19901 8857 19935 8891
rect 22569 8857 22603 8891
rect 25789 8857 25823 8891
rect 25881 8857 25915 8891
rect 26019 8857 26053 8891
rect 26525 8857 26559 8891
rect 28181 8857 28215 8891
rect 28549 8857 28583 8891
rect 6101 8789 6135 8823
rect 7987 8789 8021 8823
rect 10747 8789 10781 8823
rect 11529 8789 11563 8823
rect 13651 8789 13685 8823
rect 13737 8789 13771 8823
rect 15209 8789 15243 8823
rect 18521 8789 18555 8823
rect 21741 8789 21775 8823
rect 25513 8789 25547 8823
rect 5457 8585 5491 8619
rect 5641 8585 5675 8619
rect 13369 8585 13403 8619
rect 20637 8585 20671 8619
rect 26801 8585 26835 8619
rect 4261 8517 4295 8551
rect 4997 8517 5031 8551
rect 7665 8517 7699 8551
rect 8309 8517 8343 8551
rect 9045 8517 9079 8551
rect 9229 8517 9263 8551
rect 13737 8517 13771 8551
rect 15485 8517 15519 8551
rect 23397 8517 23431 8551
rect 27077 8517 27111 8551
rect 27813 8517 27847 8551
rect 2145 8449 2179 8483
rect 3985 8449 4019 8483
rect 4169 8449 4203 8483
rect 4353 8449 4387 8483
rect 5273 8449 5307 8483
rect 6837 8449 6871 8483
rect 7297 8449 7331 8483
rect 13093 8449 13127 8483
rect 16865 8449 16899 8483
rect 17049 8449 17083 8483
rect 17141 8449 17175 8483
rect 17289 8449 17323 8483
rect 17417 8449 17451 8483
rect 17509 8449 17543 8483
rect 17647 8449 17681 8483
rect 18889 8449 18923 8483
rect 21097 8449 21131 8483
rect 22845 8449 22879 8483
rect 23029 8449 23063 8483
rect 23489 8449 23523 8483
rect 23949 8449 23983 8483
rect 24133 8449 24167 8483
rect 26065 8449 26099 8483
rect 26985 8449 27019 8483
rect 27261 8449 27295 8483
rect 27445 8449 27479 8483
rect 2421 8381 2455 8415
rect 5181 8381 5215 8415
rect 5825 8381 5859 8415
rect 5917 8381 5951 8415
rect 6009 8381 6043 8415
rect 6101 8381 6135 8415
rect 6561 8381 6595 8415
rect 6653 8381 6687 8415
rect 6745 8381 6779 8415
rect 8769 8381 8803 8415
rect 8861 8381 8895 8415
rect 9965 8381 9999 8415
rect 13369 8381 13403 8415
rect 13461 8381 13495 8415
rect 16681 8381 16715 8415
rect 19165 8381 19199 8415
rect 23765 8381 23799 8415
rect 25881 8381 25915 8415
rect 26341 8381 26375 8415
rect 3893 8313 3927 8347
rect 4537 8313 4571 8347
rect 8309 8313 8343 8347
rect 13185 8313 13219 8347
rect 23673 8313 23707 8347
rect 23949 8313 23983 8347
rect 26617 8313 26651 8347
rect 5273 8245 5307 8279
rect 6377 8245 6411 8279
rect 17785 8245 17819 8279
rect 20913 8245 20947 8279
rect 23213 8245 23247 8279
rect 23857 8245 23891 8279
rect 26249 8245 26283 8279
rect 5181 8041 5215 8075
rect 5549 8041 5583 8075
rect 6101 8041 6135 8075
rect 13737 8041 13771 8075
rect 22385 8041 22419 8075
rect 23213 8041 23247 8075
rect 25237 8041 25271 8075
rect 27629 8041 27663 8075
rect 6745 7973 6779 8007
rect 27813 7973 27847 8007
rect 1961 7905 1995 7939
rect 5733 7905 5767 7939
rect 6285 7905 6319 7939
rect 20361 7905 20395 7939
rect 24777 7905 24811 7939
rect 26249 7905 26283 7939
rect 27169 7905 27203 7939
rect 27537 7905 27571 7939
rect 1685 7837 1719 7871
rect 3985 7837 4019 7871
rect 4537 7837 4571 7871
rect 4629 7837 4663 7871
rect 4997 7837 5031 7871
rect 5825 7837 5859 7871
rect 5917 7837 5951 7871
rect 6377 7837 6411 7871
rect 7481 7837 7515 7871
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 14565 7837 14599 7871
rect 14749 7837 14783 7871
rect 16405 7837 16439 7871
rect 16589 7837 16623 7871
rect 16865 7837 16899 7871
rect 17049 7837 17083 7871
rect 17417 7837 17451 7871
rect 17509 7837 17543 7871
rect 17785 7837 17819 7871
rect 17933 7837 17967 7871
rect 18061 7837 18095 7871
rect 18153 7837 18187 7871
rect 18250 7837 18284 7871
rect 20085 7837 20119 7871
rect 22017 7837 22051 7871
rect 22293 7837 22327 7871
rect 22569 7837 22603 7871
rect 22891 7837 22925 7871
rect 22983 7837 23017 7871
rect 23127 7837 23161 7871
rect 23305 7837 23339 7871
rect 23673 7837 23707 7871
rect 23765 7837 23799 7871
rect 23857 7837 23891 7871
rect 24041 7837 24075 7871
rect 24409 7837 24443 7871
rect 24593 7837 24627 7871
rect 24869 7837 24903 7871
rect 25053 7837 25087 7871
rect 25789 7837 25823 7871
rect 25973 7837 26007 7871
rect 26525 7837 26559 7871
rect 27261 7837 27295 7871
rect 4813 7769 4847 7803
rect 4905 7769 4939 7803
rect 6101 7769 6135 7803
rect 6745 7769 6779 7803
rect 7297 7769 7331 7803
rect 13553 7769 13587 7803
rect 13769 7769 13803 7803
rect 17233 7769 17267 7803
rect 22201 7769 22235 7803
rect 22661 7769 22695 7803
rect 22753 7769 22787 7803
rect 23397 7769 23431 7803
rect 25881 7769 25915 7803
rect 26091 7769 26125 7803
rect 3433 7701 3467 7735
rect 6561 7701 6595 7735
rect 7205 7701 7239 7735
rect 13921 7701 13955 7735
rect 14473 7701 14507 7735
rect 14657 7701 14691 7735
rect 16773 7701 16807 7735
rect 18429 7701 18463 7735
rect 21833 7701 21867 7735
rect 22293 7701 22327 7735
rect 25605 7701 25639 7735
rect 5641 7497 5675 7531
rect 16957 7497 16991 7531
rect 22569 7497 22603 7531
rect 22937 7497 22971 7531
rect 27169 7497 27203 7531
rect 27629 7497 27663 7531
rect 11529 7429 11563 7463
rect 13001 7429 13035 7463
rect 13829 7429 13863 7463
rect 18337 7429 18371 7463
rect 22477 7429 22511 7463
rect 23765 7429 23799 7463
rect 24133 7429 24167 7463
rect 25237 7429 25271 7463
rect 6009 7361 6043 7395
rect 10333 7361 10367 7395
rect 10609 7361 10643 7395
rect 10885 7361 10919 7395
rect 11805 7361 11839 7395
rect 12265 7361 12299 7395
rect 13185 7361 13219 7395
rect 13369 7361 13403 7395
rect 13553 7361 13587 7395
rect 16773 7361 16807 7395
rect 17049 7361 17083 7395
rect 17141 7361 17175 7395
rect 17289 7361 17323 7395
rect 17417 7361 17451 7395
rect 17509 7361 17543 7395
rect 17601 7361 17635 7395
rect 17877 7361 17911 7395
rect 18061 7361 18095 7395
rect 18245 7361 18279 7395
rect 18429 7361 18463 7395
rect 22753 7361 22787 7395
rect 23029 7361 23063 7395
rect 23857 7361 23891 7395
rect 24041 7361 24075 7395
rect 24225 7361 24259 7395
rect 24501 7361 24535 7395
rect 24685 7361 24719 7395
rect 24961 7361 24995 7395
rect 26985 7361 27019 7395
rect 27261 7361 27295 7395
rect 27445 7361 27479 7395
rect 27537 7361 27571 7395
rect 27721 7361 27755 7395
rect 28733 7361 28767 7395
rect 5825 7293 5859 7327
rect 5917 7293 5951 7327
rect 11069 7293 11103 7327
rect 13461 7293 13495 7327
rect 15577 7293 15611 7327
rect 21925 7293 21959 7327
rect 23213 7293 23247 7327
rect 26709 7293 26743 7327
rect 12081 7225 12115 7259
rect 24501 7225 24535 7259
rect 11897 7157 11931 7191
rect 11989 7157 12023 7191
rect 16773 7157 16807 7191
rect 17141 7157 17175 7191
rect 17877 7157 17911 7191
rect 24409 7157 24443 7191
rect 29009 7157 29043 7191
rect 11161 6953 11195 6987
rect 11345 6953 11379 6987
rect 14473 6953 14507 6987
rect 20808 6953 20842 6987
rect 22293 6953 22327 6987
rect 22740 6953 22774 6987
rect 8033 6885 8067 6919
rect 12173 6885 12207 6919
rect 24225 6885 24259 6919
rect 5365 6817 5399 6851
rect 11989 6817 12023 6851
rect 14565 6817 14599 6851
rect 20545 6817 20579 6851
rect 22477 6817 22511 6851
rect 24501 6817 24535 6851
rect 4537 6749 4571 6783
rect 4721 6749 4755 6783
rect 4905 6749 4939 6783
rect 6009 6749 6043 6783
rect 6193 6749 6227 6783
rect 6377 6749 6411 6783
rect 6837 6749 6871 6783
rect 7021 6749 7055 6783
rect 7205 6749 7239 6783
rect 7481 6749 7515 6783
rect 7665 6749 7699 6783
rect 7849 6749 7883 6783
rect 9965 6749 9999 6783
rect 10057 6749 10091 6783
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 10793 6749 10827 6783
rect 11621 6749 11655 6783
rect 12081 6749 12115 6783
rect 13737 6749 13771 6783
rect 13921 6749 13955 6783
rect 14289 6749 14323 6783
rect 17049 6749 17083 6783
rect 17325 6749 17359 6783
rect 17417 6749 17451 6783
rect 17877 6749 17911 6783
rect 18061 6749 18095 6783
rect 24409 6749 24443 6783
rect 24593 6749 24627 6783
rect 4813 6681 4847 6715
rect 6285 6681 6319 6715
rect 7113 6681 7147 6715
rect 7757 6681 7791 6715
rect 10517 6681 10551 6715
rect 11437 6681 11471 6715
rect 11713 6681 11747 6715
rect 13829 6681 13863 6715
rect 17601 6681 17635 6715
rect 5089 6613 5123 6647
rect 5917 6613 5951 6647
rect 6561 6613 6595 6647
rect 7389 6613 7423 6647
rect 11161 6613 11195 6647
rect 11805 6613 11839 6647
rect 14105 6613 14139 6647
rect 16865 6613 16899 6647
rect 17233 6613 17267 6647
rect 17785 6613 17819 6647
rect 17969 6613 18003 6647
rect 5641 6409 5675 6443
rect 7021 6409 7055 6443
rect 8769 6409 8803 6443
rect 10885 6409 10919 6443
rect 11069 6409 11103 6443
rect 17141 6409 17175 6443
rect 20085 6409 20119 6443
rect 20453 6409 20487 6443
rect 20637 6409 20671 6443
rect 4169 6341 4203 6375
rect 8033 6341 8067 6375
rect 10057 6341 10091 6375
rect 10517 6341 10551 6375
rect 13737 6341 13771 6375
rect 15485 6341 15519 6375
rect 16957 6341 16991 6375
rect 21005 6341 21039 6375
rect 3893 6273 3927 6307
rect 7389 6273 7423 6307
rect 8125 6273 8159 6307
rect 9965 6273 9999 6307
rect 10241 6273 10275 6307
rect 10609 6273 10643 6307
rect 10977 6273 11011 6307
rect 11161 6273 11195 6307
rect 11529 6273 11563 6307
rect 17233 6273 17267 6307
rect 20269 6273 20303 6307
rect 20545 6273 20579 6307
rect 20821 6273 20855 6307
rect 21097 6273 21131 6307
rect 6377 6205 6411 6239
rect 10726 6205 10760 6239
rect 11713 6205 11747 6239
rect 13461 6205 13495 6239
rect 16957 6069 16991 6103
rect 4248 5865 4282 5899
rect 8033 5865 8067 5899
rect 10793 5865 10827 5899
rect 11069 5865 11103 5899
rect 17693 5865 17727 5899
rect 5733 5797 5767 5831
rect 17877 5797 17911 5831
rect 6285 5729 6319 5763
rect 6561 5729 6595 5763
rect 10885 5729 10919 5763
rect 3985 5661 4019 5695
rect 9413 5661 9447 5695
rect 9689 5661 9723 5695
rect 9965 5661 9999 5695
rect 10057 5661 10091 5695
rect 10149 5661 10183 5695
rect 10241 5661 10275 5695
rect 10425 5661 10459 5695
rect 10609 5661 10643 5695
rect 10977 5661 11011 5695
rect 11161 5661 11195 5695
rect 11253 5661 11287 5695
rect 11529 5661 11563 5695
rect 11621 5661 11655 5695
rect 17601 5661 17635 5695
rect 18153 5661 18187 5695
rect 18245 5661 18279 5695
rect 18429 5661 18463 5695
rect 9597 5593 9631 5627
rect 11437 5593 11471 5627
rect 17417 5593 17451 5627
rect 17877 5593 17911 5627
rect 9229 5525 9263 5559
rect 9781 5525 9815 5559
rect 11805 5525 11839 5559
rect 18061 5525 18095 5559
rect 18337 5525 18371 5559
rect 8125 5321 8159 5355
rect 16891 5321 16925 5355
rect 17325 5321 17359 5355
rect 20361 5321 20395 5355
rect 28273 5321 28307 5355
rect 6653 5253 6687 5287
rect 11069 5253 11103 5287
rect 13323 5253 13357 5287
rect 16681 5253 16715 5287
rect 6377 5185 6411 5219
rect 8493 5185 8527 5219
rect 10517 5185 10551 5219
rect 11529 5185 11563 5219
rect 11897 5185 11931 5219
rect 17141 5185 17175 5219
rect 17509 5185 17543 5219
rect 17785 5185 17819 5219
rect 17969 5185 18003 5219
rect 18245 5185 18279 5219
rect 18521 5185 18555 5219
rect 18705 5185 18739 5219
rect 18981 5185 19015 5219
rect 19165 5185 19199 5219
rect 19625 5185 19659 5219
rect 20269 5185 20303 5219
rect 28089 5185 28123 5219
rect 8861 5117 8895 5151
rect 10333 5117 10367 5151
rect 20085 5117 20119 5151
rect 18981 5049 19015 5083
rect 16865 4981 16899 5015
rect 17049 4981 17083 5015
rect 17509 4981 17543 5015
rect 17877 4981 17911 5015
rect 18889 4981 18923 5015
rect 19717 4981 19751 5015
rect 10701 4777 10735 4811
rect 11345 4777 11379 4811
rect 16957 4777 16991 4811
rect 17601 4777 17635 4811
rect 19993 4777 20027 4811
rect 20453 4777 20487 4811
rect 16221 4709 16255 4743
rect 18797 4709 18831 4743
rect 8953 4641 8987 4675
rect 9321 4641 9355 4675
rect 11161 4641 11195 4675
rect 13369 4641 13403 4675
rect 16037 4641 16071 4675
rect 17693 4641 17727 4675
rect 18153 4641 18187 4675
rect 18429 4641 18463 4675
rect 18889 4641 18923 4675
rect 19533 4641 19567 4675
rect 19625 4641 19659 4675
rect 11069 4573 11103 4607
rect 13093 4573 13127 4607
rect 13277 4573 13311 4607
rect 15945 4573 15979 4607
rect 16129 4573 16163 4607
rect 16497 4573 16531 4607
rect 16589 4573 16623 4607
rect 17417 4573 17451 4607
rect 17969 4573 18003 4607
rect 18245 4573 18279 4607
rect 18613 4573 18647 4607
rect 19441 4573 19475 4607
rect 19717 4573 19751 4607
rect 19901 4573 19935 4607
rect 20177 4573 20211 4607
rect 20545 4573 20579 4607
rect 20729 4573 20763 4607
rect 16221 4505 16255 4539
rect 17785 4505 17819 4539
rect 20637 4505 20671 4539
rect 12909 4437 12943 4471
rect 16405 4437 16439 4471
rect 16957 4437 16991 4471
rect 17141 4437 17175 4471
rect 17233 4437 17267 4471
rect 19257 4437 19291 4471
rect 13185 4233 13219 4267
rect 13921 4233 13955 4267
rect 14473 4233 14507 4267
rect 15761 4233 15795 4267
rect 19993 4233 20027 4267
rect 24041 4165 24075 4199
rect 24225 4165 24259 4199
rect 24777 4165 24811 4199
rect 2421 4097 2455 4131
rect 13123 4097 13157 4131
rect 13645 4097 13679 4131
rect 13737 4097 13771 4131
rect 14381 4097 14415 4131
rect 14565 4097 14599 4131
rect 15577 4097 15611 4131
rect 15761 4097 15795 4131
rect 16037 4097 16071 4131
rect 16313 4097 16347 4131
rect 16681 4097 16715 4131
rect 17325 4097 17359 4131
rect 17601 4097 17635 4131
rect 18797 4097 18831 4131
rect 19257 4097 19291 4131
rect 19717 4097 19751 4131
rect 19809 4097 19843 4131
rect 20085 4097 20119 4131
rect 24593 4097 24627 4131
rect 14059 4029 14093 4063
rect 16221 4029 16255 4063
rect 17417 4029 17451 4063
rect 19533 4029 19567 4063
rect 19993 4029 20027 4063
rect 13001 3961 13035 3995
rect 2237 3893 2271 3927
rect 13553 3893 13587 3927
rect 14289 3893 14323 3927
rect 15853 3893 15887 3927
rect 20177 3893 20211 3927
rect 24409 3893 24443 3927
rect 24961 3893 24995 3927
rect 12633 3689 12667 3723
rect 14289 3689 14323 3723
rect 14749 3689 14783 3723
rect 15485 3689 15519 3723
rect 15117 3621 15151 3655
rect 18061 3553 18095 3587
rect 18981 3553 19015 3587
rect 1501 3485 1535 3519
rect 2421 3485 2455 3519
rect 12541 3485 12575 3519
rect 13001 3485 13035 3519
rect 13277 3485 13311 3519
rect 13461 3485 13495 3519
rect 13737 3485 13771 3519
rect 14473 3485 14507 3519
rect 14565 3485 14599 3519
rect 15393 3485 15427 3519
rect 15577 3485 15611 3519
rect 16681 3485 16715 3519
rect 16773 3485 16807 3519
rect 16865 3485 16899 3519
rect 17049 3485 17083 3519
rect 18705 3485 18739 3519
rect 25421 3485 25455 3519
rect 14105 3417 14139 3451
rect 14841 3417 14875 3451
rect 16405 3417 16439 3451
rect 17877 3417 17911 3451
rect 1593 3349 1627 3383
rect 2237 3349 2271 3383
rect 12817 3349 12851 3383
rect 13829 3349 13863 3383
rect 15301 3349 15335 3383
rect 17509 3349 17543 3383
rect 17969 3349 18003 3383
rect 18337 3349 18371 3383
rect 18797 3349 18831 3383
rect 25237 3349 25271 3383
rect 13001 3145 13035 3179
rect 14565 3145 14599 3179
rect 17601 3145 17635 3179
rect 17969 3145 18003 3179
rect 12909 3009 12943 3043
rect 13093 3009 13127 3043
rect 13369 3009 13403 3043
rect 13461 3009 13495 3043
rect 13645 3009 13679 3043
rect 13737 3009 13771 3043
rect 14013 3009 14047 3043
rect 14197 3009 14231 3043
rect 14289 3009 14323 3043
rect 14381 3009 14415 3043
rect 14565 3009 14599 3043
rect 16865 3009 16899 3043
rect 17049 3009 17083 3043
rect 17141 3009 17175 3043
rect 17233 3009 17267 3043
rect 17693 3009 17727 3043
rect 17785 3009 17819 3043
rect 18061 3009 18095 3043
rect 18245 3009 18279 3043
rect 28825 3009 28859 3043
rect 16957 2941 16991 2975
rect 17417 2941 17451 2975
rect 17509 2941 17543 2975
rect 17969 2941 18003 2975
rect 13829 2873 13863 2907
rect 13185 2805 13219 2839
rect 18061 2805 18095 2839
rect 29009 2805 29043 2839
rect 13461 2601 13495 2635
rect 1501 2397 1535 2431
rect 3893 2397 3927 2431
rect 13461 2397 13495 2431
rect 13645 2397 13679 2431
rect 15025 2397 15059 2431
rect 19349 2397 19383 2431
rect 22109 2397 22143 2431
rect 25973 2397 26007 2431
rect 28733 2397 28767 2431
rect 7297 2329 7331 2363
rect 11621 2329 11655 2363
rect 29101 2329 29135 2363
rect 1593 2261 1627 2295
rect 4169 2261 4203 2295
rect 7389 2261 7423 2295
rect 11713 2261 11747 2295
rect 15301 2261 15335 2295
rect 19441 2261 19475 2295
rect 22201 2261 22235 2295
rect 26249 2261 26283 2295
<< metal1 >>
rect 1104 30490 29595 30512
rect 1104 30438 8032 30490
rect 8084 30438 8096 30490
rect 8148 30438 8160 30490
rect 8212 30438 8224 30490
rect 8276 30438 8288 30490
rect 8340 30438 15115 30490
rect 15167 30438 15179 30490
rect 15231 30438 15243 30490
rect 15295 30438 15307 30490
rect 15359 30438 15371 30490
rect 15423 30438 22198 30490
rect 22250 30438 22262 30490
rect 22314 30438 22326 30490
rect 22378 30438 22390 30490
rect 22442 30438 22454 30490
rect 22506 30438 29281 30490
rect 29333 30438 29345 30490
rect 29397 30438 29409 30490
rect 29461 30438 29473 30490
rect 29525 30438 29537 30490
rect 29589 30438 29595 30490
rect 1104 30416 29595 30438
rect 6730 30336 6736 30388
rect 6788 30336 6794 30388
rect 9674 30268 9680 30320
rect 9732 30308 9738 30320
rect 10229 30311 10287 30317
rect 10229 30308 10241 30311
rect 9732 30280 10241 30308
rect 9732 30268 9738 30280
rect 10229 30277 10241 30280
rect 10275 30277 10287 30311
rect 10229 30271 10287 30277
rect 21266 30268 21272 30320
rect 21324 30308 21330 30320
rect 22281 30311 22339 30317
rect 22281 30308 22293 30311
rect 21324 30280 22293 30308
rect 21324 30268 21330 30280
rect 22281 30277 22293 30280
rect 22327 30277 22339 30311
rect 22281 30271 22339 30277
rect 25406 30268 25412 30320
rect 25464 30308 25470 30320
rect 25685 30311 25743 30317
rect 25685 30308 25697 30311
rect 25464 30280 25697 30308
rect 25464 30268 25470 30280
rect 25685 30277 25697 30280
rect 25731 30277 25743 30311
rect 28994 30308 29000 30320
rect 25685 30271 25743 30277
rect 28368 30280 29000 30308
rect 1578 30200 1584 30252
rect 1636 30200 1642 30252
rect 2777 30243 2835 30249
rect 2777 30209 2789 30243
rect 2823 30240 2835 30243
rect 3418 30240 3424 30252
rect 2823 30212 3424 30240
rect 2823 30209 2835 30212
rect 2777 30203 2835 30209
rect 3418 30200 3424 30212
rect 3476 30200 3482 30252
rect 6086 30200 6092 30252
rect 6144 30240 6150 30252
rect 6641 30243 6699 30249
rect 6641 30240 6653 30243
rect 6144 30212 6653 30240
rect 6144 30200 6150 30212
rect 6641 30209 6653 30212
rect 6687 30209 6699 30243
rect 6641 30203 6699 30209
rect 9858 30200 9864 30252
rect 9916 30200 9922 30252
rect 14182 30200 14188 30252
rect 14240 30200 14246 30252
rect 17586 30200 17592 30252
rect 17644 30200 17650 30252
rect 21910 30200 21916 30252
rect 21968 30200 21974 30252
rect 25314 30200 25320 30252
rect 25372 30200 25378 30252
rect 28368 30249 28396 30280
rect 28994 30268 29000 30280
rect 29052 30268 29058 30320
rect 28353 30243 28411 30249
rect 28353 30209 28365 30243
rect 28399 30209 28411 30243
rect 28353 30203 28411 30209
rect 28718 30200 28724 30252
rect 28776 30200 28782 30252
rect 28902 30132 28908 30184
rect 28960 30172 28966 30184
rect 28997 30175 29055 30181
rect 28997 30172 29009 30175
rect 28960 30144 29009 30172
rect 28960 30132 28966 30144
rect 28997 30141 29009 30144
rect 29043 30141 29055 30175
rect 28997 30135 29055 30141
rect 2774 30064 2780 30116
rect 2832 30104 2838 30116
rect 2961 30107 3019 30113
rect 2961 30104 2973 30107
rect 2832 30076 2973 30104
rect 2832 30064 2838 30076
rect 2961 30073 2973 30076
rect 3007 30073 3019 30107
rect 2961 30067 3019 30073
rect 13814 30064 13820 30116
rect 13872 30104 13878 30116
rect 14369 30107 14427 30113
rect 14369 30104 14381 30107
rect 13872 30076 14381 30104
rect 13872 30064 13878 30076
rect 14369 30073 14381 30076
rect 14415 30073 14427 30107
rect 14369 30067 14427 30073
rect 17402 30064 17408 30116
rect 17460 30104 17466 30116
rect 17773 30107 17831 30113
rect 17773 30104 17785 30107
rect 17460 30076 17785 30104
rect 17460 30064 17466 30076
rect 17773 30073 17785 30076
rect 17819 30073 17831 30107
rect 17773 30067 17831 30073
rect 1397 30039 1455 30045
rect 1397 30005 1409 30039
rect 1443 30036 1455 30039
rect 1578 30036 1584 30048
rect 1443 30008 1584 30036
rect 1443 30005 1455 30008
rect 1397 29999 1455 30005
rect 1578 29996 1584 30008
rect 1636 29996 1642 30048
rect 28534 29996 28540 30048
rect 28592 29996 28598 30048
rect 1104 29946 29440 29968
rect 1104 29894 4491 29946
rect 4543 29894 4555 29946
rect 4607 29894 4619 29946
rect 4671 29894 4683 29946
rect 4735 29894 4747 29946
rect 4799 29894 11574 29946
rect 11626 29894 11638 29946
rect 11690 29894 11702 29946
rect 11754 29894 11766 29946
rect 11818 29894 11830 29946
rect 11882 29894 18657 29946
rect 18709 29894 18721 29946
rect 18773 29894 18785 29946
rect 18837 29894 18849 29946
rect 18901 29894 18913 29946
rect 18965 29894 25740 29946
rect 25792 29894 25804 29946
rect 25856 29894 25868 29946
rect 25920 29894 25932 29946
rect 25984 29894 25996 29946
rect 26048 29894 29440 29946
rect 1104 29872 29440 29894
rect 21910 29792 21916 29844
rect 21968 29832 21974 29844
rect 23661 29835 23719 29841
rect 23661 29832 23673 29835
rect 21968 29804 23673 29832
rect 21968 29792 21974 29804
rect 23661 29801 23673 29804
rect 23707 29801 23719 29835
rect 23661 29795 23719 29801
rect 5074 29724 5080 29776
rect 5132 29724 5138 29776
rect 5442 29724 5448 29776
rect 5500 29764 5506 29776
rect 5500 29736 5672 29764
rect 5500 29724 5506 29736
rect 5092 29696 5120 29724
rect 5644 29705 5672 29736
rect 14752 29736 19288 29764
rect 5629 29699 5687 29705
rect 5092 29668 5580 29696
rect 5077 29631 5135 29637
rect 5077 29597 5089 29631
rect 5123 29597 5135 29631
rect 5077 29591 5135 29597
rect 5092 29560 5120 29591
rect 5350 29588 5356 29640
rect 5408 29628 5414 29640
rect 5552 29637 5580 29668
rect 5629 29665 5641 29699
rect 5675 29665 5687 29699
rect 14090 29696 14096 29708
rect 5629 29659 5687 29665
rect 9048 29668 14096 29696
rect 9048 29640 9076 29668
rect 14090 29656 14096 29668
rect 14148 29696 14154 29708
rect 14752 29696 14780 29736
rect 14148 29668 14780 29696
rect 14148 29656 14154 29668
rect 5445 29631 5503 29637
rect 5445 29628 5457 29631
rect 5408 29600 5457 29628
rect 5408 29588 5414 29600
rect 5445 29597 5457 29600
rect 5491 29597 5503 29631
rect 5445 29591 5503 29597
rect 5537 29631 5595 29637
rect 5537 29597 5549 29631
rect 5583 29597 5595 29631
rect 5537 29591 5595 29597
rect 5718 29588 5724 29640
rect 5776 29588 5782 29640
rect 9030 29588 9036 29640
rect 9088 29588 9094 29640
rect 11241 29631 11299 29637
rect 11241 29597 11253 29631
rect 11287 29628 11299 29631
rect 11330 29628 11336 29640
rect 11287 29600 11336 29628
rect 11287 29597 11299 29600
rect 11241 29591 11299 29597
rect 11330 29588 11336 29600
rect 11388 29628 11394 29640
rect 13262 29628 13268 29640
rect 11388 29600 13268 29628
rect 11388 29588 11394 29600
rect 13262 29588 13268 29600
rect 13320 29588 13326 29640
rect 14752 29637 14780 29668
rect 16206 29656 16212 29708
rect 16264 29696 16270 29708
rect 16761 29699 16819 29705
rect 16761 29696 16773 29699
rect 16264 29668 16773 29696
rect 16264 29656 16270 29668
rect 16761 29665 16773 29668
rect 16807 29665 16819 29699
rect 19150 29696 19156 29708
rect 16761 29659 16819 29665
rect 16868 29668 19156 29696
rect 16868 29637 16896 29668
rect 19150 29656 19156 29668
rect 19208 29656 19214 29708
rect 14737 29631 14795 29637
rect 14737 29597 14749 29631
rect 14783 29597 14795 29631
rect 14737 29591 14795 29597
rect 16853 29631 16911 29637
rect 16853 29597 16865 29631
rect 16899 29597 16911 29631
rect 16853 29591 16911 29597
rect 17497 29631 17555 29637
rect 17497 29597 17509 29631
rect 17543 29597 17555 29631
rect 17497 29591 17555 29597
rect 5994 29560 6000 29572
rect 5092 29532 6000 29560
rect 5994 29520 6000 29532
rect 6052 29520 6058 29572
rect 7374 29520 7380 29572
rect 7432 29520 7438 29572
rect 7558 29520 7564 29572
rect 7616 29520 7622 29572
rect 9398 29520 9404 29572
rect 9456 29520 9462 29572
rect 12250 29560 12256 29572
rect 11072 29532 12256 29560
rect 11072 29504 11100 29532
rect 12250 29520 12256 29532
rect 12308 29520 12314 29572
rect 14274 29520 14280 29572
rect 14332 29560 14338 29572
rect 15105 29563 15163 29569
rect 15105 29560 15117 29563
rect 14332 29532 15117 29560
rect 14332 29520 14338 29532
rect 15105 29529 15117 29532
rect 15151 29529 15163 29563
rect 15105 29523 15163 29529
rect 16482 29520 16488 29572
rect 16540 29560 16546 29572
rect 17512 29560 17540 29591
rect 16540 29532 17540 29560
rect 16540 29520 16546 29532
rect 19260 29504 19288 29736
rect 20806 29588 20812 29640
rect 20864 29588 20870 29640
rect 23845 29631 23903 29637
rect 23845 29597 23857 29631
rect 23891 29628 23903 29631
rect 25222 29628 25228 29640
rect 23891 29600 25228 29628
rect 23891 29597 23903 29600
rect 23845 29591 23903 29597
rect 25222 29588 25228 29600
rect 25280 29588 25286 29640
rect 4890 29452 4896 29504
rect 4948 29452 4954 29504
rect 5261 29495 5319 29501
rect 5261 29461 5273 29495
rect 5307 29492 5319 29495
rect 5810 29492 5816 29504
rect 5307 29464 5816 29492
rect 5307 29461 5319 29464
rect 5261 29455 5319 29461
rect 5810 29452 5816 29464
rect 5868 29452 5874 29504
rect 7742 29452 7748 29504
rect 7800 29452 7806 29504
rect 11054 29452 11060 29504
rect 11112 29452 11118 29504
rect 11238 29452 11244 29504
rect 11296 29492 11302 29504
rect 11793 29495 11851 29501
rect 11793 29492 11805 29495
rect 11296 29464 11805 29492
rect 11296 29452 11302 29464
rect 11793 29461 11805 29464
rect 11839 29461 11851 29495
rect 11793 29455 11851 29461
rect 17126 29452 17132 29504
rect 17184 29492 17190 29504
rect 17221 29495 17279 29501
rect 17221 29492 17233 29495
rect 17184 29464 17233 29492
rect 17184 29452 17190 29464
rect 17221 29461 17233 29464
rect 17267 29461 17279 29495
rect 17221 29455 17279 29461
rect 17310 29452 17316 29504
rect 17368 29452 17374 29504
rect 19242 29452 19248 29504
rect 19300 29452 19306 29504
rect 20438 29452 20444 29504
rect 20496 29492 20502 29504
rect 20625 29495 20683 29501
rect 20625 29492 20637 29495
rect 20496 29464 20637 29492
rect 20496 29452 20502 29464
rect 20625 29461 20637 29464
rect 20671 29461 20683 29495
rect 20625 29455 20683 29461
rect 1104 29402 29595 29424
rect 1104 29350 8032 29402
rect 8084 29350 8096 29402
rect 8148 29350 8160 29402
rect 8212 29350 8224 29402
rect 8276 29350 8288 29402
rect 8340 29350 15115 29402
rect 15167 29350 15179 29402
rect 15231 29350 15243 29402
rect 15295 29350 15307 29402
rect 15359 29350 15371 29402
rect 15423 29350 22198 29402
rect 22250 29350 22262 29402
rect 22314 29350 22326 29402
rect 22378 29350 22390 29402
rect 22442 29350 22454 29402
rect 22506 29350 29281 29402
rect 29333 29350 29345 29402
rect 29397 29350 29409 29402
rect 29461 29350 29473 29402
rect 29525 29350 29537 29402
rect 29589 29350 29595 29402
rect 1104 29328 29595 29350
rect 3234 29288 3240 29300
rect 1412 29260 3240 29288
rect 1412 29161 1440 29260
rect 3234 29248 3240 29260
rect 3292 29288 3298 29300
rect 3292 29260 6914 29288
rect 3292 29248 3298 29260
rect 1578 29180 1584 29232
rect 1636 29220 1642 29232
rect 1673 29223 1731 29229
rect 1673 29220 1685 29223
rect 1636 29192 1685 29220
rect 1636 29180 1642 29192
rect 1673 29189 1685 29192
rect 1719 29189 1731 29223
rect 3970 29220 3976 29232
rect 2898 29192 3976 29220
rect 1673 29183 1731 29189
rect 3970 29180 3976 29192
rect 4028 29180 4034 29232
rect 6886 29220 6914 29260
rect 7098 29248 7104 29300
rect 7156 29288 7162 29300
rect 9398 29288 9404 29300
rect 7156 29260 9404 29288
rect 7156 29248 7162 29260
rect 8496 29232 8524 29260
rect 9398 29248 9404 29260
rect 9456 29248 9462 29300
rect 11238 29248 11244 29300
rect 11296 29248 11302 29300
rect 12618 29288 12624 29300
rect 11348 29260 12624 29288
rect 7466 29220 7472 29232
rect 6886 29192 7472 29220
rect 1397 29155 1455 29161
rect 1397 29121 1409 29155
rect 1443 29121 1455 29155
rect 1397 29115 1455 29121
rect 3234 29112 3240 29164
rect 3292 29112 3298 29164
rect 6822 29112 6828 29164
rect 6880 29112 6886 29164
rect 3510 29044 3516 29096
rect 3568 29044 3574 29096
rect 5077 29087 5135 29093
rect 5077 29053 5089 29087
rect 5123 29084 5135 29087
rect 5442 29084 5448 29096
rect 5123 29056 5448 29084
rect 5123 29053 5135 29056
rect 5077 29047 5135 29053
rect 5442 29044 5448 29056
rect 5500 29044 5506 29096
rect 6932 29093 6960 29192
rect 7466 29180 7472 29192
rect 7524 29180 7530 29232
rect 8478 29220 8484 29232
rect 8418 29192 8484 29220
rect 8478 29180 8484 29192
rect 8536 29180 8542 29232
rect 8757 29223 8815 29229
rect 8757 29189 8769 29223
rect 8803 29220 8815 29223
rect 9766 29220 9772 29232
rect 8803 29192 9772 29220
rect 8803 29189 8815 29192
rect 8757 29183 8815 29189
rect 9766 29180 9772 29192
rect 9824 29180 9830 29232
rect 8941 29155 8999 29161
rect 8941 29152 8953 29155
rect 8680 29124 8953 29152
rect 6917 29087 6975 29093
rect 6917 29053 6929 29087
rect 6963 29053 6975 29087
rect 7193 29087 7251 29093
rect 7193 29084 7205 29087
rect 6917 29047 6975 29053
rect 7024 29056 7205 29084
rect 3142 28976 3148 29028
rect 3200 28976 3206 29028
rect 4985 29019 5043 29025
rect 4985 28985 4997 29019
rect 5031 28985 5043 29019
rect 4985 28979 5043 28985
rect 4154 28908 4160 28960
rect 4212 28948 4218 28960
rect 5000 28948 5028 28979
rect 5166 28976 5172 29028
rect 5224 29016 5230 29028
rect 5721 29019 5779 29025
rect 5721 29016 5733 29019
rect 5224 28988 5733 29016
rect 5224 28976 5230 28988
rect 5721 28985 5733 28988
rect 5767 28985 5779 29019
rect 5721 28979 5779 28985
rect 6641 29019 6699 29025
rect 6641 28985 6653 29019
rect 6687 29016 6699 29019
rect 7024 29016 7052 29056
rect 7193 29053 7205 29056
rect 7239 29053 7251 29087
rect 7193 29047 7251 29053
rect 7558 29044 7564 29096
rect 7616 29084 7622 29096
rect 8680 29093 8708 29124
rect 8941 29121 8953 29124
rect 8987 29121 8999 29155
rect 8941 29115 8999 29121
rect 9033 29155 9091 29161
rect 9033 29121 9045 29155
rect 9079 29121 9091 29155
rect 9033 29115 9091 29121
rect 10689 29155 10747 29161
rect 10689 29121 10701 29155
rect 10735 29152 10747 29155
rect 11256 29152 11284 29248
rect 11348 29161 11376 29260
rect 12618 29248 12624 29260
rect 12676 29248 12682 29300
rect 13262 29248 13268 29300
rect 13320 29248 13326 29300
rect 16482 29248 16488 29300
rect 16540 29248 16546 29300
rect 17310 29288 17316 29300
rect 16960 29260 17316 29288
rect 12250 29180 12256 29232
rect 12308 29180 12314 29232
rect 14274 29180 14280 29232
rect 14332 29180 14338 29232
rect 16666 29220 16672 29232
rect 16316 29192 16672 29220
rect 10735 29124 11284 29152
rect 11333 29155 11391 29161
rect 10735 29121 10747 29124
rect 10689 29115 10747 29121
rect 11333 29121 11345 29155
rect 11379 29121 11391 29155
rect 11333 29115 11391 29121
rect 8665 29087 8723 29093
rect 8665 29084 8677 29087
rect 7616 29056 8677 29084
rect 7616 29044 7622 29056
rect 8665 29053 8677 29056
rect 8711 29053 8723 29087
rect 8665 29047 8723 29053
rect 9048 29016 9076 29115
rect 16206 29112 16212 29164
rect 16264 29112 16270 29164
rect 16316 29161 16344 29192
rect 16666 29180 16672 29192
rect 16724 29180 16730 29232
rect 16960 29229 16988 29260
rect 17310 29248 17316 29260
rect 17368 29248 17374 29300
rect 19150 29248 19156 29300
rect 19208 29248 19214 29300
rect 19242 29248 19248 29300
rect 19300 29288 19306 29300
rect 19300 29260 24164 29288
rect 19300 29248 19306 29260
rect 16945 29223 17003 29229
rect 16945 29189 16957 29223
rect 16991 29189 17003 29223
rect 16945 29183 17003 29189
rect 20165 29223 20223 29229
rect 20165 29189 20177 29223
rect 20211 29220 20223 29223
rect 20438 29220 20444 29232
rect 20211 29192 20444 29220
rect 20211 29189 20223 29192
rect 20165 29183 20223 29189
rect 20438 29180 20444 29192
rect 20496 29180 20502 29232
rect 20714 29180 20720 29232
rect 20772 29180 20778 29232
rect 24029 29223 24087 29229
rect 24029 29220 24041 29223
rect 22664 29192 24041 29220
rect 16301 29155 16359 29161
rect 16301 29121 16313 29155
rect 16347 29121 16359 29155
rect 16301 29115 16359 29121
rect 18046 29112 18052 29164
rect 18104 29112 18110 29164
rect 22664 29161 22692 29192
rect 24029 29189 24041 29192
rect 24075 29189 24087 29223
rect 24029 29183 24087 29189
rect 19889 29155 19947 29161
rect 19889 29121 19901 29155
rect 19935 29121 19947 29155
rect 19889 29115 19947 29121
rect 22649 29155 22707 29161
rect 22649 29121 22661 29155
rect 22695 29121 22707 29155
rect 22649 29115 22707 29121
rect 10781 29087 10839 29093
rect 10781 29053 10793 29087
rect 10827 29084 10839 29087
rect 11238 29084 11244 29096
rect 10827 29056 11244 29084
rect 10827 29053 10839 29056
rect 10781 29047 10839 29053
rect 11238 29044 11244 29056
rect 11296 29044 11302 29096
rect 11517 29087 11575 29093
rect 11517 29053 11529 29087
rect 11563 29084 11575 29087
rect 13446 29084 13452 29096
rect 11563 29056 13452 29084
rect 11563 29053 11575 29056
rect 11517 29047 11575 29053
rect 13446 29044 13452 29056
rect 13504 29044 13510 29096
rect 13722 29044 13728 29096
rect 13780 29044 13786 29096
rect 15289 29087 15347 29093
rect 15289 29053 15301 29087
rect 15335 29053 15347 29087
rect 15289 29047 15347 29053
rect 6687 28988 7052 29016
rect 8220 28988 9076 29016
rect 11057 29019 11115 29025
rect 6687 28985 6699 28988
rect 6641 28979 6699 28985
rect 5074 28948 5080 28960
rect 4212 28920 5080 28948
rect 4212 28908 4218 28920
rect 5074 28908 5080 28920
rect 5132 28908 5138 28960
rect 5258 28908 5264 28960
rect 5316 28948 5322 28960
rect 6914 28948 6920 28960
rect 5316 28920 6920 28948
rect 5316 28908 5322 28920
rect 6914 28908 6920 28920
rect 6972 28908 6978 28960
rect 7190 28908 7196 28960
rect 7248 28948 7254 28960
rect 7374 28948 7380 28960
rect 7248 28920 7380 28948
rect 7248 28908 7254 28920
rect 7374 28908 7380 28920
rect 7432 28948 7438 28960
rect 7834 28948 7840 28960
rect 7432 28920 7840 28948
rect 7432 28908 7438 28920
rect 7834 28908 7840 28920
rect 7892 28948 7898 28960
rect 8220 28948 8248 28988
rect 11057 28985 11069 29019
rect 11103 29016 11115 29019
rect 11103 28988 11376 29016
rect 11103 28985 11115 28988
rect 11057 28979 11115 28985
rect 7892 28920 8248 28948
rect 7892 28908 7898 28920
rect 8754 28908 8760 28960
rect 8812 28908 8818 28960
rect 11146 28908 11152 28960
rect 11204 28908 11210 28960
rect 11348 28948 11376 28988
rect 11774 28951 11832 28957
rect 11774 28948 11786 28951
rect 11348 28920 11786 28948
rect 11774 28917 11786 28920
rect 11820 28917 11832 28951
rect 11774 28911 11832 28917
rect 15197 28951 15255 28957
rect 15197 28917 15209 28951
rect 15243 28948 15255 28951
rect 15304 28948 15332 29047
rect 16574 29044 16580 29096
rect 16632 29084 16638 29096
rect 16669 29087 16727 29093
rect 16669 29084 16681 29087
rect 16632 29056 16681 29084
rect 16632 29044 16638 29056
rect 16669 29053 16681 29056
rect 16715 29053 16727 29087
rect 16669 29047 16727 29053
rect 18414 29044 18420 29096
rect 18472 29084 18478 29096
rect 18509 29087 18567 29093
rect 18509 29084 18521 29087
rect 18472 29056 18521 29084
rect 18472 29044 18478 29056
rect 18509 29053 18521 29056
rect 18555 29053 18567 29087
rect 19904 29084 19932 29115
rect 22830 29112 22836 29164
rect 22888 29152 22894 29164
rect 23109 29155 23167 29161
rect 23109 29152 23121 29155
rect 22888 29124 23121 29152
rect 22888 29112 22894 29124
rect 23109 29121 23121 29124
rect 23155 29121 23167 29155
rect 23109 29115 23167 29121
rect 23293 29155 23351 29161
rect 23293 29121 23305 29155
rect 23339 29121 23351 29155
rect 23293 29115 23351 29121
rect 20162 29084 20168 29096
rect 19904 29056 20168 29084
rect 18509 29047 18567 29053
rect 20162 29044 20168 29056
rect 20220 29044 20226 29096
rect 22094 29044 22100 29096
rect 22152 29084 22158 29096
rect 22557 29087 22615 29093
rect 22557 29084 22569 29087
rect 22152 29056 22569 29084
rect 22152 29044 22158 29056
rect 22557 29053 22569 29056
rect 22603 29084 22615 29087
rect 23308 29084 23336 29115
rect 22603 29056 23336 29084
rect 22603 29053 22615 29056
rect 22557 29047 22615 29053
rect 23382 29044 23388 29096
rect 23440 29044 23446 29096
rect 24136 29084 24164 29260
rect 28534 29248 28540 29300
rect 28592 29248 28598 29300
rect 24397 29155 24455 29161
rect 24397 29121 24409 29155
rect 24443 29152 24455 29155
rect 28552 29152 28580 29248
rect 24443 29124 28580 29152
rect 24443 29121 24455 29124
rect 24397 29115 24455 29121
rect 24486 29084 24492 29096
rect 24136 29056 24492 29084
rect 24486 29044 24492 29056
rect 24544 29084 24550 29096
rect 24673 29087 24731 29093
rect 24673 29084 24685 29087
rect 24544 29056 24685 29084
rect 24544 29044 24550 29056
rect 24673 29053 24685 29056
rect 24719 29053 24731 29087
rect 24673 29047 24731 29053
rect 23198 29016 23204 29028
rect 21284 28988 22094 29016
rect 15562 28948 15568 28960
rect 15243 28920 15568 28948
rect 15243 28917 15255 28920
rect 15197 28911 15255 28917
rect 15562 28908 15568 28920
rect 15620 28908 15626 28960
rect 15930 28908 15936 28960
rect 15988 28908 15994 28960
rect 18322 28908 18328 28960
rect 18380 28948 18386 28960
rect 18417 28951 18475 28957
rect 18417 28948 18429 28951
rect 18380 28920 18429 28948
rect 18380 28908 18386 28920
rect 18417 28917 18429 28920
rect 18463 28917 18475 28951
rect 18417 28911 18475 28917
rect 20714 28908 20720 28960
rect 20772 28948 20778 28960
rect 21284 28948 21312 28988
rect 20772 28920 21312 28948
rect 20772 28908 20778 28920
rect 21358 28908 21364 28960
rect 21416 28948 21422 28960
rect 21637 28951 21695 28957
rect 21637 28948 21649 28951
rect 21416 28920 21649 28948
rect 21416 28908 21422 28920
rect 21637 28917 21649 28920
rect 21683 28917 21695 28951
rect 22066 28948 22094 28988
rect 23032 28988 23204 29016
rect 22922 28948 22928 28960
rect 22066 28920 22928 28948
rect 21637 28911 21695 28917
rect 22922 28908 22928 28920
rect 22980 28908 22986 28960
rect 23032 28957 23060 28988
rect 23198 28976 23204 28988
rect 23256 28976 23262 29028
rect 23017 28951 23075 28957
rect 23017 28917 23029 28951
rect 23063 28917 23075 28951
rect 23017 28911 23075 28917
rect 23106 28908 23112 28960
rect 23164 28908 23170 28960
rect 1104 28858 29440 28880
rect 1104 28806 4491 28858
rect 4543 28806 4555 28858
rect 4607 28806 4619 28858
rect 4671 28806 4683 28858
rect 4735 28806 4747 28858
rect 4799 28806 11574 28858
rect 11626 28806 11638 28858
rect 11690 28806 11702 28858
rect 11754 28806 11766 28858
rect 11818 28806 11830 28858
rect 11882 28806 18657 28858
rect 18709 28806 18721 28858
rect 18773 28806 18785 28858
rect 18837 28806 18849 28858
rect 18901 28806 18913 28858
rect 18965 28806 25740 28858
rect 25792 28806 25804 28858
rect 25856 28806 25868 28858
rect 25920 28806 25932 28858
rect 25984 28806 25996 28858
rect 26048 28806 29440 28858
rect 1104 28784 29440 28806
rect 5166 28744 5172 28756
rect 3252 28716 5172 28744
rect 3252 28549 3280 28716
rect 5166 28704 5172 28716
rect 5224 28704 5230 28756
rect 5718 28704 5724 28756
rect 5776 28744 5782 28756
rect 6089 28747 6147 28753
rect 6089 28744 6101 28747
rect 5776 28716 6101 28744
rect 5776 28704 5782 28716
rect 6089 28713 6101 28716
rect 6135 28744 6147 28747
rect 7377 28747 7435 28753
rect 6135 28716 6500 28744
rect 6135 28713 6147 28716
rect 6089 28707 6147 28713
rect 3329 28611 3387 28617
rect 3329 28577 3341 28611
rect 3375 28608 3387 28611
rect 4246 28608 4252 28620
rect 3375 28580 4252 28608
rect 3375 28577 3387 28580
rect 3329 28571 3387 28577
rect 4246 28568 4252 28580
rect 4304 28568 4310 28620
rect 4341 28611 4399 28617
rect 4341 28577 4353 28611
rect 4387 28608 4399 28611
rect 4982 28608 4988 28620
rect 4387 28580 4988 28608
rect 4387 28577 4399 28580
rect 4341 28571 4399 28577
rect 4982 28568 4988 28580
rect 5040 28568 5046 28620
rect 6362 28568 6368 28620
rect 6420 28568 6426 28620
rect 3237 28543 3295 28549
rect 3237 28509 3249 28543
rect 3283 28509 3295 28543
rect 3237 28503 3295 28509
rect 4065 28543 4123 28549
rect 4065 28509 4077 28543
rect 4111 28540 4123 28543
rect 4154 28540 4160 28552
rect 4111 28512 4160 28540
rect 4111 28509 4123 28512
rect 4065 28503 4123 28509
rect 4154 28500 4160 28512
rect 4212 28500 4218 28552
rect 3881 28475 3939 28481
rect 3881 28441 3893 28475
rect 3927 28472 3939 28475
rect 4617 28475 4675 28481
rect 3927 28444 4568 28472
rect 3927 28441 3939 28444
rect 3881 28435 3939 28441
rect 4172 28416 4200 28444
rect 3602 28364 3608 28416
rect 3660 28364 3666 28416
rect 4154 28364 4160 28416
rect 4212 28364 4218 28416
rect 4249 28407 4307 28413
rect 4249 28373 4261 28407
rect 4295 28404 4307 28407
rect 4338 28404 4344 28416
rect 4295 28376 4344 28404
rect 4295 28373 4307 28376
rect 4249 28367 4307 28373
rect 4338 28364 4344 28376
rect 4396 28364 4402 28416
rect 4540 28404 4568 28444
rect 4617 28441 4629 28475
rect 4663 28472 4675 28475
rect 4890 28472 4896 28484
rect 4663 28444 4896 28472
rect 4663 28441 4675 28444
rect 4617 28435 4675 28441
rect 4890 28432 4896 28444
rect 4948 28432 4954 28484
rect 5258 28432 5264 28484
rect 5316 28432 5322 28484
rect 6178 28432 6184 28484
rect 6236 28432 6242 28484
rect 6380 28481 6408 28568
rect 6472 28552 6500 28716
rect 7377 28713 7389 28747
rect 7423 28744 7435 28747
rect 7742 28744 7748 28756
rect 7423 28716 7748 28744
rect 7423 28713 7435 28716
rect 7377 28707 7435 28713
rect 7742 28704 7748 28716
rect 7800 28704 7806 28756
rect 7837 28747 7895 28753
rect 7837 28713 7849 28747
rect 7883 28744 7895 28747
rect 7883 28716 9076 28744
rect 7883 28713 7895 28716
rect 7837 28707 7895 28713
rect 6932 28648 8064 28676
rect 6454 28500 6460 28552
rect 6512 28500 6518 28552
rect 6932 28549 6960 28648
rect 7116 28580 7972 28608
rect 7116 28549 7144 28580
rect 6917 28543 6975 28549
rect 6917 28509 6929 28543
rect 6963 28509 6975 28543
rect 6917 28503 6975 28509
rect 7101 28543 7159 28549
rect 7101 28509 7113 28543
rect 7147 28509 7159 28543
rect 7101 28503 7159 28509
rect 7282 28500 7288 28552
rect 7340 28500 7346 28552
rect 7558 28500 7564 28552
rect 7616 28540 7622 28552
rect 7616 28512 7696 28540
rect 7616 28500 7622 28512
rect 6365 28475 6423 28481
rect 6365 28441 6377 28475
rect 6411 28441 6423 28475
rect 6365 28435 6423 28441
rect 6932 28444 7144 28472
rect 5350 28404 5356 28416
rect 4540 28376 5356 28404
rect 5350 28364 5356 28376
rect 5408 28404 5414 28416
rect 6549 28407 6607 28413
rect 6549 28404 6561 28407
rect 5408 28376 6561 28404
rect 5408 28364 5414 28376
rect 6549 28373 6561 28376
rect 6595 28373 6607 28407
rect 6549 28367 6607 28373
rect 6733 28407 6791 28413
rect 6733 28373 6745 28407
rect 6779 28404 6791 28407
rect 6932 28404 6960 28444
rect 7116 28416 7144 28444
rect 7190 28432 7196 28484
rect 7248 28432 7254 28484
rect 7300 28472 7328 28500
rect 7668 28481 7696 28512
rect 7653 28475 7711 28481
rect 7300 28444 7604 28472
rect 6779 28376 6960 28404
rect 6779 28373 6791 28376
rect 6733 28367 6791 28373
rect 7006 28364 7012 28416
rect 7064 28364 7070 28416
rect 7098 28364 7104 28416
rect 7156 28364 7162 28416
rect 7282 28364 7288 28416
rect 7340 28404 7346 28416
rect 7576 28413 7604 28444
rect 7653 28441 7665 28475
rect 7699 28441 7711 28475
rect 7653 28435 7711 28441
rect 7834 28432 7840 28484
rect 7892 28481 7898 28484
rect 7892 28475 7911 28481
rect 7899 28441 7911 28475
rect 7892 28435 7911 28441
rect 7892 28432 7898 28435
rect 7393 28407 7451 28413
rect 7393 28404 7405 28407
rect 7340 28376 7405 28404
rect 7340 28364 7346 28376
rect 7393 28373 7405 28376
rect 7439 28373 7451 28407
rect 7393 28367 7451 28373
rect 7561 28407 7619 28413
rect 7561 28373 7573 28407
rect 7607 28373 7619 28407
rect 7944 28404 7972 28580
rect 8036 28472 8064 28648
rect 8205 28611 8263 28617
rect 8205 28577 8217 28611
rect 8251 28608 8263 28611
rect 8754 28608 8760 28620
rect 8251 28580 8760 28608
rect 8251 28577 8263 28580
rect 8205 28571 8263 28577
rect 8754 28568 8760 28580
rect 8812 28568 8818 28620
rect 9048 28608 9076 28716
rect 9766 28704 9772 28756
rect 9824 28704 9830 28756
rect 10321 28747 10379 28753
rect 10321 28713 10333 28747
rect 10367 28744 10379 28747
rect 12437 28747 12495 28753
rect 12437 28744 12449 28747
rect 10367 28716 12449 28744
rect 10367 28713 10379 28716
rect 10321 28707 10379 28713
rect 12437 28713 12449 28716
rect 12483 28713 12495 28747
rect 12437 28707 12495 28713
rect 12618 28704 12624 28756
rect 12676 28704 12682 28756
rect 12894 28704 12900 28756
rect 12952 28744 12958 28756
rect 13449 28747 13507 28753
rect 13449 28744 13461 28747
rect 12952 28716 13461 28744
rect 12952 28704 12958 28716
rect 13449 28713 13461 28716
rect 13495 28713 13507 28747
rect 13449 28707 13507 28713
rect 13722 28704 13728 28756
rect 13780 28744 13786 28756
rect 14921 28747 14979 28753
rect 14921 28744 14933 28747
rect 13780 28716 14933 28744
rect 13780 28704 13786 28716
rect 14921 28713 14933 28716
rect 14967 28713 14979 28747
rect 14921 28707 14979 28713
rect 16117 28747 16175 28753
rect 16117 28713 16129 28747
rect 16163 28744 16175 28747
rect 16206 28744 16212 28756
rect 16163 28716 16212 28744
rect 16163 28713 16175 28716
rect 16117 28707 16175 28713
rect 16206 28704 16212 28716
rect 16264 28704 16270 28756
rect 16666 28704 16672 28756
rect 16724 28704 16730 28756
rect 20349 28747 20407 28753
rect 20349 28713 20361 28747
rect 20395 28713 20407 28747
rect 20349 28707 20407 28713
rect 20533 28747 20591 28753
rect 20533 28713 20545 28747
rect 20579 28744 20591 28747
rect 20806 28744 20812 28756
rect 20579 28716 20812 28744
rect 20579 28713 20591 28716
rect 20533 28707 20591 28713
rect 15841 28679 15899 28685
rect 15841 28676 15853 28679
rect 13188 28648 15853 28676
rect 9125 28611 9183 28617
rect 9125 28608 9137 28611
rect 9048 28580 9137 28608
rect 9125 28577 9137 28580
rect 9171 28608 9183 28611
rect 9398 28608 9404 28620
rect 9171 28580 9404 28608
rect 9171 28577 9183 28580
rect 9125 28571 9183 28577
rect 9398 28568 9404 28580
rect 9456 28568 9462 28620
rect 10689 28611 10747 28617
rect 10689 28577 10701 28611
rect 10735 28608 10747 28611
rect 11146 28608 11152 28620
rect 10735 28580 11152 28608
rect 10735 28577 10747 28580
rect 10689 28571 10747 28577
rect 11146 28568 11152 28580
rect 11204 28568 11210 28620
rect 11238 28568 11244 28620
rect 11296 28608 11302 28620
rect 11296 28580 12388 28608
rect 11296 28568 11302 28580
rect 10410 28500 10416 28552
rect 10468 28500 10474 28552
rect 8757 28475 8815 28481
rect 8757 28472 8769 28475
rect 8036 28444 8769 28472
rect 8757 28441 8769 28444
rect 8803 28441 8815 28475
rect 8757 28435 8815 28441
rect 9950 28432 9956 28484
rect 10008 28432 10014 28484
rect 10137 28475 10195 28481
rect 10137 28441 10149 28475
rect 10183 28441 10195 28475
rect 10137 28435 10195 28441
rect 8021 28407 8079 28413
rect 8021 28404 8033 28407
rect 7944 28376 8033 28404
rect 7561 28367 7619 28373
rect 8021 28373 8033 28376
rect 8067 28404 8079 28407
rect 8570 28404 8576 28416
rect 8067 28376 8576 28404
rect 8067 28373 8079 28376
rect 8021 28367 8079 28373
rect 8570 28364 8576 28376
rect 8628 28364 8634 28416
rect 10152 28404 10180 28435
rect 11146 28432 11152 28484
rect 11204 28432 11210 28484
rect 12253 28475 12311 28481
rect 12253 28441 12265 28475
rect 12299 28441 12311 28475
rect 12360 28472 12388 28580
rect 13188 28549 13216 28648
rect 15841 28645 15853 28648
rect 15887 28676 15899 28679
rect 15887 28648 16068 28676
rect 15887 28645 15899 28648
rect 15841 28639 15899 28645
rect 13630 28568 13636 28620
rect 13688 28568 13694 28620
rect 15381 28611 15439 28617
rect 15381 28577 15393 28611
rect 15427 28608 15439 28611
rect 15930 28608 15936 28620
rect 15427 28580 15936 28608
rect 15427 28577 15439 28580
rect 15381 28571 15439 28577
rect 15930 28568 15936 28580
rect 15988 28568 15994 28620
rect 13173 28543 13231 28549
rect 13173 28509 13185 28543
rect 13219 28509 13231 28543
rect 13173 28503 13231 28509
rect 13354 28500 13360 28552
rect 13412 28500 13418 28552
rect 13725 28543 13783 28549
rect 13725 28509 13737 28543
rect 13771 28540 13783 28543
rect 13998 28540 14004 28552
rect 13771 28512 14004 28540
rect 13771 28509 13783 28512
rect 13725 28503 13783 28509
rect 13998 28500 14004 28512
rect 14056 28500 14062 28552
rect 14185 28543 14243 28549
rect 14185 28509 14197 28543
rect 14231 28540 14243 28543
rect 14458 28540 14464 28552
rect 14231 28512 14464 28540
rect 14231 28509 14243 28512
rect 14185 28503 14243 28509
rect 14458 28500 14464 28512
rect 14516 28500 14522 28552
rect 15105 28543 15163 28549
rect 15105 28509 15117 28543
rect 15151 28509 15163 28543
rect 15105 28503 15163 28509
rect 15289 28543 15347 28549
rect 15289 28509 15301 28543
rect 15335 28509 15347 28543
rect 15289 28503 15347 28509
rect 12453 28475 12511 28481
rect 12453 28472 12465 28475
rect 12360 28444 12465 28472
rect 12253 28435 12311 28441
rect 12453 28441 12465 28444
rect 12499 28441 12511 28475
rect 12453 28435 12511 28441
rect 13449 28475 13507 28481
rect 13449 28441 13461 28475
rect 13495 28472 13507 28475
rect 13630 28472 13636 28484
rect 13495 28444 13636 28472
rect 13495 28441 13507 28444
rect 13449 28435 13507 28441
rect 12158 28404 12164 28416
rect 10152 28376 12164 28404
rect 12158 28364 12164 28376
rect 12216 28364 12222 28416
rect 12268 28404 12296 28435
rect 13630 28432 13636 28444
rect 13688 28432 13694 28484
rect 15120 28472 15148 28503
rect 13832 28444 15148 28472
rect 15304 28472 15332 28503
rect 15562 28500 15568 28552
rect 15620 28500 15626 28552
rect 16040 28549 16068 28648
rect 18138 28636 18144 28688
rect 18196 28676 18202 28688
rect 19242 28676 19248 28688
rect 18196 28648 19248 28676
rect 18196 28636 18202 28648
rect 19242 28636 19248 28648
rect 19300 28636 19306 28688
rect 19334 28636 19340 28688
rect 19392 28676 19398 28688
rect 20364 28676 20392 28707
rect 20806 28704 20812 28716
rect 20864 28704 20870 28756
rect 20916 28716 21220 28744
rect 20916 28676 20944 28716
rect 19392 28648 19564 28676
rect 20364 28648 20944 28676
rect 21192 28676 21220 28716
rect 21266 28704 21272 28756
rect 21324 28744 21330 28756
rect 21821 28747 21879 28753
rect 21821 28744 21833 28747
rect 21324 28716 21833 28744
rect 21324 28704 21330 28716
rect 21821 28713 21833 28716
rect 21867 28744 21879 28747
rect 22370 28744 22376 28756
rect 21867 28716 22376 28744
rect 21867 28713 21879 28716
rect 21821 28707 21879 28713
rect 22370 28704 22376 28716
rect 22428 28704 22434 28756
rect 22922 28704 22928 28756
rect 22980 28744 22986 28756
rect 22980 28716 23888 28744
rect 22980 28704 22986 28716
rect 22189 28679 22247 28685
rect 22189 28676 22201 28679
rect 21192 28648 22201 28676
rect 19392 28636 19398 28648
rect 17037 28611 17095 28617
rect 17037 28577 17049 28611
rect 17083 28608 17095 28611
rect 17126 28608 17132 28620
rect 17083 28580 17132 28608
rect 17083 28577 17095 28580
rect 17037 28571 17095 28577
rect 17126 28568 17132 28580
rect 17184 28568 17190 28620
rect 15657 28543 15715 28549
rect 15657 28509 15669 28543
rect 15703 28509 15715 28543
rect 15657 28503 15715 28509
rect 16025 28543 16083 28549
rect 16025 28509 16037 28543
rect 16071 28509 16083 28543
rect 16025 28503 16083 28509
rect 16209 28543 16267 28549
rect 16209 28509 16221 28543
rect 16255 28540 16267 28543
rect 16482 28540 16488 28552
rect 16255 28512 16488 28540
rect 16255 28509 16267 28512
rect 16209 28503 16267 28509
rect 15672 28472 15700 28503
rect 15304 28444 15700 28472
rect 16040 28472 16068 28503
rect 16482 28500 16488 28512
rect 16540 28500 16546 28552
rect 16574 28500 16580 28552
rect 16632 28540 16638 28552
rect 16761 28543 16819 28549
rect 16761 28540 16773 28543
rect 16632 28512 16773 28540
rect 16632 28500 16638 28512
rect 16761 28509 16773 28512
rect 16807 28509 16819 28543
rect 18156 28526 18184 28636
rect 19536 28617 19564 28648
rect 22189 28645 22201 28648
rect 22235 28645 22247 28679
rect 22189 28639 22247 28645
rect 19521 28611 19579 28617
rect 19521 28577 19533 28611
rect 19567 28577 19579 28611
rect 19521 28571 19579 28577
rect 19245 28543 19303 28549
rect 16761 28503 16819 28509
rect 19245 28509 19257 28543
rect 19291 28509 19303 28543
rect 19245 28503 19303 28509
rect 19337 28543 19395 28549
rect 19337 28509 19349 28543
rect 19383 28540 19395 28543
rect 19426 28540 19432 28552
rect 19383 28512 19432 28540
rect 19383 28509 19395 28512
rect 19337 28503 19395 28509
rect 16298 28472 16304 28484
rect 16040 28444 16304 28472
rect 12342 28404 12348 28416
rect 12268 28376 12348 28404
rect 12342 28364 12348 28376
rect 12400 28364 12406 28416
rect 13265 28407 13323 28413
rect 13265 28373 13277 28407
rect 13311 28404 13323 28407
rect 13832 28404 13860 28444
rect 13311 28376 13860 28404
rect 13311 28373 13323 28376
rect 13265 28367 13323 28373
rect 13906 28364 13912 28416
rect 13964 28364 13970 28416
rect 14734 28364 14740 28416
rect 14792 28364 14798 28416
rect 15010 28364 15016 28416
rect 15068 28404 15074 28416
rect 15304 28404 15332 28444
rect 16298 28432 16304 28444
rect 16356 28432 16362 28484
rect 19260 28472 19288 28503
rect 19426 28500 19432 28512
rect 19484 28500 19490 28552
rect 19536 28540 19564 28571
rect 20162 28568 20168 28620
rect 20220 28608 20226 28620
rect 21008 28608 21128 28616
rect 22465 28611 22523 28617
rect 22465 28608 22477 28611
rect 20220 28588 22477 28608
rect 20220 28580 21036 28588
rect 21100 28580 22477 28588
rect 20220 28568 20226 28580
rect 22465 28577 22477 28580
rect 22511 28577 22523 28611
rect 22465 28571 22523 28577
rect 22741 28611 22799 28617
rect 22741 28577 22753 28611
rect 22787 28608 22799 28611
rect 23106 28608 23112 28620
rect 22787 28580 23112 28608
rect 22787 28577 22799 28580
rect 22741 28571 22799 28577
rect 19536 28512 20208 28540
rect 20180 28481 20208 28512
rect 20806 28500 20812 28552
rect 20864 28500 20870 28552
rect 20901 28543 20959 28549
rect 20901 28509 20913 28543
rect 20947 28509 20959 28543
rect 20901 28503 20959 28509
rect 20994 28543 21052 28549
rect 20994 28509 21006 28543
rect 21040 28509 21052 28543
rect 20994 28503 21052 28509
rect 21085 28543 21143 28549
rect 21085 28509 21097 28543
rect 21131 28540 21143 28543
rect 21358 28540 21364 28552
rect 21131 28512 21364 28540
rect 21131 28509 21143 28512
rect 21085 28503 21143 28509
rect 20165 28475 20223 28481
rect 19260 28444 19656 28472
rect 15068 28376 15332 28404
rect 16316 28404 16344 28432
rect 18046 28404 18052 28416
rect 16316 28376 18052 28404
rect 15068 28364 15074 28376
rect 18046 28364 18052 28376
rect 18104 28364 18110 28416
rect 18414 28364 18420 28416
rect 18472 28404 18478 28416
rect 18509 28407 18567 28413
rect 18509 28404 18521 28407
rect 18472 28376 18521 28404
rect 18472 28364 18478 28376
rect 18509 28373 18521 28376
rect 18555 28373 18567 28407
rect 18509 28367 18567 28373
rect 19426 28364 19432 28416
rect 19484 28404 19490 28416
rect 19521 28407 19579 28413
rect 19521 28404 19533 28407
rect 19484 28376 19533 28404
rect 19484 28364 19490 28376
rect 19521 28373 19533 28376
rect 19567 28373 19579 28407
rect 19628 28404 19656 28444
rect 20165 28441 20177 28475
rect 20211 28441 20223 28475
rect 20165 28435 20223 28441
rect 20381 28475 20439 28481
rect 20381 28441 20393 28475
rect 20427 28472 20439 28475
rect 20427 28444 20668 28472
rect 20427 28441 20439 28444
rect 20381 28435 20439 28441
rect 20254 28404 20260 28416
rect 19628 28376 20260 28404
rect 19521 28367 19579 28373
rect 20254 28364 20260 28376
rect 20312 28364 20318 28416
rect 20640 28413 20668 28444
rect 20625 28407 20683 28413
rect 20625 28373 20637 28407
rect 20671 28373 20683 28407
rect 20916 28404 20944 28503
rect 21024 28472 21052 28503
rect 21358 28500 21364 28512
rect 21416 28500 21422 28552
rect 21453 28543 21511 28549
rect 21453 28509 21465 28543
rect 21499 28540 21511 28543
rect 21634 28540 21640 28552
rect 21499 28512 21640 28540
rect 21499 28509 21511 28512
rect 21453 28503 21511 28509
rect 21634 28500 21640 28512
rect 21692 28500 21698 28552
rect 21818 28549 21824 28552
rect 21811 28543 21824 28549
rect 21811 28540 21823 28543
rect 21744 28512 21823 28540
rect 21744 28472 21772 28512
rect 21811 28509 21823 28512
rect 21811 28503 21824 28509
rect 21818 28500 21824 28503
rect 21876 28500 21882 28552
rect 22281 28543 22339 28549
rect 22281 28540 22293 28543
rect 21928 28512 22293 28540
rect 21024 28444 21772 28472
rect 21266 28404 21272 28416
rect 20916 28376 21272 28404
rect 20625 28367 20683 28373
rect 21266 28364 21272 28376
rect 21324 28364 21330 28416
rect 21358 28364 21364 28416
rect 21416 28404 21422 28416
rect 21928 28404 21956 28512
rect 22281 28509 22293 28512
rect 22327 28509 22339 28543
rect 22281 28503 22339 28509
rect 22370 28500 22376 28552
rect 22428 28500 22434 28552
rect 22094 28432 22100 28484
rect 22152 28432 22158 28484
rect 21416 28376 21956 28404
rect 21416 28364 21422 28376
rect 22002 28364 22008 28416
rect 22060 28364 22066 28416
rect 22388 28404 22416 28500
rect 22480 28472 22508 28571
rect 23106 28568 23112 28580
rect 23164 28568 23170 28620
rect 23860 28608 23888 28716
rect 24210 28636 24216 28688
rect 24268 28676 24274 28688
rect 24268 28648 25268 28676
rect 24268 28636 24274 28648
rect 25240 28617 25268 28648
rect 24765 28611 24823 28617
rect 24765 28608 24777 28611
rect 23860 28580 24777 28608
rect 23860 28526 23888 28580
rect 24765 28577 24777 28580
rect 24811 28577 24823 28611
rect 24765 28571 24823 28577
rect 25225 28611 25283 28617
rect 25225 28577 25237 28611
rect 25271 28577 25283 28611
rect 25225 28571 25283 28577
rect 24026 28500 24032 28552
rect 24084 28540 24090 28552
rect 24486 28540 24492 28552
rect 24084 28512 24492 28540
rect 24084 28500 24090 28512
rect 24486 28500 24492 28512
rect 24544 28500 24550 28552
rect 22646 28472 22652 28484
rect 22480 28444 22652 28472
rect 22646 28432 22652 28444
rect 22704 28432 22710 28484
rect 24670 28472 24676 28484
rect 24044 28444 24676 28472
rect 23382 28404 23388 28416
rect 22388 28376 23388 28404
rect 23382 28364 23388 28376
rect 23440 28404 23446 28416
rect 24044 28404 24072 28444
rect 24670 28432 24676 28444
rect 24728 28432 24734 28484
rect 23440 28376 24072 28404
rect 23440 28364 23446 28376
rect 24394 28364 24400 28416
rect 24452 28404 24458 28416
rect 25869 28407 25927 28413
rect 25869 28404 25881 28407
rect 24452 28376 25881 28404
rect 24452 28364 24458 28376
rect 25869 28373 25881 28376
rect 25915 28373 25927 28407
rect 25869 28367 25927 28373
rect 1104 28314 29595 28336
rect 1104 28262 8032 28314
rect 8084 28262 8096 28314
rect 8148 28262 8160 28314
rect 8212 28262 8224 28314
rect 8276 28262 8288 28314
rect 8340 28262 15115 28314
rect 15167 28262 15179 28314
rect 15231 28262 15243 28314
rect 15295 28262 15307 28314
rect 15359 28262 15371 28314
rect 15423 28262 22198 28314
rect 22250 28262 22262 28314
rect 22314 28262 22326 28314
rect 22378 28262 22390 28314
rect 22442 28262 22454 28314
rect 22506 28262 29281 28314
rect 29333 28262 29345 28314
rect 29397 28262 29409 28314
rect 29461 28262 29473 28314
rect 29525 28262 29537 28314
rect 29589 28262 29595 28314
rect 1104 28240 29595 28262
rect 3421 28203 3479 28209
rect 3421 28169 3433 28203
rect 3467 28200 3479 28203
rect 3510 28200 3516 28212
rect 3467 28172 3516 28200
rect 3467 28169 3479 28172
rect 3421 28163 3479 28169
rect 3510 28160 3516 28172
rect 3568 28160 3574 28212
rect 3602 28160 3608 28212
rect 3660 28160 3666 28212
rect 5258 28200 5264 28212
rect 4356 28172 5264 28200
rect 3620 28132 3648 28160
rect 3973 28135 4031 28141
rect 3973 28132 3985 28135
rect 3620 28104 3985 28132
rect 3973 28101 3985 28104
rect 4019 28101 4031 28135
rect 4356 28132 4384 28172
rect 5258 28160 5264 28172
rect 5316 28160 5322 28212
rect 5442 28160 5448 28212
rect 5500 28160 5506 28212
rect 5994 28160 6000 28212
rect 6052 28160 6058 28212
rect 7006 28160 7012 28212
rect 7064 28160 7070 28212
rect 7282 28160 7288 28212
rect 7340 28160 7346 28212
rect 8570 28160 8576 28212
rect 8628 28200 8634 28212
rect 8628 28172 9260 28200
rect 8628 28160 8634 28172
rect 4430 28132 4436 28144
rect 4356 28104 4436 28132
rect 3973 28095 4031 28101
rect 4430 28092 4436 28104
rect 4488 28092 4494 28144
rect 5460 28132 5488 28160
rect 6178 28132 6184 28144
rect 5460 28104 6184 28132
rect 6178 28092 6184 28104
rect 6236 28132 6242 28144
rect 7024 28132 7052 28160
rect 7929 28135 7987 28141
rect 7929 28132 7941 28135
rect 6236 28104 6868 28132
rect 7024 28104 7941 28132
rect 6236 28092 6242 28104
rect 3602 28024 3608 28076
rect 3660 28024 3666 28076
rect 6840 28073 6868 28104
rect 7929 28101 7941 28104
rect 7975 28101 7987 28135
rect 7929 28095 7987 28101
rect 6365 28067 6423 28073
rect 6365 28033 6377 28067
rect 6411 28064 6423 28067
rect 6825 28067 6883 28073
rect 6411 28036 6776 28064
rect 6411 28033 6423 28036
rect 6365 28027 6423 28033
rect 3697 27999 3755 28005
rect 3697 27965 3709 27999
rect 3743 27996 3755 27999
rect 4982 27996 4988 28008
rect 3743 27968 4988 27996
rect 3743 27965 3755 27968
rect 3697 27959 3755 27965
rect 4982 27956 4988 27968
rect 5040 27956 5046 28008
rect 5537 27999 5595 28005
rect 5537 27965 5549 27999
rect 5583 27996 5595 27999
rect 5583 27968 6224 27996
rect 5583 27965 5595 27968
rect 5537 27959 5595 27965
rect 5810 27888 5816 27940
rect 5868 27888 5874 27940
rect 6196 27928 6224 27968
rect 6454 27956 6460 28008
rect 6512 27996 6518 28008
rect 6641 27999 6699 28005
rect 6641 27996 6653 27999
rect 6512 27968 6653 27996
rect 6512 27956 6518 27968
rect 6641 27965 6653 27968
rect 6687 27965 6699 27999
rect 6748 27996 6776 28036
rect 6825 28033 6837 28067
rect 6871 28033 6883 28067
rect 6825 28027 6883 28033
rect 7098 28024 7104 28076
rect 7156 28024 7162 28076
rect 7285 28067 7343 28073
rect 7285 28033 7297 28067
rect 7331 28064 7343 28067
rect 7558 28064 7564 28076
rect 7331 28036 7564 28064
rect 7331 28033 7343 28036
rect 7285 28027 7343 28033
rect 7300 27996 7328 28027
rect 7558 28024 7564 28036
rect 7616 28024 7622 28076
rect 9030 28024 9036 28076
rect 9088 28024 9094 28076
rect 9232 28064 9260 28172
rect 9398 28160 9404 28212
rect 9456 28160 9462 28212
rect 9861 28203 9919 28209
rect 9861 28169 9873 28203
rect 9907 28200 9919 28203
rect 9950 28200 9956 28212
rect 9907 28172 9956 28200
rect 9907 28169 9919 28172
rect 9861 28163 9919 28169
rect 9950 28160 9956 28172
rect 10008 28200 10014 28212
rect 10008 28172 11100 28200
rect 10008 28160 10014 28172
rect 9416 28132 9444 28160
rect 11072 28132 11100 28172
rect 11238 28160 11244 28212
rect 11296 28160 11302 28212
rect 11701 28203 11759 28209
rect 11701 28169 11713 28203
rect 11747 28200 11759 28203
rect 12158 28200 12164 28212
rect 11747 28172 12164 28200
rect 11747 28169 11759 28172
rect 11701 28163 11759 28169
rect 11885 28135 11943 28141
rect 11885 28132 11897 28135
rect 9416 28104 10824 28132
rect 9306 28064 9312 28076
rect 9232 28036 9312 28064
rect 9306 28024 9312 28036
rect 9364 28064 9370 28076
rect 10796 28073 10824 28104
rect 11072 28104 11897 28132
rect 11072 28073 11100 28104
rect 11885 28101 11897 28104
rect 11931 28101 11943 28135
rect 11885 28095 11943 28101
rect 9677 28067 9735 28073
rect 9677 28064 9689 28067
rect 9364 28036 9689 28064
rect 9364 28024 9370 28036
rect 9677 28033 9689 28036
rect 9723 28033 9735 28067
rect 10413 28067 10471 28073
rect 10413 28064 10425 28067
rect 9677 28027 9735 28033
rect 9784 28036 10425 28064
rect 9784 28008 9812 28036
rect 10413 28033 10425 28036
rect 10459 28033 10471 28067
rect 10413 28027 10471 28033
rect 10781 28067 10839 28073
rect 10781 28033 10793 28067
rect 10827 28033 10839 28067
rect 10781 28027 10839 28033
rect 11057 28067 11115 28073
rect 11057 28033 11069 28067
rect 11103 28033 11115 28067
rect 11057 28027 11115 28033
rect 11241 28067 11299 28073
rect 11241 28033 11253 28067
rect 11287 28033 11299 28067
rect 11241 28027 11299 28033
rect 6748 27968 7328 27996
rect 6641 27959 6699 27965
rect 7466 27956 7472 28008
rect 7524 27996 7530 28008
rect 7650 27996 7656 28008
rect 7524 27968 7656 27996
rect 7524 27956 7530 27968
rect 7650 27956 7656 27968
rect 7708 27956 7714 28008
rect 9493 27999 9551 28005
rect 9493 27965 9505 27999
rect 9539 27996 9551 27999
rect 9766 27996 9772 28008
rect 9539 27968 9772 27996
rect 9539 27965 9551 27968
rect 9493 27959 9551 27965
rect 9766 27956 9772 27968
rect 9824 27956 9830 28008
rect 10321 27999 10379 28005
rect 10321 27965 10333 27999
rect 10367 27996 10379 27999
rect 11256 27996 11284 28027
rect 11330 28024 11336 28076
rect 11388 28064 11394 28076
rect 11517 28067 11575 28073
rect 11517 28064 11529 28067
rect 11388 28036 11529 28064
rect 11388 28024 11394 28036
rect 11517 28033 11529 28036
rect 11563 28033 11575 28067
rect 11517 28027 11575 28033
rect 11793 28067 11851 28073
rect 11793 28033 11805 28067
rect 11839 28064 11851 28067
rect 11974 28064 11980 28076
rect 11839 28036 11980 28064
rect 11839 28033 11851 28036
rect 11793 28027 11851 28033
rect 11974 28024 11980 28036
rect 12032 28024 12038 28076
rect 11422 27996 11428 28008
rect 10367 27968 11428 27996
rect 10367 27965 10379 27968
rect 10321 27959 10379 27965
rect 11422 27956 11428 27968
rect 11480 27996 11486 28008
rect 12084 27996 12112 28172
rect 12158 28160 12164 28172
rect 12216 28160 12222 28212
rect 12894 28200 12900 28212
rect 12406 28172 12900 28200
rect 11480 27968 12112 27996
rect 11480 27956 11486 27968
rect 7098 27928 7104 27940
rect 6196 27900 7104 27928
rect 7098 27888 7104 27900
rect 7156 27888 7162 27940
rect 11330 27928 11336 27940
rect 10796 27900 11336 27928
rect 5074 27820 5080 27872
rect 5132 27860 5138 27872
rect 5442 27860 5448 27872
rect 5132 27832 5448 27860
rect 5132 27820 5138 27832
rect 5442 27820 5448 27832
rect 5500 27860 5506 27872
rect 6362 27860 6368 27872
rect 5500 27832 6368 27860
rect 5500 27820 5506 27832
rect 6362 27820 6368 27832
rect 6420 27860 6426 27872
rect 6457 27863 6515 27869
rect 6457 27860 6469 27863
rect 6420 27832 6469 27860
rect 6420 27820 6426 27832
rect 6457 27829 6469 27832
rect 6503 27829 6515 27863
rect 6457 27823 6515 27829
rect 6546 27820 6552 27872
rect 6604 27860 6610 27872
rect 10796 27869 10824 27900
rect 11330 27888 11336 27900
rect 11388 27888 11394 27940
rect 12406 27928 12434 28172
rect 12894 28160 12900 28172
rect 12952 28160 12958 28212
rect 13357 28203 13415 28209
rect 13357 28169 13369 28203
rect 13403 28200 13415 28203
rect 15010 28200 15016 28212
rect 13403 28172 15016 28200
rect 13403 28169 13415 28172
rect 13357 28163 13415 28169
rect 15010 28160 15016 28172
rect 15068 28160 15074 28212
rect 16298 28160 16304 28212
rect 16356 28200 16362 28212
rect 17037 28203 17095 28209
rect 17037 28200 17049 28203
rect 16356 28172 17049 28200
rect 16356 28160 16362 28172
rect 17037 28169 17049 28172
rect 17083 28169 17095 28203
rect 17037 28163 17095 28169
rect 17236 28172 17816 28200
rect 12989 28135 13047 28141
rect 12989 28101 13001 28135
rect 13035 28132 13047 28135
rect 13078 28132 13084 28144
rect 13035 28104 13084 28132
rect 13035 28101 13047 28104
rect 12989 28095 13047 28101
rect 13078 28092 13084 28104
rect 13136 28092 13142 28144
rect 13189 28135 13247 28141
rect 13189 28132 13201 28135
rect 13188 28101 13201 28132
rect 13235 28101 13247 28135
rect 13188 28095 13247 28101
rect 13188 28064 13216 28095
rect 14274 28092 14280 28144
rect 14332 28092 14338 28144
rect 15028 28132 15056 28160
rect 16669 28135 16727 28141
rect 15028 28104 16252 28132
rect 11992 27900 12434 27928
rect 13096 28036 13216 28064
rect 7009 27863 7067 27869
rect 7009 27860 7021 27863
rect 6604 27832 7021 27860
rect 6604 27820 6610 27832
rect 7009 27829 7021 27832
rect 7055 27829 7067 27863
rect 7009 27823 7067 27829
rect 10781 27863 10839 27869
rect 10781 27829 10793 27863
rect 10827 27829 10839 27863
rect 10781 27823 10839 27829
rect 10965 27863 11023 27869
rect 10965 27829 10977 27863
rect 11011 27860 11023 27863
rect 11992 27860 12020 27900
rect 11011 27832 12020 27860
rect 11011 27829 11023 27832
rect 10965 27823 11023 27829
rect 12066 27820 12072 27872
rect 12124 27820 12130 27872
rect 12434 27820 12440 27872
rect 12492 27860 12498 27872
rect 13096 27860 13124 28036
rect 13446 28024 13452 28076
rect 13504 28024 13510 28076
rect 16224 28073 16252 28104
rect 16669 28101 16681 28135
rect 16715 28132 16727 28135
rect 17236 28132 17264 28172
rect 16715 28104 17264 28132
rect 17788 28132 17816 28172
rect 17862 28160 17868 28212
rect 17920 28200 17926 28212
rect 20717 28203 20775 28209
rect 20717 28200 20729 28203
rect 17920 28172 20729 28200
rect 17920 28160 17926 28172
rect 20717 28169 20729 28172
rect 20763 28169 20775 28203
rect 20717 28163 20775 28169
rect 18414 28132 18420 28144
rect 17788 28104 18420 28132
rect 16715 28101 16727 28104
rect 16669 28095 16727 28101
rect 15933 28067 15991 28073
rect 15933 28033 15945 28067
rect 15979 28064 15991 28067
rect 16025 28067 16083 28073
rect 16025 28064 16037 28067
rect 15979 28036 16037 28064
rect 15979 28033 15991 28036
rect 15933 28027 15991 28033
rect 16025 28033 16037 28036
rect 16071 28033 16083 28067
rect 16025 28027 16083 28033
rect 16209 28067 16267 28073
rect 16209 28033 16221 28067
rect 16255 28033 16267 28067
rect 16209 28027 16267 28033
rect 16482 28024 16488 28076
rect 16540 28064 16546 28076
rect 16853 28067 16911 28073
rect 16853 28064 16865 28067
rect 16540 28036 16865 28064
rect 16540 28024 16546 28036
rect 16853 28033 16865 28036
rect 16899 28033 16911 28067
rect 16853 28027 16911 28033
rect 16945 28067 17003 28073
rect 16945 28033 16957 28067
rect 16991 28033 17003 28067
rect 16945 28027 17003 28033
rect 17313 28067 17371 28073
rect 17313 28033 17325 28067
rect 17359 28064 17371 28067
rect 17678 28064 17684 28076
rect 17359 28036 17684 28064
rect 17359 28033 17371 28036
rect 17313 28027 17371 28033
rect 13725 27999 13783 28005
rect 13725 27965 13737 27999
rect 13771 27996 13783 27999
rect 15381 27999 15439 28005
rect 13771 27968 14964 27996
rect 13771 27965 13783 27968
rect 13725 27959 13783 27965
rect 14936 27928 14964 27968
rect 15381 27965 15393 27999
rect 15427 27996 15439 27999
rect 15470 27996 15476 28008
rect 15427 27968 15476 27996
rect 15427 27965 15439 27968
rect 15381 27959 15439 27965
rect 15470 27956 15476 27968
rect 15528 27956 15534 28008
rect 16025 27931 16083 27937
rect 16025 27928 16037 27931
rect 13188 27900 13584 27928
rect 14936 27900 16037 27928
rect 13188 27869 13216 27900
rect 12492 27832 13124 27860
rect 13173 27863 13231 27869
rect 12492 27820 12498 27832
rect 13173 27829 13185 27863
rect 13219 27829 13231 27863
rect 13556 27860 13584 27900
rect 16025 27897 16037 27900
rect 16071 27897 16083 27931
rect 16868 27928 16896 28027
rect 16960 27996 16988 28027
rect 17678 28024 17684 28036
rect 17736 28024 17742 28076
rect 17788 28073 17816 28104
rect 18414 28092 18420 28104
rect 18472 28132 18478 28144
rect 18472 28104 18644 28132
rect 18472 28092 18478 28104
rect 17773 28067 17831 28073
rect 17773 28033 17785 28067
rect 17819 28033 17831 28067
rect 18138 28064 18144 28076
rect 17773 28027 17831 28033
rect 17880 28036 18144 28064
rect 17589 27999 17647 28005
rect 17589 27996 17601 27999
rect 16960 27968 17601 27996
rect 17589 27965 17601 27968
rect 17635 27996 17647 27999
rect 17880 27996 17908 28036
rect 18138 28024 18144 28036
rect 18196 28064 18202 28076
rect 18509 28067 18567 28073
rect 18509 28064 18521 28067
rect 18196 28036 18521 28064
rect 18196 28024 18202 28036
rect 18509 28033 18521 28036
rect 18555 28033 18567 28067
rect 18509 28027 18567 28033
rect 17635 27968 17908 27996
rect 17635 27965 17647 27968
rect 17589 27959 17647 27965
rect 18046 27956 18052 28008
rect 18104 27996 18110 28008
rect 18233 27999 18291 28005
rect 18233 27996 18245 27999
rect 18104 27968 18245 27996
rect 18104 27956 18110 27968
rect 18233 27965 18245 27968
rect 18279 27965 18291 27999
rect 18233 27959 18291 27965
rect 18322 27956 18328 28008
rect 18380 27956 18386 28008
rect 18417 27999 18475 28005
rect 18417 27965 18429 27999
rect 18463 27996 18475 27999
rect 18616 27996 18644 28104
rect 19242 28092 19248 28144
rect 19300 28132 19306 28144
rect 19300 28104 19734 28132
rect 19300 28092 19306 28104
rect 20732 28064 20760 28163
rect 21818 28160 21824 28212
rect 21876 28200 21882 28212
rect 22278 28200 22284 28212
rect 21876 28172 22284 28200
rect 21876 28160 21882 28172
rect 22278 28160 22284 28172
rect 22336 28200 22342 28212
rect 24210 28200 24216 28212
rect 22336 28172 24216 28200
rect 22336 28160 22342 28172
rect 24210 28160 24216 28172
rect 24268 28160 24274 28212
rect 24670 28160 24676 28212
rect 24728 28160 24734 28212
rect 22066 28104 22876 28132
rect 20806 28064 20812 28076
rect 20732 28036 20812 28064
rect 20806 28024 20812 28036
rect 20864 28024 20870 28076
rect 22066 28064 22094 28104
rect 21284 28036 22094 28064
rect 21284 28008 21312 28036
rect 22370 28024 22376 28076
rect 22428 28064 22434 28076
rect 22557 28067 22615 28073
rect 22557 28064 22569 28067
rect 22428 28036 22569 28064
rect 22428 28024 22434 28036
rect 22557 28033 22569 28036
rect 22603 28033 22615 28067
rect 22557 28027 22615 28033
rect 22646 28024 22652 28076
rect 22704 28024 22710 28076
rect 22848 28073 22876 28104
rect 23198 28092 23204 28144
rect 23256 28092 23262 28144
rect 23750 28092 23756 28144
rect 23808 28092 23814 28144
rect 22833 28067 22891 28073
rect 22833 28033 22845 28067
rect 22879 28033 22891 28067
rect 22833 28027 22891 28033
rect 18463 27968 18644 27996
rect 18969 27999 19027 28005
rect 18463 27965 18475 27968
rect 18417 27959 18475 27965
rect 18969 27965 18981 27999
rect 19015 27965 19027 27999
rect 18969 27959 19027 27965
rect 19245 27999 19303 28005
rect 19245 27965 19257 27999
rect 19291 27996 19303 27999
rect 19334 27996 19340 28008
rect 19291 27968 19340 27996
rect 19291 27965 19303 27968
rect 19245 27959 19303 27965
rect 18340 27928 18368 27956
rect 16868 27900 18368 27928
rect 16025 27891 16083 27897
rect 14458 27860 14464 27872
rect 13556 27832 14464 27860
rect 13173 27823 13231 27829
rect 14458 27820 14464 27832
rect 14516 27860 14522 27872
rect 15197 27863 15255 27869
rect 15197 27860 15209 27863
rect 14516 27832 15209 27860
rect 14516 27820 14522 27832
rect 15197 27829 15209 27832
rect 15243 27829 15255 27863
rect 15197 27823 15255 27829
rect 17126 27820 17132 27872
rect 17184 27860 17190 27872
rect 17788 27869 17816 27900
rect 17221 27863 17279 27869
rect 17221 27860 17233 27863
rect 17184 27832 17233 27860
rect 17184 27820 17190 27832
rect 17221 27829 17233 27832
rect 17267 27829 17279 27863
rect 17221 27823 17279 27829
rect 17773 27863 17831 27869
rect 17773 27829 17785 27863
rect 17819 27829 17831 27863
rect 17773 27823 17831 27829
rect 17954 27820 17960 27872
rect 18012 27820 18018 27872
rect 18046 27820 18052 27872
rect 18104 27820 18110 27872
rect 18984 27860 19012 27959
rect 19334 27956 19340 27968
rect 19392 27956 19398 28008
rect 21266 27956 21272 28008
rect 21324 27956 21330 28008
rect 21634 27956 21640 28008
rect 21692 27996 21698 28008
rect 21821 27999 21879 28005
rect 21821 27996 21833 27999
rect 21692 27968 21833 27996
rect 21692 27956 21698 27968
rect 21821 27965 21833 27968
rect 21867 27965 21879 27999
rect 22664 27996 22692 28024
rect 22925 27999 22983 28005
rect 22925 27996 22937 27999
rect 22664 27968 22937 27996
rect 21821 27959 21879 27965
rect 22925 27965 22937 27968
rect 22971 27965 22983 27999
rect 22925 27959 22983 27965
rect 20254 27888 20260 27940
rect 20312 27928 20318 27940
rect 21453 27931 21511 27937
rect 21453 27928 21465 27931
rect 20312 27900 21465 27928
rect 20312 27888 20318 27900
rect 21453 27897 21465 27900
rect 21499 27897 21511 27931
rect 21453 27891 21511 27897
rect 22646 27888 22652 27940
rect 22704 27888 22710 27940
rect 19886 27860 19892 27872
rect 18984 27832 19892 27860
rect 19886 27820 19892 27832
rect 19944 27820 19950 27872
rect 22186 27820 22192 27872
rect 22244 27860 22250 27872
rect 22465 27863 22523 27869
rect 22465 27860 22477 27863
rect 22244 27832 22477 27860
rect 22244 27820 22250 27832
rect 22465 27829 22477 27832
rect 22511 27829 22523 27863
rect 22465 27823 22523 27829
rect 22554 27820 22560 27872
rect 22612 27820 22618 27872
rect 1104 27770 29440 27792
rect 1104 27718 4491 27770
rect 4543 27718 4555 27770
rect 4607 27718 4619 27770
rect 4671 27718 4683 27770
rect 4735 27718 4747 27770
rect 4799 27718 11574 27770
rect 11626 27718 11638 27770
rect 11690 27718 11702 27770
rect 11754 27718 11766 27770
rect 11818 27718 11830 27770
rect 11882 27718 18657 27770
rect 18709 27718 18721 27770
rect 18773 27718 18785 27770
rect 18837 27718 18849 27770
rect 18901 27718 18913 27770
rect 18965 27718 25740 27770
rect 25792 27718 25804 27770
rect 25856 27718 25868 27770
rect 25920 27718 25932 27770
rect 25984 27718 25996 27770
rect 26048 27718 29440 27770
rect 1104 27696 29440 27718
rect 3602 27616 3608 27668
rect 3660 27656 3666 27668
rect 3660 27628 4660 27656
rect 3660 27616 3666 27628
rect 4632 27597 4660 27628
rect 9306 27616 9312 27668
rect 9364 27616 9370 27668
rect 11054 27616 11060 27668
rect 11112 27616 11118 27668
rect 11330 27616 11336 27668
rect 11388 27616 11394 27668
rect 13354 27656 13360 27668
rect 12084 27628 13360 27656
rect 4617 27591 4675 27597
rect 4617 27557 4629 27591
rect 4663 27557 4675 27591
rect 4617 27551 4675 27557
rect 7190 27548 7196 27600
rect 7248 27588 7254 27600
rect 8113 27591 8171 27597
rect 8113 27588 8125 27591
rect 7248 27560 8125 27588
rect 7248 27548 7254 27560
rect 8113 27557 8125 27560
rect 8159 27588 8171 27591
rect 11072 27588 11100 27616
rect 8159 27560 11100 27588
rect 11348 27588 11376 27616
rect 11348 27560 11744 27588
rect 8159 27557 8171 27560
rect 8113 27551 8171 27557
rect 2685 27523 2743 27529
rect 2685 27489 2697 27523
rect 2731 27520 2743 27523
rect 3142 27520 3148 27532
rect 2731 27492 3148 27520
rect 2731 27489 2743 27492
rect 2685 27483 2743 27489
rect 3142 27480 3148 27492
rect 3200 27480 3206 27532
rect 4246 27480 4252 27532
rect 4304 27520 4310 27532
rect 4801 27523 4859 27529
rect 4801 27520 4813 27523
rect 4304 27492 4813 27520
rect 4304 27480 4310 27492
rect 4801 27489 4813 27492
rect 4847 27489 4859 27523
rect 4801 27483 4859 27489
rect 4338 27412 4344 27464
rect 4396 27452 4402 27464
rect 4433 27455 4491 27461
rect 4433 27452 4445 27455
rect 4396 27424 4445 27452
rect 4396 27412 4402 27424
rect 4433 27421 4445 27424
rect 4479 27421 4491 27455
rect 4433 27415 4491 27421
rect 4709 27455 4767 27461
rect 4709 27421 4721 27455
rect 4755 27421 4767 27455
rect 4709 27415 4767 27421
rect 4893 27455 4951 27461
rect 4893 27421 4905 27455
rect 4939 27452 4951 27455
rect 5442 27452 5448 27464
rect 4939 27424 5448 27452
rect 4939 27421 4951 27424
rect 4893 27415 4951 27421
rect 1486 27344 1492 27396
rect 1544 27344 1550 27396
rect 4154 27344 4160 27396
rect 4212 27384 4218 27396
rect 4724 27384 4752 27415
rect 5442 27412 5448 27424
rect 5500 27412 5506 27464
rect 8496 27461 8524 27560
rect 11716 27529 11744 27560
rect 9401 27523 9459 27529
rect 9401 27489 9413 27523
rect 9447 27520 9459 27523
rect 10229 27523 10287 27529
rect 10229 27520 10241 27523
rect 9447 27492 10241 27520
rect 9447 27489 9459 27492
rect 9401 27483 9459 27489
rect 10229 27489 10241 27492
rect 10275 27489 10287 27523
rect 11517 27523 11575 27529
rect 11517 27520 11529 27523
rect 10229 27483 10287 27489
rect 10336 27492 11529 27520
rect 7745 27455 7803 27461
rect 7745 27421 7757 27455
rect 7791 27452 7803 27455
rect 8481 27455 8539 27461
rect 7791 27424 8432 27452
rect 7791 27421 7803 27424
rect 7745 27415 7803 27421
rect 5166 27384 5172 27396
rect 4212 27356 5172 27384
rect 4212 27344 4218 27356
rect 5166 27344 5172 27356
rect 5224 27344 5230 27396
rect 7926 27344 7932 27396
rect 7984 27344 7990 27396
rect 8404 27384 8432 27424
rect 8481 27421 8493 27455
rect 8527 27421 8539 27455
rect 8481 27415 8539 27421
rect 9125 27455 9183 27461
rect 9125 27421 9137 27455
rect 9171 27421 9183 27455
rect 9125 27415 9183 27421
rect 9677 27455 9735 27461
rect 9677 27421 9689 27455
rect 9723 27452 9735 27455
rect 9766 27452 9772 27464
rect 9723 27424 9772 27452
rect 9723 27421 9735 27424
rect 9677 27415 9735 27421
rect 9140 27384 9168 27415
rect 9766 27412 9772 27424
rect 9824 27412 9830 27464
rect 9950 27412 9956 27464
rect 10008 27452 10014 27464
rect 10336 27461 10364 27492
rect 11517 27489 11529 27492
rect 11563 27489 11575 27523
rect 11517 27483 11575 27489
rect 11701 27523 11759 27529
rect 11701 27489 11713 27523
rect 11747 27489 11759 27523
rect 12084 27520 12112 27628
rect 13354 27616 13360 27628
rect 13412 27616 13418 27668
rect 13998 27616 14004 27668
rect 14056 27616 14062 27668
rect 14458 27616 14464 27668
rect 14516 27656 14522 27668
rect 14553 27659 14611 27665
rect 14553 27656 14565 27659
rect 14516 27628 14565 27656
rect 14516 27616 14522 27628
rect 14553 27625 14565 27628
rect 14599 27625 14611 27659
rect 14553 27619 14611 27625
rect 18138 27616 18144 27668
rect 18196 27656 18202 27668
rect 18233 27659 18291 27665
rect 18233 27656 18245 27659
rect 18196 27628 18245 27656
rect 18196 27616 18202 27628
rect 18233 27625 18245 27628
rect 18279 27625 18291 27659
rect 18233 27619 18291 27625
rect 19245 27659 19303 27665
rect 19245 27625 19257 27659
rect 19291 27656 19303 27659
rect 19334 27656 19340 27668
rect 19291 27628 19340 27656
rect 19291 27625 19303 27628
rect 19245 27619 19303 27625
rect 19334 27616 19340 27628
rect 19392 27616 19398 27668
rect 20152 27659 20210 27665
rect 20152 27625 20164 27659
rect 20198 27656 20210 27659
rect 22554 27656 22560 27668
rect 20198 27628 22560 27656
rect 20198 27625 20210 27628
rect 20152 27619 20210 27625
rect 22554 27616 22560 27628
rect 22612 27616 22618 27668
rect 12161 27591 12219 27597
rect 12161 27557 12173 27591
rect 12207 27588 12219 27591
rect 13909 27591 13967 27597
rect 13909 27588 13921 27591
rect 12207 27560 12434 27588
rect 12207 27557 12219 27560
rect 12161 27551 12219 27557
rect 12406 27532 12434 27560
rect 12636 27560 13921 27588
rect 12084 27492 12204 27520
rect 12406 27492 12440 27532
rect 11701 27483 11759 27489
rect 10321 27455 10379 27461
rect 10321 27452 10333 27455
rect 10008 27424 10333 27452
rect 10008 27412 10014 27424
rect 10321 27421 10333 27424
rect 10367 27421 10379 27455
rect 10321 27415 10379 27421
rect 10505 27455 10563 27461
rect 10505 27421 10517 27455
rect 10551 27421 10563 27455
rect 10505 27415 10563 27421
rect 10413 27387 10471 27393
rect 10413 27384 10425 27387
rect 8404 27356 9076 27384
rect 9140 27356 10425 27384
rect 934 27276 940 27328
rect 992 27316 998 27328
rect 1581 27319 1639 27325
rect 1581 27316 1593 27319
rect 992 27288 1593 27316
rect 992 27276 998 27288
rect 1581 27285 1593 27288
rect 1627 27285 1639 27319
rect 1581 27279 1639 27285
rect 2774 27276 2780 27328
rect 2832 27316 2838 27328
rect 3329 27319 3387 27325
rect 3329 27316 3341 27319
rect 2832 27288 3341 27316
rect 2832 27276 2838 27288
rect 3329 27285 3341 27288
rect 3375 27285 3387 27319
rect 3329 27279 3387 27285
rect 8570 27276 8576 27328
rect 8628 27276 8634 27328
rect 8938 27276 8944 27328
rect 8996 27276 9002 27328
rect 9048 27316 9076 27356
rect 10413 27353 10425 27356
rect 10459 27353 10471 27387
rect 10520 27384 10548 27415
rect 11422 27412 11428 27464
rect 11480 27452 11486 27464
rect 11609 27455 11667 27461
rect 11609 27452 11621 27455
rect 11480 27424 11621 27452
rect 11480 27412 11486 27424
rect 11609 27421 11621 27424
rect 11655 27421 11667 27455
rect 11609 27415 11667 27421
rect 11793 27455 11851 27461
rect 11793 27421 11805 27455
rect 11839 27452 11851 27455
rect 11882 27452 11888 27464
rect 11839 27424 11888 27452
rect 11839 27421 11851 27424
rect 11793 27415 11851 27421
rect 11882 27412 11888 27424
rect 11940 27412 11946 27464
rect 11977 27455 12035 27461
rect 11977 27421 11989 27455
rect 12023 27452 12035 27455
rect 12066 27452 12072 27464
rect 12023 27424 12072 27452
rect 12023 27421 12035 27424
rect 11977 27415 12035 27421
rect 12066 27412 12072 27424
rect 12124 27412 12130 27464
rect 11514 27384 11520 27396
rect 10520 27356 11520 27384
rect 10413 27347 10471 27353
rect 11514 27344 11520 27356
rect 11572 27384 11578 27396
rect 12176 27384 12204 27492
rect 12434 27480 12440 27492
rect 12492 27520 12498 27532
rect 12529 27523 12587 27529
rect 12529 27520 12541 27523
rect 12492 27492 12541 27520
rect 12492 27480 12498 27492
rect 12529 27489 12541 27492
rect 12575 27489 12587 27523
rect 12529 27483 12587 27489
rect 12636 27461 12664 27560
rect 13909 27557 13921 27560
rect 13955 27557 13967 27591
rect 14016 27588 14044 27616
rect 14829 27591 14887 27597
rect 14829 27588 14841 27591
rect 14016 27560 14841 27588
rect 13909 27551 13967 27557
rect 14829 27557 14841 27560
rect 14875 27557 14887 27591
rect 14829 27551 14887 27557
rect 21729 27591 21787 27597
rect 21729 27557 21741 27591
rect 21775 27588 21787 27591
rect 22646 27588 22652 27600
rect 21775 27560 22652 27588
rect 21775 27557 21787 27560
rect 21729 27551 21787 27557
rect 22646 27548 22652 27560
rect 22704 27548 22710 27600
rect 22830 27548 22836 27600
rect 22888 27548 22894 27600
rect 12989 27523 13047 27529
rect 12989 27520 13001 27523
rect 12820 27492 13001 27520
rect 12820 27464 12848 27492
rect 12989 27489 13001 27492
rect 13035 27489 13047 27523
rect 12989 27483 13047 27489
rect 13078 27480 13084 27532
rect 13136 27520 13142 27532
rect 13265 27523 13323 27529
rect 13265 27520 13277 27523
rect 13136 27492 13277 27520
rect 13136 27480 13142 27492
rect 13265 27489 13277 27492
rect 13311 27520 13323 27523
rect 13998 27520 14004 27532
rect 13311 27492 14004 27520
rect 13311 27489 13323 27492
rect 13265 27483 13323 27489
rect 13998 27480 14004 27492
rect 14056 27480 14062 27532
rect 14185 27523 14243 27529
rect 14185 27489 14197 27523
rect 14231 27520 14243 27523
rect 15562 27520 15568 27532
rect 14231 27492 15568 27520
rect 14231 27489 14243 27492
rect 14185 27483 14243 27489
rect 15562 27480 15568 27492
rect 15620 27480 15626 27532
rect 16482 27480 16488 27532
rect 16540 27480 16546 27532
rect 17126 27480 17132 27532
rect 17184 27520 17190 27532
rect 17184 27492 19656 27520
rect 17184 27480 17190 27492
rect 12621 27455 12679 27461
rect 12621 27421 12633 27455
rect 12667 27421 12679 27455
rect 12621 27415 12679 27421
rect 12802 27412 12808 27464
rect 12860 27412 12866 27464
rect 14277 27455 14335 27461
rect 14277 27452 14289 27455
rect 13372 27424 14289 27452
rect 11572 27356 12204 27384
rect 11572 27344 11578 27356
rect 10778 27316 10784 27328
rect 9048 27288 10784 27316
rect 10778 27276 10784 27288
rect 10836 27276 10842 27328
rect 11333 27319 11391 27325
rect 11333 27285 11345 27319
rect 11379 27316 11391 27319
rect 11882 27316 11888 27328
rect 11379 27288 11888 27316
rect 11379 27285 11391 27288
rect 11333 27279 11391 27285
rect 11882 27276 11888 27288
rect 11940 27276 11946 27328
rect 11974 27276 11980 27328
rect 12032 27316 12038 27328
rect 12526 27316 12532 27328
rect 12032 27288 12532 27316
rect 12032 27276 12038 27288
rect 12526 27276 12532 27288
rect 12584 27316 12590 27328
rect 13372 27316 13400 27424
rect 14277 27421 14289 27424
rect 14323 27421 14335 27455
rect 14277 27415 14335 27421
rect 14645 27455 14703 27461
rect 14645 27421 14657 27455
rect 14691 27421 14703 27455
rect 14645 27415 14703 27421
rect 12584 27288 13400 27316
rect 12584 27276 12590 27288
rect 13998 27276 14004 27328
rect 14056 27316 14062 27328
rect 14458 27316 14464 27328
rect 14056 27288 14464 27316
rect 14056 27276 14062 27288
rect 14458 27276 14464 27288
rect 14516 27316 14522 27328
rect 14660 27316 14688 27415
rect 16390 27412 16396 27464
rect 16448 27412 16454 27464
rect 19245 27455 19303 27461
rect 19245 27421 19257 27455
rect 19291 27452 19303 27455
rect 19426 27452 19432 27464
rect 19291 27424 19432 27452
rect 19291 27421 19303 27424
rect 19245 27415 19303 27421
rect 19426 27412 19432 27424
rect 19484 27412 19490 27464
rect 19518 27412 19524 27464
rect 19576 27452 19582 27464
rect 19628 27452 19656 27492
rect 20806 27480 20812 27532
rect 20864 27520 20870 27532
rect 20864 27492 21956 27520
rect 20864 27480 20870 27492
rect 19576 27424 19656 27452
rect 19576 27412 19582 27424
rect 19886 27412 19892 27464
rect 19944 27412 19950 27464
rect 21928 27461 21956 27492
rect 22094 27480 22100 27532
rect 22152 27520 22158 27532
rect 22557 27523 22615 27529
rect 22557 27520 22569 27523
rect 22152 27492 22569 27520
rect 22152 27480 22158 27492
rect 22557 27489 22569 27492
rect 22603 27489 22615 27523
rect 22557 27483 22615 27489
rect 22741 27523 22799 27529
rect 22741 27489 22753 27523
rect 22787 27520 22799 27523
rect 22848 27520 22876 27548
rect 22787 27492 22876 27520
rect 22787 27489 22799 27492
rect 22741 27483 22799 27489
rect 21913 27455 21971 27461
rect 21913 27421 21925 27455
rect 21959 27421 21971 27455
rect 21913 27415 21971 27421
rect 22002 27412 22008 27464
rect 22060 27412 22066 27464
rect 22278 27412 22284 27464
rect 22336 27412 22342 27464
rect 22370 27412 22376 27464
rect 22428 27452 22434 27464
rect 22649 27455 22707 27461
rect 22649 27452 22661 27455
rect 22428 27424 22661 27452
rect 22428 27412 22434 27424
rect 22649 27421 22661 27424
rect 22695 27421 22707 27455
rect 22649 27415 22707 27421
rect 22833 27455 22891 27461
rect 22833 27421 22845 27455
rect 22879 27452 22891 27455
rect 24394 27452 24400 27464
rect 22879 27424 24400 27452
rect 22879 27421 22891 27424
rect 22833 27415 22891 27421
rect 24394 27412 24400 27424
rect 24452 27412 24458 27464
rect 16761 27387 16819 27393
rect 16761 27353 16773 27387
rect 16807 27353 16819 27387
rect 16761 27347 16819 27353
rect 14516 27288 14688 27316
rect 16209 27319 16267 27325
rect 14516 27276 14522 27288
rect 16209 27285 16221 27319
rect 16255 27316 16267 27319
rect 16776 27316 16804 27347
rect 17218 27344 17224 27396
rect 17276 27344 17282 27396
rect 19904 27384 19932 27412
rect 20070 27384 20076 27396
rect 19904 27356 20076 27384
rect 20070 27344 20076 27356
rect 20128 27344 20134 27396
rect 20254 27344 20260 27396
rect 20312 27344 20318 27396
rect 20714 27344 20720 27396
rect 20772 27344 20778 27396
rect 21729 27387 21787 27393
rect 21729 27353 21741 27387
rect 21775 27384 21787 27387
rect 22186 27384 22192 27396
rect 21775 27356 22192 27384
rect 21775 27353 21787 27356
rect 21729 27347 21787 27353
rect 22186 27344 22192 27356
rect 22244 27344 22250 27396
rect 16255 27288 16804 27316
rect 19429 27319 19487 27325
rect 16255 27285 16267 27288
rect 16209 27279 16267 27285
rect 19429 27285 19441 27319
rect 19475 27316 19487 27319
rect 20272 27316 20300 27344
rect 19475 27288 20300 27316
rect 19475 27285 19487 27288
rect 19429 27279 19487 27285
rect 20990 27276 20996 27328
rect 21048 27316 21054 27328
rect 21634 27316 21640 27328
rect 21048 27288 21640 27316
rect 21048 27276 21054 27288
rect 21634 27276 21640 27288
rect 21692 27276 21698 27328
rect 22002 27276 22008 27328
rect 22060 27316 22066 27328
rect 22388 27316 22416 27412
rect 22060 27288 22416 27316
rect 22060 27276 22066 27288
rect 1104 27226 29595 27248
rect 1104 27174 8032 27226
rect 8084 27174 8096 27226
rect 8148 27174 8160 27226
rect 8212 27174 8224 27226
rect 8276 27174 8288 27226
rect 8340 27174 15115 27226
rect 15167 27174 15179 27226
rect 15231 27174 15243 27226
rect 15295 27174 15307 27226
rect 15359 27174 15371 27226
rect 15423 27174 22198 27226
rect 22250 27174 22262 27226
rect 22314 27174 22326 27226
rect 22378 27174 22390 27226
rect 22442 27174 22454 27226
rect 22506 27174 29281 27226
rect 29333 27174 29345 27226
rect 29397 27174 29409 27226
rect 29461 27174 29473 27226
rect 29525 27174 29537 27226
rect 29589 27174 29595 27226
rect 1104 27152 29595 27174
rect 8938 27112 8944 27124
rect 8220 27084 8944 27112
rect 8220 27053 8248 27084
rect 8938 27072 8944 27084
rect 8996 27072 9002 27124
rect 9677 27115 9735 27121
rect 9677 27081 9689 27115
rect 9723 27112 9735 27115
rect 9766 27112 9772 27124
rect 9723 27084 9772 27112
rect 9723 27081 9735 27084
rect 9677 27075 9735 27081
rect 9766 27072 9772 27084
rect 9824 27072 9830 27124
rect 10778 27072 10784 27124
rect 10836 27112 10842 27124
rect 13630 27112 13636 27124
rect 10836 27084 13636 27112
rect 10836 27072 10842 27084
rect 13630 27072 13636 27084
rect 13688 27072 13694 27124
rect 14277 27115 14335 27121
rect 14277 27081 14289 27115
rect 14323 27112 14335 27115
rect 14458 27112 14464 27124
rect 14323 27084 14464 27112
rect 14323 27081 14335 27084
rect 14277 27075 14335 27081
rect 14458 27072 14464 27084
rect 14516 27112 14522 27124
rect 14553 27115 14611 27121
rect 14553 27112 14565 27115
rect 14516 27084 14565 27112
rect 14516 27072 14522 27084
rect 14553 27081 14565 27084
rect 14599 27081 14611 27115
rect 14553 27075 14611 27081
rect 16390 27072 16396 27124
rect 16448 27112 16454 27124
rect 17589 27115 17647 27121
rect 17589 27112 17601 27115
rect 16448 27084 17601 27112
rect 16448 27072 16454 27084
rect 17589 27081 17601 27084
rect 17635 27081 17647 27115
rect 17589 27075 17647 27081
rect 19518 27072 19524 27124
rect 19576 27072 19582 27124
rect 20898 27072 20904 27124
rect 20956 27112 20962 27124
rect 21177 27115 21235 27121
rect 21177 27112 21189 27115
rect 20956 27084 21189 27112
rect 20956 27072 20962 27084
rect 21177 27081 21189 27084
rect 21223 27112 21235 27115
rect 22002 27112 22008 27124
rect 21223 27084 22008 27112
rect 21223 27081 21235 27084
rect 21177 27075 21235 27081
rect 22002 27072 22008 27084
rect 22060 27072 22066 27124
rect 8205 27047 8263 27053
rect 8205 27013 8217 27047
rect 8251 27013 8263 27047
rect 8205 27007 8263 27013
rect 11146 27004 11152 27056
rect 11204 27044 11210 27056
rect 12710 27044 12716 27056
rect 11204 27016 12716 27044
rect 11204 27004 11210 27016
rect 12710 27004 12716 27016
rect 12768 27004 12774 27056
rect 12802 27004 12808 27056
rect 12860 27004 12866 27056
rect 14369 27047 14427 27053
rect 14369 27013 14381 27047
rect 14415 27044 14427 27047
rect 14734 27044 14740 27056
rect 14415 27016 14740 27044
rect 14415 27013 14427 27016
rect 14369 27007 14427 27013
rect 14734 27004 14740 27016
rect 14792 27004 14798 27056
rect 17126 27004 17132 27056
rect 17184 27004 17190 27056
rect 9214 26936 9220 26988
rect 9272 26976 9278 26988
rect 11793 26979 11851 26985
rect 11793 26976 11805 26979
rect 9272 26948 9338 26976
rect 11624 26948 11805 26976
rect 9272 26936 9278 26948
rect 7650 26868 7656 26920
rect 7708 26908 7714 26920
rect 7929 26911 7987 26917
rect 7929 26908 7941 26911
rect 7708 26880 7941 26908
rect 7708 26868 7714 26880
rect 7929 26877 7941 26880
rect 7975 26877 7987 26911
rect 7929 26871 7987 26877
rect 8570 26868 8576 26920
rect 8628 26908 8634 26920
rect 8628 26880 9260 26908
rect 8628 26868 8634 26880
rect 9232 26840 9260 26880
rect 11514 26868 11520 26920
rect 11572 26908 11578 26920
rect 11624 26908 11652 26948
rect 11793 26945 11805 26948
rect 11839 26945 11851 26979
rect 11793 26939 11851 26945
rect 12250 26936 12256 26988
rect 12308 26976 12314 26988
rect 12529 26979 12587 26985
rect 12529 26976 12541 26979
rect 12308 26948 12541 26976
rect 12308 26936 12314 26948
rect 12529 26945 12541 26948
rect 12575 26945 12587 26979
rect 12529 26939 12587 26945
rect 13906 26936 13912 26988
rect 13964 26936 13970 26988
rect 14645 26979 14703 26985
rect 14645 26976 14657 26979
rect 14016 26948 14657 26976
rect 11572 26880 11652 26908
rect 11708 26911 11766 26917
rect 11572 26868 11578 26880
rect 11708 26877 11720 26911
rect 11754 26877 11766 26911
rect 11708 26871 11766 26877
rect 11532 26840 11560 26868
rect 9232 26812 11560 26840
rect 11716 26840 11744 26871
rect 11882 26868 11888 26920
rect 11940 26868 11946 26920
rect 12434 26908 12440 26920
rect 11992 26880 12440 26908
rect 11992 26840 12020 26880
rect 12434 26868 12440 26880
rect 12492 26908 12498 26920
rect 14016 26908 14044 26948
rect 14645 26945 14657 26948
rect 14691 26945 14703 26979
rect 19536 26976 19564 27072
rect 20806 27004 20812 27056
rect 20864 27004 20870 27056
rect 21039 27013 21097 27019
rect 21039 27010 21051 27013
rect 21024 26979 21051 27010
rect 21085 26979 21097 27013
rect 21024 26976 21097 26979
rect 21910 26976 21916 26988
rect 19536 26948 21916 26976
rect 14645 26939 14703 26945
rect 21910 26936 21916 26948
rect 21968 26936 21974 26988
rect 28258 26936 28264 26988
rect 28316 26976 28322 26988
rect 28813 26979 28871 26985
rect 28813 26976 28825 26979
rect 28316 26948 28825 26976
rect 28316 26936 28322 26948
rect 28813 26945 28825 26948
rect 28859 26945 28871 26979
rect 28813 26939 28871 26945
rect 15470 26908 15476 26920
rect 12492 26880 14044 26908
rect 14384 26880 15476 26908
rect 12492 26868 12498 26880
rect 11716 26812 12020 26840
rect 13906 26800 13912 26852
rect 13964 26840 13970 26852
rect 14274 26840 14280 26852
rect 13964 26812 14280 26840
rect 13964 26800 13970 26812
rect 14274 26800 14280 26812
rect 14332 26800 14338 26852
rect 14384 26849 14412 26880
rect 15470 26868 15476 26880
rect 15528 26868 15534 26920
rect 14369 26843 14427 26849
rect 14369 26809 14381 26843
rect 14415 26809 14427 26843
rect 14369 26803 14427 26809
rect 17497 26843 17555 26849
rect 17497 26809 17509 26843
rect 17543 26840 17555 26843
rect 18046 26840 18052 26852
rect 17543 26812 18052 26840
rect 17543 26809 17555 26812
rect 17497 26803 17555 26809
rect 18046 26800 18052 26812
rect 18104 26800 18110 26852
rect 11238 26732 11244 26784
rect 11296 26772 11302 26784
rect 11517 26775 11575 26781
rect 11517 26772 11529 26775
rect 11296 26744 11529 26772
rect 11296 26732 11302 26744
rect 11517 26741 11529 26744
rect 11563 26741 11575 26775
rect 11517 26735 11575 26741
rect 12802 26732 12808 26784
rect 12860 26772 12866 26784
rect 13924 26772 13952 26800
rect 12860 26744 13952 26772
rect 12860 26732 12866 26744
rect 20990 26732 20996 26784
rect 21048 26732 21054 26784
rect 28994 26732 29000 26784
rect 29052 26732 29058 26784
rect 1104 26682 29440 26704
rect 1104 26630 4491 26682
rect 4543 26630 4555 26682
rect 4607 26630 4619 26682
rect 4671 26630 4683 26682
rect 4735 26630 4747 26682
rect 4799 26630 11574 26682
rect 11626 26630 11638 26682
rect 11690 26630 11702 26682
rect 11754 26630 11766 26682
rect 11818 26630 11830 26682
rect 11882 26630 18657 26682
rect 18709 26630 18721 26682
rect 18773 26630 18785 26682
rect 18837 26630 18849 26682
rect 18901 26630 18913 26682
rect 18965 26630 25740 26682
rect 25792 26630 25804 26682
rect 25856 26630 25868 26682
rect 25920 26630 25932 26682
rect 25984 26630 25996 26682
rect 26048 26630 29440 26682
rect 1104 26608 29440 26630
rect 1486 26528 1492 26580
rect 1544 26568 1550 26580
rect 2225 26571 2283 26577
rect 2225 26568 2237 26571
rect 1544 26540 2237 26568
rect 1544 26528 1550 26540
rect 2225 26537 2237 26540
rect 2271 26537 2283 26571
rect 2225 26531 2283 26537
rect 11044 26571 11102 26577
rect 11044 26537 11056 26571
rect 11090 26568 11102 26571
rect 11238 26568 11244 26580
rect 11090 26540 11244 26568
rect 11090 26537 11102 26540
rect 11044 26531 11102 26537
rect 11238 26528 11244 26540
rect 11296 26528 11302 26580
rect 12526 26528 12532 26580
rect 12584 26528 12590 26580
rect 7006 26432 7012 26444
rect 5736 26404 7012 26432
rect 2406 26324 2412 26376
rect 2464 26324 2470 26376
rect 5736 26373 5764 26404
rect 7006 26392 7012 26404
rect 7064 26392 7070 26444
rect 10410 26392 10416 26444
rect 10468 26432 10474 26444
rect 10781 26435 10839 26441
rect 10781 26432 10793 26435
rect 10468 26404 10793 26432
rect 10468 26392 10474 26404
rect 10781 26401 10793 26404
rect 10827 26432 10839 26435
rect 11422 26432 11428 26444
rect 10827 26404 11428 26432
rect 10827 26401 10839 26404
rect 10781 26395 10839 26401
rect 11422 26392 11428 26404
rect 11480 26432 11486 26444
rect 12250 26432 12256 26444
rect 11480 26404 12256 26432
rect 11480 26392 11486 26404
rect 12250 26392 12256 26404
rect 12308 26392 12314 26444
rect 5721 26367 5779 26373
rect 5721 26333 5733 26367
rect 5767 26333 5779 26367
rect 5721 26327 5779 26333
rect 5905 26367 5963 26373
rect 5905 26333 5917 26367
rect 5951 26333 5963 26367
rect 5905 26327 5963 26333
rect 5920 26296 5948 26327
rect 6270 26324 6276 26376
rect 6328 26324 6334 26376
rect 9214 26324 9220 26376
rect 9272 26324 9278 26376
rect 17954 26324 17960 26376
rect 18012 26364 18018 26376
rect 19613 26367 19671 26373
rect 19613 26364 19625 26367
rect 18012 26336 19625 26364
rect 18012 26324 18018 26336
rect 19613 26333 19625 26336
rect 19659 26333 19671 26367
rect 19613 26327 19671 26333
rect 6825 26299 6883 26305
rect 6825 26296 6837 26299
rect 5920 26268 6837 26296
rect 6825 26265 6837 26268
rect 6871 26265 6883 26299
rect 9232 26296 9260 26324
rect 11146 26296 11152 26308
rect 9232 26268 11152 26296
rect 6825 26259 6883 26265
rect 11146 26256 11152 26268
rect 11204 26296 11210 26308
rect 19245 26299 19303 26305
rect 11204 26268 11546 26296
rect 11204 26256 11210 26268
rect 19245 26265 19257 26299
rect 19291 26265 19303 26299
rect 19245 26259 19303 26265
rect 5810 26188 5816 26240
rect 5868 26188 5874 26240
rect 19260 26228 19288 26259
rect 19426 26256 19432 26308
rect 19484 26256 19490 26308
rect 19794 26256 19800 26308
rect 19852 26256 19858 26308
rect 19812 26228 19840 26256
rect 19260 26200 19840 26228
rect 1104 26138 29595 26160
rect 1104 26086 8032 26138
rect 8084 26086 8096 26138
rect 8148 26086 8160 26138
rect 8212 26086 8224 26138
rect 8276 26086 8288 26138
rect 8340 26086 15115 26138
rect 15167 26086 15179 26138
rect 15231 26086 15243 26138
rect 15295 26086 15307 26138
rect 15359 26086 15371 26138
rect 15423 26086 22198 26138
rect 22250 26086 22262 26138
rect 22314 26086 22326 26138
rect 22378 26086 22390 26138
rect 22442 26086 22454 26138
rect 22506 26086 29281 26138
rect 29333 26086 29345 26138
rect 29397 26086 29409 26138
rect 29461 26086 29473 26138
rect 29525 26086 29537 26138
rect 29589 26086 29595 26138
rect 1104 26064 29595 26086
rect 6181 26027 6239 26033
rect 6181 25993 6193 26027
rect 6227 26024 6239 26027
rect 7926 26024 7932 26036
rect 6227 25996 7932 26024
rect 6227 25993 6239 25996
rect 6181 25987 6239 25993
rect 7926 25984 7932 25996
rect 7984 25984 7990 26036
rect 20714 26024 20720 26036
rect 19444 25996 20720 26024
rect 5810 25956 5816 25968
rect 5000 25928 5816 25956
rect 5000 25897 5028 25928
rect 5810 25916 5816 25928
rect 5868 25916 5874 25968
rect 6454 25956 6460 25968
rect 6012 25928 6460 25956
rect 4985 25891 5043 25897
rect 4985 25857 4997 25891
rect 5031 25857 5043 25891
rect 4985 25851 5043 25857
rect 5166 25848 5172 25900
rect 5224 25848 5230 25900
rect 5261 25891 5319 25897
rect 5261 25857 5273 25891
rect 5307 25857 5319 25891
rect 5261 25851 5319 25857
rect 5276 25820 5304 25851
rect 5350 25848 5356 25900
rect 5408 25888 5414 25900
rect 6012 25897 6040 25928
rect 6454 25916 6460 25928
rect 6512 25916 6518 25968
rect 8570 25956 8576 25968
rect 8220 25928 8576 25956
rect 5445 25891 5503 25897
rect 5445 25888 5457 25891
rect 5408 25860 5457 25888
rect 5408 25848 5414 25860
rect 5445 25857 5457 25860
rect 5491 25857 5503 25891
rect 5721 25891 5779 25897
rect 5721 25888 5733 25891
rect 5445 25851 5503 25857
rect 5644 25860 5733 25888
rect 5534 25820 5540 25832
rect 4356 25792 5540 25820
rect 4356 25696 4384 25792
rect 5534 25780 5540 25792
rect 5592 25780 5598 25832
rect 5644 25696 5672 25860
rect 5721 25857 5733 25860
rect 5767 25857 5779 25891
rect 5721 25851 5779 25857
rect 5997 25891 6055 25897
rect 5997 25857 6009 25891
rect 6043 25857 6055 25891
rect 6546 25888 6552 25900
rect 5997 25851 6055 25857
rect 6104 25860 6552 25888
rect 5905 25823 5963 25829
rect 5905 25789 5917 25823
rect 5951 25820 5963 25823
rect 6104 25820 6132 25860
rect 6546 25848 6552 25860
rect 6604 25848 6610 25900
rect 6914 25848 6920 25900
rect 6972 25888 6978 25900
rect 7101 25891 7159 25897
rect 7101 25888 7113 25891
rect 6972 25860 7113 25888
rect 6972 25848 6978 25860
rect 7101 25857 7113 25860
rect 7147 25857 7159 25891
rect 7101 25851 7159 25857
rect 7282 25848 7288 25900
rect 7340 25848 7346 25900
rect 8220 25897 8248 25928
rect 8570 25916 8576 25928
rect 8628 25916 8634 25968
rect 18230 25916 18236 25968
rect 18288 25956 18294 25968
rect 19061 25959 19119 25965
rect 19061 25956 19073 25959
rect 18288 25928 19073 25956
rect 18288 25916 18294 25928
rect 19061 25925 19073 25928
rect 19107 25925 19119 25959
rect 19061 25919 19119 25925
rect 19334 25916 19340 25968
rect 19392 25956 19398 25968
rect 19444 25956 19472 25996
rect 20714 25984 20720 25996
rect 20772 25984 20778 26036
rect 19392 25928 19550 25956
rect 19392 25916 19398 25928
rect 7377 25891 7435 25897
rect 7377 25857 7389 25891
rect 7423 25888 7435 25891
rect 8113 25891 8171 25897
rect 8113 25888 8125 25891
rect 7423 25860 8125 25888
rect 7423 25857 7435 25860
rect 7377 25851 7435 25857
rect 8113 25857 8125 25860
rect 8159 25857 8171 25891
rect 8113 25851 8171 25857
rect 8205 25891 8263 25897
rect 8205 25857 8217 25891
rect 8251 25857 8263 25891
rect 8205 25851 8263 25857
rect 8389 25891 8447 25897
rect 8389 25857 8401 25891
rect 8435 25857 8447 25891
rect 8389 25851 8447 25857
rect 5951 25792 6132 25820
rect 6457 25823 6515 25829
rect 5951 25789 5963 25792
rect 5905 25783 5963 25789
rect 6457 25789 6469 25823
rect 6503 25789 6515 25823
rect 6457 25783 6515 25789
rect 6472 25752 6500 25783
rect 6730 25780 6736 25832
rect 6788 25820 6794 25832
rect 7561 25823 7619 25829
rect 7561 25820 7573 25823
rect 6788 25792 7573 25820
rect 6788 25780 6794 25792
rect 7561 25789 7573 25792
rect 7607 25820 7619 25823
rect 8128 25820 8156 25851
rect 8404 25820 8432 25851
rect 7607 25792 7696 25820
rect 8128 25792 8432 25820
rect 7607 25789 7619 25792
rect 7561 25783 7619 25789
rect 7101 25755 7159 25761
rect 7101 25752 7113 25755
rect 6472 25724 7113 25752
rect 7101 25721 7113 25724
rect 7147 25721 7159 25755
rect 7101 25715 7159 25721
rect 4338 25644 4344 25696
rect 4396 25644 4402 25696
rect 4985 25687 5043 25693
rect 4985 25653 4997 25687
rect 5031 25684 5043 25687
rect 5074 25684 5080 25696
rect 5031 25656 5080 25684
rect 5031 25653 5043 25656
rect 4985 25647 5043 25653
rect 5074 25644 5080 25656
rect 5132 25644 5138 25696
rect 5626 25644 5632 25696
rect 5684 25644 5690 25696
rect 5718 25644 5724 25696
rect 5776 25644 5782 25696
rect 7009 25687 7067 25693
rect 7009 25653 7021 25687
rect 7055 25684 7067 25687
rect 7190 25684 7196 25696
rect 7055 25656 7196 25684
rect 7055 25653 7067 25656
rect 7009 25647 7067 25653
rect 7190 25644 7196 25656
rect 7248 25644 7254 25696
rect 7668 25684 7696 25792
rect 17862 25780 17868 25832
rect 17920 25820 17926 25832
rect 18785 25823 18843 25829
rect 18785 25820 18797 25823
rect 17920 25792 18797 25820
rect 17920 25780 17926 25792
rect 18785 25789 18797 25792
rect 18831 25789 18843 25823
rect 18785 25783 18843 25789
rect 7742 25712 7748 25764
rect 7800 25752 7806 25764
rect 8205 25755 8263 25761
rect 8205 25752 8217 25755
rect 7800 25724 8217 25752
rect 7800 25712 7806 25724
rect 8205 25721 8217 25724
rect 8251 25721 8263 25755
rect 8205 25715 8263 25721
rect 8754 25684 8760 25696
rect 7668 25656 8760 25684
rect 8754 25644 8760 25656
rect 8812 25644 8818 25696
rect 20533 25687 20591 25693
rect 20533 25653 20545 25687
rect 20579 25684 20591 25687
rect 20714 25684 20720 25696
rect 20579 25656 20720 25684
rect 20579 25653 20591 25656
rect 20533 25647 20591 25653
rect 20714 25644 20720 25656
rect 20772 25644 20778 25696
rect 1104 25594 29440 25616
rect 1104 25542 4491 25594
rect 4543 25542 4555 25594
rect 4607 25542 4619 25594
rect 4671 25542 4683 25594
rect 4735 25542 4747 25594
rect 4799 25542 11574 25594
rect 11626 25542 11638 25594
rect 11690 25542 11702 25594
rect 11754 25542 11766 25594
rect 11818 25542 11830 25594
rect 11882 25542 18657 25594
rect 18709 25542 18721 25594
rect 18773 25542 18785 25594
rect 18837 25542 18849 25594
rect 18901 25542 18913 25594
rect 18965 25542 25740 25594
rect 25792 25542 25804 25594
rect 25856 25542 25868 25594
rect 25920 25542 25932 25594
rect 25984 25542 25996 25594
rect 26048 25542 29440 25594
rect 1104 25520 29440 25542
rect 4972 25483 5030 25489
rect 4972 25449 4984 25483
rect 5018 25480 5030 25483
rect 5074 25480 5080 25492
rect 5018 25452 5080 25480
rect 5018 25449 5030 25452
rect 4972 25443 5030 25449
rect 5074 25440 5080 25452
rect 5132 25440 5138 25492
rect 5534 25440 5540 25492
rect 5592 25480 5598 25492
rect 5592 25452 6408 25480
rect 5592 25440 5598 25452
rect 6380 25412 6408 25452
rect 6454 25440 6460 25492
rect 6512 25440 6518 25492
rect 6730 25440 6736 25492
rect 6788 25440 6794 25492
rect 6917 25483 6975 25489
rect 6917 25449 6929 25483
rect 6963 25480 6975 25483
rect 7006 25480 7012 25492
rect 6963 25452 7012 25480
rect 6963 25449 6975 25452
rect 6917 25443 6975 25449
rect 7006 25440 7012 25452
rect 7064 25440 7070 25492
rect 7272 25483 7330 25489
rect 7272 25449 7284 25483
rect 7318 25480 7330 25483
rect 7742 25480 7748 25492
rect 7318 25452 7748 25480
rect 7318 25449 7330 25452
rect 7272 25443 7330 25449
rect 7742 25440 7748 25452
rect 7800 25440 7806 25492
rect 8754 25440 8760 25492
rect 8812 25440 8818 25492
rect 18874 25480 18880 25492
rect 18156 25452 18880 25480
rect 6748 25412 6776 25440
rect 18156 25424 18184 25452
rect 18874 25440 18880 25452
rect 18932 25440 18938 25492
rect 6380 25384 6776 25412
rect 18138 25372 18144 25424
rect 18196 25372 18202 25424
rect 18616 25384 19932 25412
rect 1857 25347 1915 25353
rect 1857 25313 1869 25347
rect 1903 25344 1915 25347
rect 4709 25347 4767 25353
rect 4709 25344 4721 25347
rect 1903 25316 4721 25344
rect 1903 25313 1915 25316
rect 1857 25307 1915 25313
rect 4709 25313 4721 25316
rect 4755 25344 4767 25347
rect 4982 25344 4988 25356
rect 4755 25316 4988 25344
rect 4755 25313 4767 25316
rect 4709 25307 4767 25313
rect 4982 25304 4988 25316
rect 5040 25304 5046 25356
rect 5350 25304 5356 25356
rect 5408 25344 5414 25356
rect 7009 25347 7067 25353
rect 5408 25316 6776 25344
rect 5408 25304 5414 25316
rect 4338 25236 4344 25288
rect 4396 25276 4402 25288
rect 4433 25279 4491 25285
rect 4433 25276 4445 25279
rect 4396 25248 4445 25276
rect 4396 25236 4402 25248
rect 4433 25245 4445 25248
rect 4479 25245 4491 25279
rect 4433 25239 4491 25245
rect 4614 25236 4620 25288
rect 4672 25236 4678 25288
rect 2133 25211 2191 25217
rect 2133 25177 2145 25211
rect 2179 25177 2191 25211
rect 3510 25208 3516 25220
rect 3358 25180 3516 25208
rect 2133 25171 2191 25177
rect 2148 25140 2176 25171
rect 3510 25168 3516 25180
rect 3568 25168 3574 25220
rect 5258 25208 5264 25220
rect 3620 25180 5264 25208
rect 2774 25140 2780 25152
rect 2148 25112 2780 25140
rect 2774 25100 2780 25112
rect 2832 25100 2838 25152
rect 3620 25149 3648 25180
rect 5258 25168 5264 25180
rect 5316 25168 5322 25220
rect 6549 25211 6607 25217
rect 5368 25180 5474 25208
rect 3605 25143 3663 25149
rect 3605 25109 3617 25143
rect 3651 25109 3663 25143
rect 3605 25103 3663 25109
rect 4617 25143 4675 25149
rect 4617 25109 4629 25143
rect 4663 25140 4675 25143
rect 4890 25140 4896 25152
rect 4663 25112 4896 25140
rect 4663 25109 4675 25112
rect 4617 25103 4675 25109
rect 4890 25100 4896 25112
rect 4948 25100 4954 25152
rect 5074 25100 5080 25152
rect 5132 25140 5138 25152
rect 5368 25140 5396 25180
rect 6549 25177 6561 25211
rect 6595 25208 6607 25211
rect 6748 25208 6776 25316
rect 7009 25313 7021 25347
rect 7055 25344 7067 25347
rect 17218 25344 17224 25356
rect 7055 25316 9352 25344
rect 7055 25313 7067 25316
rect 7009 25307 7067 25313
rect 9324 25288 9352 25316
rect 16408 25316 17224 25344
rect 8386 25236 8392 25288
rect 8444 25236 8450 25288
rect 9306 25236 9312 25288
rect 9364 25236 9370 25288
rect 12069 25279 12127 25285
rect 12069 25245 12081 25279
rect 12115 25276 12127 25279
rect 12986 25276 12992 25288
rect 12115 25248 12992 25276
rect 12115 25245 12127 25248
rect 12069 25239 12127 25245
rect 12986 25236 12992 25248
rect 13044 25236 13050 25288
rect 13446 25236 13452 25288
rect 13504 25276 13510 25288
rect 15010 25276 15016 25288
rect 13504 25248 15016 25276
rect 13504 25236 13510 25248
rect 15010 25236 15016 25248
rect 15068 25236 15074 25288
rect 16408 25262 16436 25316
rect 17218 25304 17224 25316
rect 17276 25304 17282 25356
rect 17862 25276 17868 25288
rect 16592 25248 17868 25276
rect 16592 25220 16620 25248
rect 17862 25236 17868 25248
rect 17920 25276 17926 25288
rect 18616 25285 18644 25384
rect 19904 25356 19932 25384
rect 19242 25344 19248 25356
rect 18708 25316 19248 25344
rect 18708 25285 18736 25316
rect 19242 25304 19248 25316
rect 19300 25304 19306 25356
rect 19352 25316 19840 25344
rect 18141 25279 18199 25285
rect 18141 25276 18153 25279
rect 17920 25248 18153 25276
rect 17920 25236 17926 25248
rect 18141 25245 18153 25248
rect 18187 25245 18199 25279
rect 18141 25239 18199 25245
rect 18601 25279 18659 25285
rect 18601 25245 18613 25279
rect 18647 25245 18659 25279
rect 18601 25239 18659 25245
rect 18693 25279 18751 25285
rect 18693 25245 18705 25279
rect 18739 25245 18751 25279
rect 18693 25239 18751 25245
rect 18874 25236 18880 25288
rect 18932 25285 18938 25288
rect 18932 25279 18961 25285
rect 18949 25245 18961 25279
rect 18932 25239 18961 25245
rect 18932 25236 18938 25239
rect 19058 25236 19064 25288
rect 19116 25236 19122 25288
rect 19352 25285 19380 25316
rect 19812 25288 19840 25316
rect 19886 25304 19892 25356
rect 19944 25304 19950 25356
rect 20625 25347 20683 25353
rect 20625 25344 20637 25347
rect 20364 25316 20637 25344
rect 19337 25279 19395 25285
rect 19337 25245 19349 25279
rect 19383 25245 19395 25279
rect 19337 25239 19395 25245
rect 19426 25236 19432 25288
rect 19484 25276 19490 25288
rect 19521 25279 19579 25285
rect 19521 25276 19533 25279
rect 19484 25248 19533 25276
rect 19484 25236 19490 25248
rect 19521 25245 19533 25248
rect 19567 25245 19579 25279
rect 19521 25239 19579 25245
rect 19794 25236 19800 25288
rect 19852 25236 19858 25288
rect 7282 25208 7288 25220
rect 6595 25180 7288 25208
rect 6595 25177 6607 25180
rect 6549 25171 6607 25177
rect 7282 25168 7288 25180
rect 7340 25168 7346 25220
rect 14918 25168 14924 25220
rect 14976 25208 14982 25220
rect 15289 25211 15347 25217
rect 15289 25208 15301 25211
rect 14976 25180 15301 25208
rect 14976 25168 14982 25180
rect 15289 25177 15301 25180
rect 15335 25177 15347 25211
rect 15289 25171 15347 25177
rect 16574 25168 16580 25220
rect 16632 25168 16638 25220
rect 16945 25211 17003 25217
rect 16945 25208 16957 25211
rect 16776 25180 16957 25208
rect 5132 25112 5396 25140
rect 5132 25100 5138 25112
rect 5718 25100 5724 25152
rect 5776 25140 5782 25152
rect 6749 25143 6807 25149
rect 6749 25140 6761 25143
rect 5776 25112 6761 25140
rect 5776 25100 5782 25112
rect 6749 25109 6761 25112
rect 6795 25140 6807 25143
rect 7466 25140 7472 25152
rect 6795 25112 7472 25140
rect 6795 25109 6807 25112
rect 6749 25103 6807 25109
rect 7466 25100 7472 25112
rect 7524 25100 7530 25152
rect 11882 25100 11888 25152
rect 11940 25100 11946 25152
rect 16776 25149 16804 25180
rect 16945 25177 16957 25180
rect 16991 25177 17003 25211
rect 16945 25171 17003 25177
rect 17402 25168 17408 25220
rect 17460 25208 17466 25220
rect 17460 25180 18552 25208
rect 17460 25168 17466 25180
rect 16761 25143 16819 25149
rect 16761 25109 16773 25143
rect 16807 25109 16819 25143
rect 16761 25103 16819 25109
rect 17034 25100 17040 25152
rect 17092 25100 17098 25152
rect 18414 25100 18420 25152
rect 18472 25100 18478 25152
rect 18524 25140 18552 25180
rect 18782 25168 18788 25220
rect 18840 25168 18846 25220
rect 19613 25211 19671 25217
rect 19613 25208 19625 25211
rect 19076 25180 19625 25208
rect 19076 25140 19104 25180
rect 19613 25177 19625 25180
rect 19659 25177 19671 25211
rect 19613 25171 19671 25177
rect 20070 25168 20076 25220
rect 20128 25208 20134 25220
rect 20364 25217 20392 25316
rect 20625 25313 20637 25316
rect 20671 25313 20683 25347
rect 20625 25307 20683 25313
rect 20901 25347 20959 25353
rect 20901 25313 20913 25347
rect 20947 25344 20959 25347
rect 21266 25344 21272 25356
rect 20947 25316 21272 25344
rect 20947 25313 20959 25316
rect 20901 25307 20959 25313
rect 21266 25304 21272 25316
rect 21324 25304 21330 25356
rect 20349 25211 20407 25217
rect 20349 25208 20361 25211
rect 20128 25180 20361 25208
rect 20128 25168 20134 25180
rect 20349 25177 20361 25180
rect 20395 25177 20407 25211
rect 20349 25171 20407 25177
rect 20806 25168 20812 25220
rect 20864 25208 20870 25220
rect 20864 25180 21390 25208
rect 20864 25168 20870 25180
rect 22646 25168 22652 25220
rect 22704 25168 22710 25220
rect 18524 25112 19104 25140
rect 19150 25100 19156 25152
rect 19208 25140 19214 25152
rect 19429 25143 19487 25149
rect 19429 25140 19441 25143
rect 19208 25112 19441 25140
rect 19208 25100 19214 25112
rect 19429 25109 19441 25112
rect 19475 25109 19487 25143
rect 19429 25103 19487 25109
rect 1104 25050 29595 25072
rect 1104 24998 8032 25050
rect 8084 24998 8096 25050
rect 8148 24998 8160 25050
rect 8212 24998 8224 25050
rect 8276 24998 8288 25050
rect 8340 24998 15115 25050
rect 15167 24998 15179 25050
rect 15231 24998 15243 25050
rect 15295 24998 15307 25050
rect 15359 24998 15371 25050
rect 15423 24998 22198 25050
rect 22250 24998 22262 25050
rect 22314 24998 22326 25050
rect 22378 24998 22390 25050
rect 22442 24998 22454 25050
rect 22506 24998 29281 25050
rect 29333 24998 29345 25050
rect 29397 24998 29409 25050
rect 29461 24998 29473 25050
rect 29525 24998 29537 25050
rect 29589 24998 29595 25050
rect 1104 24976 29595 24998
rect 3160 24908 5028 24936
rect 3160 24809 3188 24908
rect 5000 24880 5028 24908
rect 5258 24896 5264 24948
rect 5316 24896 5322 24948
rect 5353 24939 5411 24945
rect 5353 24905 5365 24939
rect 5399 24936 5411 24939
rect 5442 24936 5448 24948
rect 5399 24908 5448 24936
rect 5399 24905 5411 24908
rect 5353 24899 5411 24905
rect 5442 24896 5448 24908
rect 5500 24896 5506 24948
rect 6454 24896 6460 24948
rect 6512 24936 6518 24948
rect 7377 24939 7435 24945
rect 7377 24936 7389 24939
rect 6512 24908 7389 24936
rect 6512 24896 6518 24908
rect 7377 24905 7389 24908
rect 7423 24905 7435 24939
rect 7377 24899 7435 24905
rect 7466 24896 7472 24948
rect 7524 24896 7530 24948
rect 14918 24896 14924 24948
rect 14976 24896 14982 24948
rect 17126 24936 17132 24948
rect 15396 24908 17132 24936
rect 3510 24828 3516 24880
rect 3568 24868 3574 24880
rect 3568 24840 3910 24868
rect 3568 24828 3574 24840
rect 4890 24828 4896 24880
rect 4948 24828 4954 24880
rect 4982 24828 4988 24880
rect 5040 24828 5046 24880
rect 5276 24868 5304 24896
rect 5276 24840 6408 24868
rect 3145 24803 3203 24809
rect 3145 24769 3157 24803
rect 3191 24769 3203 24803
rect 4908 24800 4936 24828
rect 5169 24803 5227 24809
rect 5169 24800 5181 24803
rect 4908 24772 5181 24800
rect 3145 24763 3203 24769
rect 5169 24769 5181 24772
rect 5215 24769 5227 24803
rect 5626 24800 5632 24812
rect 5169 24763 5227 24769
rect 5460 24772 5632 24800
rect 3418 24692 3424 24744
rect 3476 24692 3482 24744
rect 4614 24692 4620 24744
rect 4672 24732 4678 24744
rect 4893 24735 4951 24741
rect 4893 24732 4905 24735
rect 4672 24704 4905 24732
rect 4672 24692 4678 24704
rect 4893 24701 4905 24704
rect 4939 24701 4951 24735
rect 4893 24695 4951 24701
rect 4985 24735 5043 24741
rect 4985 24701 4997 24735
rect 5031 24732 5043 24735
rect 5460 24732 5488 24772
rect 5626 24760 5632 24772
rect 5684 24760 5690 24812
rect 6380 24809 6408 24840
rect 6730 24828 6736 24880
rect 6788 24868 6794 24880
rect 7285 24871 7343 24877
rect 7285 24868 7297 24871
rect 6788 24840 7297 24868
rect 6788 24828 6794 24840
rect 7285 24837 7297 24840
rect 7331 24837 7343 24871
rect 7285 24831 7343 24837
rect 11793 24871 11851 24877
rect 11793 24837 11805 24871
rect 11839 24868 11851 24871
rect 11882 24868 11888 24880
rect 11839 24840 11888 24868
rect 11839 24837 11851 24840
rect 11793 24831 11851 24837
rect 11882 24828 11888 24840
rect 11940 24828 11946 24880
rect 14090 24868 14096 24880
rect 13018 24854 14096 24868
rect 13004 24840 14096 24854
rect 6365 24803 6423 24809
rect 6365 24769 6377 24803
rect 6411 24800 6423 24803
rect 6546 24800 6552 24812
rect 6411 24772 6552 24800
rect 6411 24769 6423 24772
rect 6365 24763 6423 24769
rect 6546 24760 6552 24772
rect 6604 24760 6610 24812
rect 7650 24760 7656 24812
rect 7708 24800 7714 24812
rect 7837 24803 7895 24809
rect 7837 24800 7849 24803
rect 7708 24772 7849 24800
rect 7708 24760 7714 24772
rect 7837 24769 7849 24772
rect 7883 24769 7895 24803
rect 7837 24763 7895 24769
rect 9214 24760 9220 24812
rect 9272 24800 9278 24812
rect 9582 24800 9588 24812
rect 9272 24772 9588 24800
rect 9272 24760 9278 24772
rect 9582 24760 9588 24772
rect 9640 24760 9646 24812
rect 9674 24760 9680 24812
rect 9732 24760 9738 24812
rect 11422 24760 11428 24812
rect 11480 24800 11486 24812
rect 11517 24803 11575 24809
rect 11517 24800 11529 24803
rect 11480 24772 11529 24800
rect 11480 24760 11486 24772
rect 11517 24769 11529 24772
rect 11563 24769 11575 24803
rect 11517 24763 11575 24769
rect 5031 24704 5488 24732
rect 5537 24735 5595 24741
rect 5031 24701 5043 24704
rect 4985 24695 5043 24701
rect 5537 24701 5549 24735
rect 5583 24732 5595 24735
rect 5718 24732 5724 24744
rect 5583 24704 5724 24732
rect 5583 24701 5595 24704
rect 5537 24695 5595 24701
rect 4908 24664 4936 24695
rect 5718 24692 5724 24704
rect 5776 24692 5782 24744
rect 6822 24692 6828 24744
rect 6880 24732 6886 24744
rect 7668 24732 7696 24760
rect 8113 24735 8171 24741
rect 8113 24732 8125 24735
rect 6880 24704 7696 24732
rect 7760 24704 8125 24732
rect 6880 24692 6886 24704
rect 5258 24664 5264 24676
rect 4908 24636 5264 24664
rect 5258 24624 5264 24636
rect 5316 24624 5322 24676
rect 5994 24664 6000 24676
rect 5368 24636 6000 24664
rect 3510 24556 3516 24608
rect 3568 24596 3574 24608
rect 5074 24596 5080 24608
rect 3568 24568 5080 24596
rect 3568 24556 3574 24568
rect 5074 24556 5080 24568
rect 5132 24596 5138 24608
rect 5368 24596 5396 24636
rect 5994 24624 6000 24636
rect 6052 24624 6058 24676
rect 6181 24667 6239 24673
rect 6181 24633 6193 24667
rect 6227 24664 6239 24667
rect 6914 24664 6920 24676
rect 6227 24636 6920 24664
rect 6227 24633 6239 24636
rect 6181 24627 6239 24633
rect 6914 24624 6920 24636
rect 6972 24624 6978 24676
rect 7101 24667 7159 24673
rect 7101 24633 7113 24667
rect 7147 24664 7159 24667
rect 7282 24664 7288 24676
rect 7147 24636 7288 24664
rect 7147 24633 7159 24636
rect 7101 24627 7159 24633
rect 7282 24624 7288 24636
rect 7340 24624 7346 24676
rect 7760 24664 7788 24704
rect 8113 24701 8125 24704
rect 8159 24701 8171 24735
rect 8113 24695 8171 24701
rect 11330 24692 11336 24744
rect 11388 24732 11394 24744
rect 13004 24732 13032 24840
rect 14090 24828 14096 24840
rect 14148 24828 14154 24880
rect 14185 24871 14243 24877
rect 14185 24837 14197 24871
rect 14231 24868 14243 24871
rect 14826 24868 14832 24880
rect 14231 24840 14832 24868
rect 14231 24837 14243 24840
rect 14185 24831 14243 24837
rect 14826 24828 14832 24840
rect 14884 24828 14890 24880
rect 15396 24868 15424 24908
rect 17126 24896 17132 24908
rect 17184 24896 17190 24948
rect 19058 24936 19064 24948
rect 17972 24908 19064 24936
rect 17034 24868 17040 24880
rect 14936 24840 15424 24868
rect 15672 24840 15976 24868
rect 14369 24803 14427 24809
rect 14369 24769 14381 24803
rect 14415 24800 14427 24803
rect 14936 24800 14964 24840
rect 15672 24812 15700 24840
rect 14415 24772 14964 24800
rect 15105 24803 15163 24809
rect 14415 24769 14427 24772
rect 14369 24763 14427 24769
rect 15105 24769 15117 24803
rect 15151 24769 15163 24803
rect 15105 24763 15163 24769
rect 15197 24803 15255 24809
rect 15197 24769 15209 24803
rect 15243 24769 15255 24803
rect 15197 24763 15255 24769
rect 11388 24704 13032 24732
rect 11388 24692 11394 24704
rect 13538 24692 13544 24744
rect 13596 24692 13602 24744
rect 14458 24692 14464 24744
rect 14516 24692 14522 24744
rect 14550 24692 14556 24744
rect 14608 24692 14614 24744
rect 7576 24636 7788 24664
rect 5132 24568 5396 24596
rect 7009 24599 7067 24605
rect 5132 24556 5138 24568
rect 7009 24565 7021 24599
rect 7055 24596 7067 24599
rect 7576 24596 7604 24636
rect 14734 24624 14740 24676
rect 14792 24664 14798 24676
rect 15120 24664 15148 24763
rect 15212 24732 15240 24763
rect 15286 24760 15292 24812
rect 15344 24760 15350 24812
rect 15470 24809 15476 24812
rect 15427 24803 15476 24809
rect 15427 24769 15439 24803
rect 15473 24769 15476 24803
rect 15427 24763 15476 24769
rect 15470 24760 15476 24763
rect 15528 24760 15534 24812
rect 15654 24760 15660 24812
rect 15712 24760 15718 24812
rect 15841 24803 15899 24809
rect 15841 24769 15853 24803
rect 15887 24769 15899 24803
rect 15841 24766 15899 24769
rect 15764 24763 15899 24766
rect 15764 24744 15884 24763
rect 15565 24735 15623 24741
rect 15212 24704 15332 24732
rect 15304 24664 15332 24704
rect 15565 24701 15577 24735
rect 15611 24732 15623 24735
rect 15746 24732 15752 24744
rect 15611 24704 15752 24732
rect 15611 24701 15623 24704
rect 15565 24695 15623 24701
rect 15746 24692 15752 24704
rect 15804 24738 15884 24744
rect 15804 24692 15810 24738
rect 15948 24732 15976 24840
rect 16040 24840 16252 24868
rect 16040 24812 16068 24840
rect 16022 24760 16028 24812
rect 16080 24760 16086 24812
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24769 16175 24803
rect 16224 24800 16252 24840
rect 16776 24840 17040 24868
rect 16301 24803 16359 24809
rect 16301 24800 16313 24803
rect 16224 24772 16313 24800
rect 16117 24763 16175 24769
rect 16301 24769 16313 24772
rect 16347 24800 16359 24803
rect 16776 24800 16804 24840
rect 17034 24828 17040 24840
rect 17092 24828 17098 24880
rect 16347 24772 16804 24800
rect 16853 24803 16911 24809
rect 16347 24769 16359 24772
rect 16301 24763 16359 24769
rect 16853 24769 16865 24803
rect 16899 24769 16911 24803
rect 16853 24763 16911 24769
rect 16132 24732 16160 24763
rect 16868 24732 16896 24763
rect 17034 24732 17040 24744
rect 15948 24704 17040 24732
rect 17034 24692 17040 24704
rect 17092 24692 17098 24744
rect 17144 24732 17172 24896
rect 17972 24868 18000 24908
rect 19058 24896 19064 24908
rect 19116 24896 19122 24948
rect 17880 24840 18000 24868
rect 18049 24871 18107 24877
rect 17880 24809 17908 24840
rect 18049 24837 18061 24871
rect 18095 24868 18107 24871
rect 18322 24868 18328 24880
rect 18095 24840 18328 24868
rect 18095 24837 18107 24840
rect 18049 24831 18107 24837
rect 18322 24828 18328 24840
rect 18380 24828 18386 24880
rect 18414 24828 18420 24880
rect 18472 24868 18478 24880
rect 18693 24871 18751 24877
rect 18693 24868 18705 24871
rect 18472 24840 18705 24868
rect 18472 24828 18478 24840
rect 18693 24837 18705 24840
rect 18739 24837 18751 24871
rect 18693 24831 18751 24837
rect 19334 24828 19340 24880
rect 19392 24828 19398 24880
rect 20254 24828 20260 24880
rect 20312 24868 20318 24880
rect 21085 24871 21143 24877
rect 21085 24868 21097 24871
rect 20312 24840 21097 24868
rect 20312 24828 20318 24840
rect 21085 24837 21097 24840
rect 21131 24837 21143 24871
rect 21085 24831 21143 24837
rect 17865 24803 17923 24809
rect 17865 24769 17877 24803
rect 17911 24769 17923 24803
rect 17865 24763 17923 24769
rect 17954 24760 17960 24812
rect 18012 24760 18018 24812
rect 18138 24760 18144 24812
rect 18196 24809 18202 24812
rect 18196 24803 18225 24809
rect 18213 24769 18225 24803
rect 20349 24803 20407 24809
rect 20349 24800 20361 24803
rect 18196 24763 18225 24769
rect 20180 24772 20361 24800
rect 18196 24760 18202 24763
rect 18325 24735 18383 24741
rect 18325 24732 18337 24735
rect 17144 24704 18337 24732
rect 18325 24701 18337 24704
rect 18371 24701 18383 24735
rect 18325 24695 18383 24701
rect 18417 24735 18475 24741
rect 18417 24701 18429 24735
rect 18463 24732 18475 24735
rect 20070 24732 20076 24744
rect 18463 24704 20076 24732
rect 18463 24701 18475 24704
rect 18417 24695 18475 24701
rect 16025 24667 16083 24673
rect 16025 24664 16037 24667
rect 14792 24636 15240 24664
rect 15304 24636 16037 24664
rect 14792 24624 14798 24636
rect 7055 24568 7604 24596
rect 7055 24565 7067 24568
rect 7009 24559 7067 24565
rect 7650 24556 7656 24608
rect 7708 24556 7714 24608
rect 9585 24599 9643 24605
rect 9585 24565 9597 24599
rect 9631 24596 9643 24599
rect 9769 24599 9827 24605
rect 9769 24596 9781 24599
rect 9631 24568 9781 24596
rect 9631 24565 9643 24568
rect 9585 24559 9643 24565
rect 9769 24565 9781 24568
rect 9815 24565 9827 24599
rect 9769 24559 9827 24565
rect 10137 24599 10195 24605
rect 10137 24565 10149 24599
rect 10183 24596 10195 24599
rect 10410 24596 10416 24608
rect 10183 24568 10416 24596
rect 10183 24565 10195 24568
rect 10137 24559 10195 24565
rect 10410 24556 10416 24568
rect 10468 24556 10474 24608
rect 15212 24596 15240 24636
rect 16025 24633 16037 24636
rect 16071 24633 16083 24667
rect 16025 24627 16083 24633
rect 16114 24624 16120 24676
rect 16172 24664 16178 24676
rect 17681 24667 17739 24673
rect 16172 24636 16988 24664
rect 16172 24624 16178 24636
rect 16960 24605 16988 24636
rect 17681 24633 17693 24667
rect 17727 24664 17739 24667
rect 18230 24664 18236 24676
rect 17727 24636 18236 24664
rect 17727 24633 17739 24636
rect 17681 24627 17739 24633
rect 18230 24624 18236 24636
rect 18288 24624 18294 24676
rect 16209 24599 16267 24605
rect 16209 24596 16221 24599
rect 15212 24568 16221 24596
rect 16209 24565 16221 24568
rect 16255 24565 16267 24599
rect 16209 24559 16267 24565
rect 16945 24599 17003 24605
rect 16945 24565 16957 24599
rect 16991 24565 17003 24599
rect 18340 24596 18368 24695
rect 20070 24692 20076 24704
rect 20128 24692 20134 24744
rect 20180 24741 20208 24772
rect 20349 24769 20361 24772
rect 20395 24769 20407 24803
rect 20349 24763 20407 24769
rect 20714 24760 20720 24812
rect 20772 24800 20778 24812
rect 20809 24803 20867 24809
rect 20809 24800 20821 24803
rect 20772 24772 20821 24800
rect 20772 24760 20778 24772
rect 20809 24769 20821 24772
rect 20855 24769 20867 24803
rect 20809 24763 20867 24769
rect 20165 24735 20223 24741
rect 20165 24701 20177 24735
rect 20211 24701 20223 24735
rect 20165 24695 20223 24701
rect 19426 24596 19432 24608
rect 18340 24568 19432 24596
rect 16945 24559 17003 24565
rect 19426 24556 19432 24568
rect 19484 24556 19490 24608
rect 20070 24556 20076 24608
rect 20128 24596 20134 24608
rect 20441 24599 20499 24605
rect 20441 24596 20453 24599
rect 20128 24568 20453 24596
rect 20128 24556 20134 24568
rect 20441 24565 20453 24568
rect 20487 24565 20499 24599
rect 20441 24559 20499 24565
rect 1104 24506 29440 24528
rect 1104 24454 4491 24506
rect 4543 24454 4555 24506
rect 4607 24454 4619 24506
rect 4671 24454 4683 24506
rect 4735 24454 4747 24506
rect 4799 24454 11574 24506
rect 11626 24454 11638 24506
rect 11690 24454 11702 24506
rect 11754 24454 11766 24506
rect 11818 24454 11830 24506
rect 11882 24454 18657 24506
rect 18709 24454 18721 24506
rect 18773 24454 18785 24506
rect 18837 24454 18849 24506
rect 18901 24454 18913 24506
rect 18965 24454 25740 24506
rect 25792 24454 25804 24506
rect 25856 24454 25868 24506
rect 25920 24454 25932 24506
rect 25984 24454 25996 24506
rect 26048 24454 29440 24506
rect 1104 24432 29440 24454
rect 3418 24352 3424 24404
rect 3476 24392 3482 24404
rect 4065 24395 4123 24401
rect 4065 24392 4077 24395
rect 3476 24364 4077 24392
rect 3476 24352 3482 24364
rect 4065 24361 4077 24364
rect 4111 24361 4123 24395
rect 4065 24355 4123 24361
rect 5350 24352 5356 24404
rect 5408 24352 5414 24404
rect 9674 24392 9680 24404
rect 6886 24364 9680 24392
rect 5368 24324 5396 24352
rect 4264 24296 5396 24324
rect 4264 24197 4292 24296
rect 6546 24284 6552 24336
rect 6604 24324 6610 24336
rect 6886 24324 6914 24364
rect 9674 24352 9680 24364
rect 9732 24352 9738 24404
rect 15286 24352 15292 24404
rect 15344 24392 15350 24404
rect 16022 24392 16028 24404
rect 15344 24364 16028 24392
rect 15344 24352 15350 24364
rect 16022 24352 16028 24364
rect 16080 24352 16086 24404
rect 19242 24352 19248 24404
rect 19300 24352 19306 24404
rect 19886 24352 19892 24404
rect 19944 24352 19950 24404
rect 6604 24296 6914 24324
rect 7009 24327 7067 24333
rect 6604 24284 6610 24296
rect 7009 24293 7021 24327
rect 7055 24324 7067 24327
rect 7466 24324 7472 24336
rect 7055 24296 7472 24324
rect 7055 24293 7067 24296
rect 7009 24287 7067 24293
rect 7466 24284 7472 24296
rect 7524 24284 7530 24336
rect 14458 24284 14464 24336
rect 14516 24324 14522 24336
rect 14516 24296 16160 24324
rect 14516 24284 14522 24296
rect 16132 24268 16160 24296
rect 19426 24284 19432 24336
rect 19484 24324 19490 24336
rect 19484 24296 20024 24324
rect 19484 24284 19490 24296
rect 4982 24216 4988 24268
rect 5040 24256 5046 24268
rect 5261 24259 5319 24265
rect 5261 24256 5273 24259
rect 5040 24228 5273 24256
rect 5040 24216 5046 24228
rect 5261 24225 5273 24228
rect 5307 24256 5319 24259
rect 6822 24256 6828 24268
rect 5307 24228 6828 24256
rect 5307 24225 5319 24228
rect 5261 24219 5319 24225
rect 6822 24216 6828 24228
rect 6880 24216 6886 24268
rect 11609 24259 11667 24265
rect 11609 24225 11621 24259
rect 11655 24256 11667 24259
rect 15010 24256 15016 24268
rect 11655 24228 15016 24256
rect 11655 24225 11667 24228
rect 11609 24219 11667 24225
rect 15010 24216 15016 24228
rect 15068 24256 15074 24268
rect 15289 24259 15347 24265
rect 15289 24256 15301 24259
rect 15068 24228 15301 24256
rect 15068 24216 15074 24228
rect 15289 24225 15301 24228
rect 15335 24225 15347 24259
rect 15930 24256 15936 24268
rect 15289 24219 15347 24225
rect 15856 24228 15936 24256
rect 4249 24191 4307 24197
rect 4249 24157 4261 24191
rect 4295 24157 4307 24191
rect 4249 24151 4307 24157
rect 7006 24148 7012 24200
rect 7064 24188 7070 24200
rect 7101 24191 7159 24197
rect 7101 24188 7113 24191
rect 7064 24160 7113 24188
rect 7064 24148 7070 24160
rect 7101 24157 7113 24160
rect 7147 24157 7159 24191
rect 7101 24151 7159 24157
rect 7190 24148 7196 24200
rect 7248 24188 7254 24200
rect 7285 24191 7343 24197
rect 7285 24188 7297 24191
rect 7248 24160 7297 24188
rect 7248 24148 7254 24160
rect 7285 24157 7297 24160
rect 7331 24157 7343 24191
rect 7285 24151 7343 24157
rect 10042 24148 10048 24200
rect 10100 24148 10106 24200
rect 13906 24188 13912 24200
rect 13556 24160 13912 24188
rect 5537 24123 5595 24129
rect 5537 24089 5549 24123
rect 5583 24120 5595 24123
rect 5583 24092 5948 24120
rect 5583 24089 5595 24092
rect 5537 24083 5595 24089
rect 5920 24052 5948 24092
rect 5994 24080 6000 24132
rect 6052 24080 6058 24132
rect 6886 24092 7236 24120
rect 6886 24052 6914 24092
rect 7208 24061 7236 24092
rect 9508 24092 11836 24120
rect 9508 24064 9536 24092
rect 5920 24024 6914 24052
rect 7193 24055 7251 24061
rect 7193 24021 7205 24055
rect 7239 24021 7251 24055
rect 7193 24015 7251 24021
rect 9490 24012 9496 24064
rect 9548 24012 9554 24064
rect 9674 24012 9680 24064
rect 9732 24052 9738 24064
rect 10597 24055 10655 24061
rect 10597 24052 10609 24055
rect 9732 24024 10609 24052
rect 9732 24012 9738 24024
rect 10597 24021 10609 24024
rect 10643 24021 10655 24055
rect 11808 24052 11836 24092
rect 11882 24080 11888 24132
rect 11940 24080 11946 24132
rect 13446 24120 13452 24132
rect 13110 24092 13452 24120
rect 13446 24080 13452 24092
rect 13504 24120 13510 24132
rect 13556 24120 13584 24160
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 15856 24197 15884 24228
rect 15930 24216 15936 24228
rect 15988 24216 15994 24268
rect 16114 24216 16120 24268
rect 16172 24216 16178 24268
rect 16390 24216 16396 24268
rect 16448 24216 16454 24268
rect 15841 24191 15899 24197
rect 15841 24157 15853 24191
rect 15887 24157 15899 24191
rect 15841 24151 15899 24157
rect 16298 24148 16304 24200
rect 16356 24148 16362 24200
rect 17954 24148 17960 24200
rect 18012 24188 18018 24200
rect 19058 24188 19064 24200
rect 18012 24160 19064 24188
rect 18012 24148 18018 24160
rect 19058 24148 19064 24160
rect 19116 24188 19122 24200
rect 19628 24197 19656 24296
rect 19429 24191 19487 24197
rect 19429 24188 19441 24191
rect 19116 24160 19441 24188
rect 19116 24148 19122 24160
rect 19429 24157 19441 24160
rect 19475 24157 19487 24191
rect 19429 24151 19487 24157
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 19705 24191 19763 24197
rect 19705 24157 19717 24191
rect 19751 24157 19763 24191
rect 19705 24151 19763 24157
rect 13504 24092 13584 24120
rect 13633 24123 13691 24129
rect 13504 24080 13510 24092
rect 13633 24089 13645 24123
rect 13679 24089 13691 24123
rect 13633 24083 13691 24089
rect 14553 24123 14611 24129
rect 14553 24089 14565 24123
rect 14599 24120 14611 24123
rect 15010 24120 15016 24132
rect 14599 24092 15016 24120
rect 14599 24089 14611 24092
rect 14553 24083 14611 24089
rect 13648 24052 13676 24083
rect 15010 24080 15016 24092
rect 15068 24080 15074 24132
rect 15930 24080 15936 24132
rect 15988 24080 15994 24132
rect 16022 24080 16028 24132
rect 16080 24080 16086 24132
rect 16206 24129 16212 24132
rect 16163 24123 16212 24129
rect 16163 24089 16175 24123
rect 16209 24089 16212 24123
rect 16163 24083 16212 24089
rect 16206 24080 16212 24083
rect 16264 24080 16270 24132
rect 16669 24123 16727 24129
rect 16669 24089 16681 24123
rect 16715 24089 16727 24123
rect 16669 24083 16727 24089
rect 14366 24052 14372 24064
rect 11808 24024 14372 24052
rect 10597 24015 10655 24021
rect 14366 24012 14372 24024
rect 14424 24012 14430 24064
rect 15657 24055 15715 24061
rect 15657 24021 15669 24055
rect 15703 24052 15715 24055
rect 16684 24052 16712 24083
rect 17218 24080 17224 24132
rect 17276 24080 17282 24132
rect 18046 24080 18052 24132
rect 18104 24120 18110 24132
rect 18417 24123 18475 24129
rect 18417 24120 18429 24123
rect 18104 24092 18429 24120
rect 18104 24080 18110 24092
rect 18417 24089 18429 24092
rect 18463 24089 18475 24123
rect 18417 24083 18475 24089
rect 15703 24024 16712 24052
rect 19444 24052 19472 24151
rect 19720 24120 19748 24151
rect 19797 24123 19855 24129
rect 19797 24120 19809 24123
rect 19720 24092 19809 24120
rect 19797 24089 19809 24092
rect 19843 24120 19855 24123
rect 19886 24120 19892 24132
rect 19843 24092 19892 24120
rect 19843 24089 19855 24092
rect 19797 24083 19855 24089
rect 19886 24080 19892 24092
rect 19944 24080 19950 24132
rect 19996 24129 20024 24296
rect 20070 24148 20076 24200
rect 20128 24148 20134 24200
rect 19981 24123 20039 24129
rect 19981 24089 19993 24123
rect 20027 24120 20039 24123
rect 20254 24120 20260 24132
rect 20027 24092 20260 24120
rect 20027 24089 20039 24092
rect 19981 24083 20039 24089
rect 20254 24080 20260 24092
rect 20312 24080 20318 24132
rect 20070 24052 20076 24064
rect 19444 24024 20076 24052
rect 15703 24021 15715 24024
rect 15657 24015 15715 24021
rect 20070 24012 20076 24024
rect 20128 24012 20134 24064
rect 1104 23962 29595 23984
rect 1104 23910 8032 23962
rect 8084 23910 8096 23962
rect 8148 23910 8160 23962
rect 8212 23910 8224 23962
rect 8276 23910 8288 23962
rect 8340 23910 15115 23962
rect 15167 23910 15179 23962
rect 15231 23910 15243 23962
rect 15295 23910 15307 23962
rect 15359 23910 15371 23962
rect 15423 23910 22198 23962
rect 22250 23910 22262 23962
rect 22314 23910 22326 23962
rect 22378 23910 22390 23962
rect 22442 23910 22454 23962
rect 22506 23910 29281 23962
rect 29333 23910 29345 23962
rect 29397 23910 29409 23962
rect 29461 23910 29473 23962
rect 29525 23910 29537 23962
rect 29589 23910 29595 23962
rect 1104 23888 29595 23910
rect 5166 23808 5172 23860
rect 5224 23848 5230 23860
rect 7650 23848 7656 23860
rect 5224 23820 7656 23848
rect 5224 23808 5230 23820
rect 7650 23808 7656 23820
rect 7708 23808 7714 23860
rect 11882 23808 11888 23860
rect 11940 23808 11946 23860
rect 12986 23808 12992 23860
rect 13044 23808 13050 23860
rect 14737 23851 14795 23857
rect 14737 23848 14749 23851
rect 13280 23820 14749 23848
rect 5718 23740 5724 23792
rect 5776 23780 5782 23792
rect 9490 23780 9496 23792
rect 5776 23752 9496 23780
rect 5776 23740 5782 23752
rect 9490 23740 9496 23752
rect 9548 23740 9554 23792
rect 10778 23780 10784 23792
rect 10718 23752 10784 23780
rect 10778 23740 10784 23752
rect 10836 23780 10842 23792
rect 11330 23780 11336 23792
rect 10836 23752 11336 23780
rect 10836 23740 10842 23752
rect 11330 23740 11336 23752
rect 11388 23740 11394 23792
rect 11900 23780 11928 23808
rect 13280 23780 13308 23820
rect 14737 23817 14749 23820
rect 14783 23817 14795 23851
rect 14737 23811 14795 23817
rect 14826 23808 14832 23860
rect 14884 23848 14890 23860
rect 14884 23820 15700 23848
rect 14884 23808 14890 23820
rect 15672 23792 15700 23820
rect 15930 23808 15936 23860
rect 15988 23848 15994 23860
rect 17589 23851 17647 23857
rect 17589 23848 17601 23851
rect 15988 23820 17601 23848
rect 15988 23808 15994 23820
rect 17589 23817 17601 23820
rect 17635 23817 17647 23851
rect 19886 23848 19892 23860
rect 17589 23811 17647 23817
rect 17926 23820 19892 23848
rect 11900 23752 13308 23780
rect 13357 23783 13415 23789
rect 13357 23749 13369 23783
rect 13403 23749 13415 23783
rect 13357 23743 13415 23749
rect 14936 23752 15608 23780
rect 1486 23672 1492 23724
rect 1544 23672 1550 23724
rect 12802 23712 12808 23724
rect 10888 23684 12808 23712
rect 9217 23647 9275 23653
rect 9217 23613 9229 23647
rect 9263 23644 9275 23647
rect 9493 23647 9551 23653
rect 9263 23616 9352 23644
rect 9263 23613 9275 23616
rect 9217 23607 9275 23613
rect 9324 23520 9352 23616
rect 9493 23613 9505 23647
rect 9539 23644 9551 23647
rect 10888 23644 10916 23684
rect 12802 23672 12808 23684
rect 12860 23672 12866 23724
rect 11517 23647 11575 23653
rect 11517 23644 11529 23647
rect 9539 23616 10916 23644
rect 10980 23616 11529 23644
rect 9539 23613 9551 23616
rect 9493 23607 9551 23613
rect 1578 23468 1584 23520
rect 1636 23468 1642 23520
rect 9306 23468 9312 23520
rect 9364 23468 9370 23520
rect 10778 23468 10784 23520
rect 10836 23508 10842 23520
rect 10980 23517 11008 23616
rect 11517 23613 11529 23616
rect 11563 23613 11575 23647
rect 13372 23644 13400 23743
rect 13449 23715 13507 23721
rect 13449 23681 13461 23715
rect 13495 23712 13507 23715
rect 14553 23715 14611 23721
rect 14553 23712 14565 23715
rect 13495 23684 14565 23712
rect 13495 23681 13507 23684
rect 13449 23675 13507 23681
rect 14553 23681 14565 23684
rect 14599 23681 14611 23715
rect 14553 23675 14611 23681
rect 14829 23715 14887 23721
rect 14829 23681 14841 23715
rect 14875 23712 14887 23715
rect 14936 23712 14964 23752
rect 15580 23724 15608 23752
rect 15654 23740 15660 23792
rect 15712 23740 15718 23792
rect 16022 23740 16028 23792
rect 16080 23740 16086 23792
rect 16298 23740 16304 23792
rect 16356 23780 16362 23792
rect 17221 23783 17279 23789
rect 17221 23780 17233 23783
rect 16356 23752 17233 23780
rect 16356 23740 16362 23752
rect 17221 23749 17233 23752
rect 17267 23780 17279 23783
rect 17494 23780 17500 23792
rect 17267 23752 17500 23780
rect 17267 23749 17279 23752
rect 17221 23743 17279 23749
rect 17494 23740 17500 23752
rect 17552 23740 17558 23792
rect 14875 23684 14964 23712
rect 15013 23715 15071 23721
rect 14875 23681 14887 23684
rect 14829 23675 14887 23681
rect 15013 23681 15025 23715
rect 15059 23712 15071 23715
rect 15289 23715 15347 23721
rect 15059 23684 15240 23712
rect 15059 23681 15071 23684
rect 15013 23675 15071 23681
rect 13372 23616 13492 23644
rect 11517 23607 11575 23613
rect 10965 23511 11023 23517
rect 10965 23508 10977 23511
rect 10836 23480 10977 23508
rect 10836 23468 10842 23480
rect 10965 23477 10977 23480
rect 11011 23477 11023 23511
rect 10965 23471 11023 23477
rect 12158 23468 12164 23520
rect 12216 23468 12222 23520
rect 13464 23508 13492 23616
rect 13538 23604 13544 23656
rect 13596 23604 13602 23656
rect 14093 23647 14151 23653
rect 14093 23613 14105 23647
rect 14139 23613 14151 23647
rect 14093 23607 14151 23613
rect 14108 23576 14136 23607
rect 14366 23604 14372 23656
rect 14424 23644 14430 23656
rect 14461 23647 14519 23653
rect 14461 23644 14473 23647
rect 14424 23616 14473 23644
rect 14424 23604 14430 23616
rect 14461 23613 14473 23616
rect 14507 23613 14519 23647
rect 14568 23644 14596 23675
rect 15212 23656 15240 23684
rect 15289 23681 15301 23715
rect 15335 23712 15347 23715
rect 15378 23712 15384 23724
rect 15335 23684 15384 23712
rect 15335 23681 15347 23684
rect 15289 23675 15347 23681
rect 15378 23672 15384 23684
rect 15436 23672 15442 23724
rect 15473 23715 15531 23721
rect 15473 23681 15485 23715
rect 15519 23681 15531 23715
rect 15473 23675 15531 23681
rect 15105 23647 15163 23653
rect 15105 23644 15117 23647
rect 14568 23616 15117 23644
rect 14461 23607 14519 23613
rect 15105 23613 15117 23616
rect 15151 23613 15163 23647
rect 15105 23607 15163 23613
rect 15194 23604 15200 23656
rect 15252 23604 15258 23656
rect 14108 23548 15240 23576
rect 15212 23520 15240 23548
rect 14829 23511 14887 23517
rect 14829 23508 14841 23511
rect 13464 23480 14841 23508
rect 14829 23477 14841 23480
rect 14875 23477 14887 23511
rect 14829 23471 14887 23477
rect 15194 23468 15200 23520
rect 15252 23468 15258 23520
rect 15396 23508 15424 23672
rect 15488 23644 15516 23675
rect 15562 23672 15568 23724
rect 15620 23672 15626 23724
rect 16040 23712 16068 23740
rect 15672 23684 16068 23712
rect 15672 23644 15700 23684
rect 16114 23672 16120 23724
rect 16172 23712 16178 23724
rect 16945 23715 17003 23721
rect 16945 23712 16957 23715
rect 16172 23684 16957 23712
rect 16172 23672 16178 23684
rect 15488 23616 15700 23644
rect 15470 23536 15476 23588
rect 15528 23576 15534 23588
rect 15746 23576 15752 23588
rect 15528 23548 15752 23576
rect 15528 23536 15534 23548
rect 15746 23536 15752 23548
rect 15804 23536 15810 23588
rect 15930 23536 15936 23588
rect 15988 23536 15994 23588
rect 16117 23511 16175 23517
rect 16117 23508 16129 23511
rect 15396 23480 16129 23508
rect 16117 23477 16129 23480
rect 16163 23508 16175 23511
rect 16206 23508 16212 23520
rect 16163 23480 16212 23508
rect 16163 23477 16175 23480
rect 16117 23471 16175 23477
rect 16206 23468 16212 23480
rect 16264 23468 16270 23520
rect 16868 23508 16896 23684
rect 16945 23681 16957 23684
rect 16991 23681 17003 23715
rect 16945 23675 17003 23681
rect 17034 23672 17040 23724
rect 17092 23672 17098 23724
rect 17126 23672 17132 23724
rect 17184 23672 17190 23724
rect 17313 23715 17371 23721
rect 17313 23681 17325 23715
rect 17359 23712 17371 23715
rect 17773 23715 17831 23721
rect 17773 23712 17785 23715
rect 17359 23684 17785 23712
rect 17359 23681 17371 23684
rect 17313 23675 17371 23681
rect 17773 23681 17785 23684
rect 17819 23712 17831 23715
rect 17926 23712 17954 23820
rect 19886 23808 19892 23820
rect 19944 23848 19950 23860
rect 22646 23848 22652 23860
rect 19944 23820 22652 23848
rect 19944 23808 19950 23820
rect 22646 23808 22652 23820
rect 22704 23808 22710 23860
rect 17819 23684 17954 23712
rect 17819 23681 17831 23684
rect 17773 23675 17831 23681
rect 17052 23644 17080 23672
rect 17497 23647 17555 23653
rect 17497 23644 17509 23647
rect 17052 23616 17509 23644
rect 17497 23613 17509 23616
rect 17543 23613 17555 23647
rect 17497 23607 17555 23613
rect 17865 23647 17923 23653
rect 17865 23613 17877 23647
rect 17911 23613 17923 23647
rect 17865 23607 17923 23613
rect 17126 23536 17132 23588
rect 17184 23576 17190 23588
rect 17880 23576 17908 23607
rect 17954 23604 17960 23656
rect 18012 23604 18018 23656
rect 18046 23604 18052 23656
rect 18104 23604 18110 23656
rect 17184 23548 17908 23576
rect 17184 23536 17190 23548
rect 17972 23508 18000 23604
rect 16868 23480 18000 23508
rect 1104 23418 29440 23440
rect 1104 23366 4491 23418
rect 4543 23366 4555 23418
rect 4607 23366 4619 23418
rect 4671 23366 4683 23418
rect 4735 23366 4747 23418
rect 4799 23366 11574 23418
rect 11626 23366 11638 23418
rect 11690 23366 11702 23418
rect 11754 23366 11766 23418
rect 11818 23366 11830 23418
rect 11882 23366 18657 23418
rect 18709 23366 18721 23418
rect 18773 23366 18785 23418
rect 18837 23366 18849 23418
rect 18901 23366 18913 23418
rect 18965 23366 25740 23418
rect 25792 23366 25804 23418
rect 25856 23366 25868 23418
rect 25920 23366 25932 23418
rect 25984 23366 25996 23418
rect 26048 23366 29440 23418
rect 1104 23344 29440 23366
rect 10042 23264 10048 23316
rect 10100 23304 10106 23316
rect 10502 23304 10508 23316
rect 10100 23276 10508 23304
rect 10100 23264 10106 23276
rect 10502 23264 10508 23276
rect 10560 23304 10566 23316
rect 10781 23307 10839 23313
rect 10781 23304 10793 23307
rect 10560 23276 10793 23304
rect 10560 23264 10566 23276
rect 10781 23273 10793 23276
rect 10827 23273 10839 23307
rect 10781 23267 10839 23273
rect 14550 23264 14556 23316
rect 14608 23304 14614 23316
rect 14645 23307 14703 23313
rect 14645 23304 14657 23307
rect 14608 23276 14657 23304
rect 14608 23264 14614 23276
rect 14645 23273 14657 23276
rect 14691 23273 14703 23307
rect 14645 23267 14703 23273
rect 14918 23264 14924 23316
rect 14976 23264 14982 23316
rect 15010 23264 15016 23316
rect 15068 23304 15074 23316
rect 16390 23304 16396 23316
rect 15068 23276 16396 23304
rect 15068 23264 15074 23276
rect 16390 23264 16396 23276
rect 16448 23304 16454 23316
rect 17402 23304 17408 23316
rect 16448 23276 17408 23304
rect 16448 23264 16454 23276
rect 17402 23264 17408 23276
rect 17460 23264 17466 23316
rect 25222 23264 25228 23316
rect 25280 23264 25286 23316
rect 15028 23236 15056 23264
rect 12406 23208 15056 23236
rect 6822 23128 6828 23180
rect 6880 23128 6886 23180
rect 9033 23171 9091 23177
rect 9033 23137 9045 23171
rect 9079 23168 9091 23171
rect 9306 23168 9312 23180
rect 9079 23140 9312 23168
rect 9079 23137 9091 23140
rect 9033 23131 9091 23137
rect 9306 23128 9312 23140
rect 9364 23168 9370 23180
rect 11422 23168 11428 23180
rect 9364 23140 11428 23168
rect 9364 23128 9370 23140
rect 11422 23128 11428 23140
rect 11480 23168 11486 23180
rect 11609 23171 11667 23177
rect 11609 23168 11621 23171
rect 11480 23140 11621 23168
rect 11480 23128 11486 23140
rect 11609 23137 11621 23140
rect 11655 23137 11667 23171
rect 11609 23131 11667 23137
rect 4525 23103 4583 23109
rect 4525 23069 4537 23103
rect 4571 23100 4583 23103
rect 6178 23100 6184 23112
rect 4571 23072 6184 23100
rect 4571 23069 4583 23072
rect 4525 23063 4583 23069
rect 6178 23060 6184 23072
rect 6236 23060 6242 23112
rect 10686 23100 10692 23112
rect 10442 23072 10692 23100
rect 10686 23060 10692 23072
rect 10744 23060 10750 23112
rect 10870 23060 10876 23112
rect 10928 23100 10934 23112
rect 12406 23100 12434 23208
rect 15194 23196 15200 23248
rect 15252 23196 15258 23248
rect 15562 23196 15568 23248
rect 15620 23196 15626 23248
rect 15930 23196 15936 23248
rect 15988 23236 15994 23248
rect 17589 23239 17647 23245
rect 17589 23236 17601 23239
rect 15988 23208 17601 23236
rect 15988 23196 15994 23208
rect 17589 23205 17601 23208
rect 17635 23236 17647 23239
rect 18138 23236 18144 23248
rect 17635 23208 18144 23236
rect 17635 23205 17647 23208
rect 17589 23199 17647 23205
rect 18138 23196 18144 23208
rect 18196 23196 18202 23248
rect 14550 23128 14556 23180
rect 14608 23168 14614 23180
rect 14829 23171 14887 23177
rect 14829 23168 14841 23171
rect 14608 23140 14841 23168
rect 14608 23128 14614 23140
rect 14829 23137 14841 23140
rect 14875 23168 14887 23171
rect 14875 23140 15884 23168
rect 14875 23137 14887 23140
rect 14829 23131 14887 23137
rect 10928 23072 12434 23100
rect 10928 23060 10934 23072
rect 13538 23060 13544 23112
rect 13596 23100 13602 23112
rect 13998 23100 14004 23112
rect 13596 23072 14004 23100
rect 13596 23060 13602 23072
rect 13998 23060 14004 23072
rect 14056 23100 14062 23112
rect 14369 23103 14427 23109
rect 14369 23100 14381 23103
rect 14056 23072 14381 23100
rect 14056 23060 14062 23072
rect 14369 23069 14381 23072
rect 14415 23069 14427 23103
rect 14369 23063 14427 23069
rect 14734 23060 14740 23112
rect 14792 23060 14798 23112
rect 15013 23103 15071 23109
rect 15013 23069 15025 23103
rect 15059 23069 15071 23103
rect 15013 23063 15071 23069
rect 15289 23103 15347 23109
rect 15289 23069 15301 23103
rect 15335 23100 15347 23103
rect 15378 23100 15384 23112
rect 15335 23072 15384 23100
rect 15335 23069 15347 23072
rect 15289 23063 15347 23069
rect 5997 23035 6055 23041
rect 5997 23032 6009 23035
rect 5276 23004 6009 23032
rect 5276 22976 5304 23004
rect 5997 23001 6009 23004
rect 6043 23001 6055 23035
rect 5997 22995 6055 23001
rect 5074 22924 5080 22976
rect 5132 22924 5138 22976
rect 5258 22924 5264 22976
rect 5316 22924 5322 22976
rect 6012 22964 6040 22995
rect 9214 22992 9220 23044
rect 9272 23032 9278 23044
rect 9309 23035 9367 23041
rect 9309 23032 9321 23035
rect 9272 23004 9321 23032
rect 9272 22992 9278 23004
rect 9309 23001 9321 23004
rect 9355 23001 9367 23035
rect 10888 23032 10916 23060
rect 9309 22995 9367 23001
rect 10704 23004 10916 23032
rect 10704 22964 10732 23004
rect 13906 22992 13912 23044
rect 13964 23032 13970 23044
rect 14093 23035 14151 23041
rect 14093 23032 14105 23035
rect 13964 23004 14105 23032
rect 13964 22992 13970 23004
rect 14093 23001 14105 23004
rect 14139 23001 14151 23035
rect 15028 23032 15056 23063
rect 15378 23060 15384 23072
rect 15436 23060 15442 23112
rect 15856 23109 15884 23140
rect 16022 23128 16028 23180
rect 16080 23168 16086 23180
rect 20993 23171 21051 23177
rect 16080 23140 18368 23168
rect 16080 23128 16086 23140
rect 17604 23109 17632 23140
rect 18340 23112 18368 23140
rect 20993 23137 21005 23171
rect 21039 23168 21051 23171
rect 21634 23168 21640 23180
rect 21039 23140 21640 23168
rect 21039 23137 21051 23140
rect 20993 23131 21051 23137
rect 21634 23128 21640 23140
rect 21692 23128 21698 23180
rect 24302 23128 24308 23180
rect 24360 23168 24366 23180
rect 25038 23168 25044 23180
rect 24360 23140 25044 23168
rect 24360 23128 24366 23140
rect 25038 23128 25044 23140
rect 25096 23128 25102 23180
rect 15657 23103 15715 23109
rect 15563 23081 15621 23087
rect 15563 23047 15575 23081
rect 15609 23047 15621 23081
rect 15657 23069 15669 23103
rect 15703 23069 15715 23103
rect 15657 23063 15715 23069
rect 15841 23103 15899 23109
rect 15841 23069 15853 23103
rect 15887 23069 15899 23103
rect 15841 23063 15899 23069
rect 17589 23103 17647 23109
rect 17589 23069 17601 23103
rect 17635 23069 17647 23103
rect 17589 23063 17647 23069
rect 17773 23103 17831 23109
rect 17773 23069 17785 23103
rect 17819 23069 17831 23103
rect 17773 23063 17831 23069
rect 15563 23044 15621 23047
rect 15470 23032 15476 23044
rect 14093 22995 14151 23001
rect 14476 23004 15476 23032
rect 6012 22936 10732 22964
rect 14274 22924 14280 22976
rect 14332 22924 14338 22976
rect 14366 22924 14372 22976
rect 14424 22964 14430 22976
rect 14476 22973 14504 23004
rect 15470 22992 15476 23004
rect 15528 22992 15534 23044
rect 15562 22992 15568 23044
rect 15620 22992 15626 23044
rect 14461 22967 14519 22973
rect 14461 22964 14473 22967
rect 14424 22936 14473 22964
rect 14424 22924 14430 22936
rect 14461 22933 14473 22936
rect 14507 22933 14519 22967
rect 14461 22927 14519 22933
rect 14918 22924 14924 22976
rect 14976 22964 14982 22976
rect 15102 22964 15108 22976
rect 14976 22936 15108 22964
rect 14976 22924 14982 22936
rect 15102 22924 15108 22936
rect 15160 22964 15166 22976
rect 15672 22964 15700 23063
rect 16758 22992 16764 23044
rect 16816 23032 16822 23044
rect 17788 23032 17816 23063
rect 18322 23060 18328 23112
rect 18380 23060 18386 23112
rect 20714 23060 20720 23112
rect 20772 23060 20778 23112
rect 20806 23060 20812 23112
rect 20864 23060 20870 23112
rect 21085 23103 21143 23109
rect 21085 23069 21097 23103
rect 21131 23100 21143 23103
rect 21726 23100 21732 23112
rect 21131 23072 21732 23100
rect 21131 23069 21143 23072
rect 21085 23063 21143 23069
rect 21726 23060 21732 23072
rect 21784 23060 21790 23112
rect 24486 23060 24492 23112
rect 24544 23060 24550 23112
rect 24581 23103 24639 23109
rect 24581 23069 24593 23103
rect 24627 23069 24639 23103
rect 24581 23063 24639 23069
rect 24765 23103 24823 23109
rect 24765 23069 24777 23103
rect 24811 23100 24823 23103
rect 24857 23103 24915 23109
rect 24857 23100 24869 23103
rect 24811 23072 24869 23100
rect 24811 23069 24823 23072
rect 24765 23063 24823 23069
rect 24857 23069 24869 23072
rect 24903 23100 24915 23103
rect 24903 23072 25544 23100
rect 24903 23069 24915 23072
rect 24857 23063 24915 23069
rect 16816 23004 17816 23032
rect 16816 22992 16822 23004
rect 21174 22992 21180 23044
rect 21232 22992 21238 23044
rect 22554 22992 22560 23044
rect 22612 23032 22618 23044
rect 24596 23032 24624 23063
rect 25516 23044 25544 23072
rect 24670 23032 24676 23044
rect 22612 23004 24676 23032
rect 22612 22992 22618 23004
rect 24670 22992 24676 23004
rect 24728 22992 24734 23044
rect 25041 23035 25099 23041
rect 25041 23001 25053 23035
rect 25087 23001 25099 23035
rect 25041 22995 25099 23001
rect 16206 22964 16212 22976
rect 15160 22936 16212 22964
rect 15160 22924 15166 22936
rect 16206 22924 16212 22936
rect 16264 22924 16270 22976
rect 17586 22924 17592 22976
rect 17644 22964 17650 22976
rect 18046 22964 18052 22976
rect 17644 22936 18052 22964
rect 17644 22924 17650 22936
rect 18046 22924 18052 22936
rect 18104 22924 18110 22976
rect 20990 22924 20996 22976
rect 21048 22924 21054 22976
rect 23474 22924 23480 22976
rect 23532 22964 23538 22976
rect 24118 22964 24124 22976
rect 23532 22936 24124 22964
rect 23532 22924 23538 22936
rect 24118 22924 24124 22936
rect 24176 22964 24182 22976
rect 24762 22964 24768 22976
rect 24176 22936 24768 22964
rect 24176 22924 24182 22936
rect 24762 22924 24768 22936
rect 24820 22924 24826 22976
rect 24946 22924 24952 22976
rect 25004 22964 25010 22976
rect 25056 22964 25084 22995
rect 25498 22992 25504 23044
rect 25556 22992 25562 23044
rect 25004 22936 25084 22964
rect 25004 22924 25010 22936
rect 1104 22874 29595 22896
rect 1104 22822 8032 22874
rect 8084 22822 8096 22874
rect 8148 22822 8160 22874
rect 8212 22822 8224 22874
rect 8276 22822 8288 22874
rect 8340 22822 15115 22874
rect 15167 22822 15179 22874
rect 15231 22822 15243 22874
rect 15295 22822 15307 22874
rect 15359 22822 15371 22874
rect 15423 22822 22198 22874
rect 22250 22822 22262 22874
rect 22314 22822 22326 22874
rect 22378 22822 22390 22874
rect 22442 22822 22454 22874
rect 22506 22822 29281 22874
rect 29333 22822 29345 22874
rect 29397 22822 29409 22874
rect 29461 22822 29473 22874
rect 29525 22822 29537 22874
rect 29589 22822 29595 22874
rect 1104 22800 29595 22822
rect 6914 22720 6920 22772
rect 6972 22760 6978 22772
rect 10226 22760 10232 22772
rect 6972 22732 10232 22760
rect 6972 22720 6978 22732
rect 10226 22720 10232 22732
rect 10284 22760 10290 22772
rect 10284 22732 12480 22760
rect 10284 22720 10290 22732
rect 5258 22652 5264 22704
rect 5316 22652 5322 22704
rect 8205 22695 8263 22701
rect 8205 22692 8217 22695
rect 6748 22664 8217 22692
rect 6748 22633 6776 22664
rect 8205 22661 8217 22664
rect 8251 22661 8263 22695
rect 8205 22655 8263 22661
rect 8941 22695 8999 22701
rect 8941 22661 8953 22695
rect 8987 22692 8999 22695
rect 9674 22692 9680 22704
rect 8987 22664 9680 22692
rect 8987 22661 8999 22664
rect 8941 22655 8999 22661
rect 9674 22652 9680 22664
rect 9732 22652 9738 22704
rect 12452 22701 12480 22732
rect 12802 22720 12808 22772
rect 12860 22720 12866 22772
rect 15010 22720 15016 22772
rect 15068 22760 15074 22772
rect 15068 22732 15424 22760
rect 15068 22720 15074 22732
rect 12437 22695 12495 22701
rect 12437 22661 12449 22695
rect 12483 22661 12495 22695
rect 12437 22655 12495 22661
rect 12526 22652 12532 22704
rect 12584 22652 12590 22704
rect 15396 22701 15424 22732
rect 20714 22720 20720 22772
rect 20772 22760 20778 22772
rect 20901 22763 20959 22769
rect 20901 22760 20913 22763
rect 20772 22732 20913 22760
rect 20772 22720 20778 22732
rect 20901 22729 20913 22732
rect 20947 22729 20959 22763
rect 23474 22760 23480 22772
rect 20901 22723 20959 22729
rect 21468 22732 23480 22760
rect 15381 22695 15439 22701
rect 15381 22661 15393 22695
rect 15427 22661 15439 22695
rect 15381 22655 15439 22661
rect 6733 22627 6791 22633
rect 6733 22593 6745 22627
rect 6779 22593 6791 22627
rect 6733 22587 6791 22593
rect 6917 22627 6975 22633
rect 6917 22593 6929 22627
rect 6963 22593 6975 22627
rect 6917 22587 6975 22593
rect 7009 22627 7067 22633
rect 7009 22593 7021 22627
rect 7055 22593 7067 22627
rect 7009 22587 7067 22593
rect 7101 22627 7159 22633
rect 7101 22593 7113 22627
rect 7147 22624 7159 22627
rect 8110 22624 8116 22636
rect 7147 22596 8116 22624
rect 7147 22593 7159 22596
rect 7101 22587 7159 22593
rect 4525 22559 4583 22565
rect 4525 22525 4537 22559
rect 4571 22556 4583 22559
rect 5626 22556 5632 22568
rect 4571 22528 5632 22556
rect 4571 22525 4583 22528
rect 4525 22519 4583 22525
rect 5626 22516 5632 22528
rect 5684 22516 5690 22568
rect 5994 22516 6000 22568
rect 6052 22516 6058 22568
rect 6932 22556 6960 22587
rect 6840 22528 6960 22556
rect 4154 22380 4160 22432
rect 4212 22420 4218 22432
rect 5077 22423 5135 22429
rect 5077 22420 5089 22423
rect 4212 22392 5089 22420
rect 4212 22380 4218 22392
rect 5077 22389 5089 22392
rect 5123 22389 5135 22423
rect 6840 22420 6868 22528
rect 7024 22488 7052 22587
rect 8110 22584 8116 22596
rect 8168 22584 8174 22636
rect 8662 22584 8668 22636
rect 8720 22584 8726 22636
rect 8846 22584 8852 22636
rect 8904 22584 8910 22636
rect 9033 22627 9091 22633
rect 9033 22593 9045 22627
rect 9079 22593 9091 22627
rect 9033 22587 9091 22593
rect 7650 22516 7656 22568
rect 7708 22516 7714 22568
rect 9048 22556 9076 22587
rect 9306 22584 9312 22636
rect 9364 22584 9370 22636
rect 10962 22624 10968 22636
rect 10718 22596 10968 22624
rect 10962 22584 10968 22596
rect 11020 22584 11026 22636
rect 12158 22584 12164 22636
rect 12216 22624 12222 22636
rect 12253 22627 12311 22633
rect 12253 22624 12265 22627
rect 12216 22596 12265 22624
rect 12216 22584 12222 22596
rect 12253 22593 12265 22596
rect 12299 22593 12311 22627
rect 12253 22587 12311 22593
rect 12618 22584 12624 22636
rect 12676 22584 12682 22636
rect 15013 22627 15071 22633
rect 15013 22593 15025 22627
rect 15059 22593 15071 22627
rect 15013 22587 15071 22593
rect 15289 22627 15347 22633
rect 15289 22593 15301 22627
rect 15335 22624 15347 22627
rect 17313 22627 17371 22633
rect 17313 22624 17325 22627
rect 15335 22596 17325 22624
rect 15335 22593 15347 22596
rect 15289 22587 15347 22593
rect 17313 22593 17325 22596
rect 17359 22593 17371 22627
rect 17313 22587 17371 22593
rect 9585 22559 9643 22565
rect 9048 22528 9444 22556
rect 7024 22460 7788 22488
rect 7760 22432 7788 22460
rect 9214 22448 9220 22500
rect 9272 22448 9278 22500
rect 9416 22432 9444 22528
rect 9585 22525 9597 22559
rect 9631 22556 9643 22559
rect 9950 22556 9956 22568
rect 9631 22528 9956 22556
rect 9631 22525 9643 22528
rect 9585 22519 9643 22525
rect 9950 22516 9956 22528
rect 10008 22516 10014 22568
rect 11057 22559 11115 22565
rect 11057 22525 11069 22559
rect 11103 22556 11115 22559
rect 11422 22556 11428 22568
rect 11103 22528 11428 22556
rect 11103 22525 11115 22528
rect 11057 22519 11115 22525
rect 11422 22516 11428 22528
rect 11480 22556 11486 22568
rect 11517 22559 11575 22565
rect 11517 22556 11529 22559
rect 11480 22528 11529 22556
rect 11480 22516 11486 22528
rect 11517 22525 11529 22528
rect 11563 22525 11575 22559
rect 11517 22519 11575 22525
rect 13906 22448 13912 22500
rect 13964 22488 13970 22500
rect 15028 22488 15056 22587
rect 20714 22584 20720 22636
rect 20772 22584 20778 22636
rect 20806 22584 20812 22636
rect 20864 22584 20870 22636
rect 20916 22624 20944 22723
rect 21468 22633 21496 22732
rect 23474 22720 23480 22732
rect 23532 22720 23538 22772
rect 24397 22763 24455 22769
rect 23768 22732 24348 22760
rect 21726 22692 21732 22704
rect 21560 22664 21732 22692
rect 21560 22633 21588 22664
rect 21726 22652 21732 22664
rect 21784 22652 21790 22704
rect 22830 22692 22836 22704
rect 22756 22664 22836 22692
rect 21269 22627 21327 22633
rect 21269 22624 21281 22627
rect 20916 22596 21281 22624
rect 21269 22593 21281 22596
rect 21315 22593 21327 22627
rect 21269 22587 21327 22593
rect 21453 22627 21511 22633
rect 21453 22593 21465 22627
rect 21499 22593 21511 22627
rect 21453 22587 21511 22593
rect 21545 22627 21603 22633
rect 21545 22593 21557 22627
rect 21591 22593 21603 22627
rect 21545 22587 21603 22593
rect 21634 22584 21640 22636
rect 21692 22624 21698 22636
rect 22756 22633 22784 22664
rect 22830 22652 22836 22664
rect 22888 22692 22894 22704
rect 23201 22695 23259 22701
rect 23201 22692 23213 22695
rect 22888 22664 23213 22692
rect 22888 22652 22894 22664
rect 23201 22661 23213 22664
rect 23247 22661 23259 22695
rect 23768 22692 23796 22732
rect 24213 22695 24271 22701
rect 24213 22692 24225 22695
rect 23201 22655 23259 22661
rect 23584 22664 23796 22692
rect 23584 22636 23612 22664
rect 21821 22627 21879 22633
rect 21821 22624 21833 22627
rect 21692 22596 21833 22624
rect 21692 22584 21698 22596
rect 21821 22593 21833 22596
rect 21867 22593 21879 22627
rect 21999 22627 22057 22633
rect 21999 22624 22011 22627
rect 21821 22587 21879 22593
rect 21928 22596 22011 22624
rect 15197 22559 15255 22565
rect 15197 22525 15209 22559
rect 15243 22556 15255 22559
rect 15654 22556 15660 22568
rect 15243 22528 15660 22556
rect 15243 22525 15255 22528
rect 15197 22519 15255 22525
rect 15654 22516 15660 22528
rect 15712 22516 15718 22568
rect 16209 22559 16267 22565
rect 16209 22525 16221 22559
rect 16255 22556 16267 22559
rect 16482 22556 16488 22568
rect 16255 22528 16488 22556
rect 16255 22525 16267 22528
rect 16209 22519 16267 22525
rect 16482 22516 16488 22528
rect 16540 22516 16546 22568
rect 16666 22516 16672 22568
rect 16724 22516 16730 22568
rect 20438 22516 20444 22568
rect 20496 22556 20502 22568
rect 20533 22559 20591 22565
rect 20533 22556 20545 22559
rect 20496 22528 20545 22556
rect 20496 22516 20502 22528
rect 20533 22525 20545 22528
rect 20579 22525 20591 22559
rect 20824 22556 20852 22584
rect 21358 22556 21364 22568
rect 20824 22528 21364 22556
rect 20533 22519 20591 22525
rect 21358 22516 21364 22528
rect 21416 22516 21422 22568
rect 21928 22556 21956 22596
rect 21999 22593 22011 22596
rect 22045 22593 22057 22627
rect 21999 22587 22057 22593
rect 22741 22627 22799 22633
rect 22741 22593 22753 22627
rect 22787 22593 22799 22627
rect 22741 22587 22799 22593
rect 22925 22627 22983 22633
rect 22925 22593 22937 22627
rect 22971 22593 22983 22627
rect 22925 22587 22983 22593
rect 22940 22556 22968 22587
rect 23014 22584 23020 22636
rect 23072 22624 23078 22636
rect 23109 22627 23167 22633
rect 23109 22624 23121 22627
rect 23072 22596 23121 22624
rect 23072 22584 23078 22596
rect 23109 22593 23121 22596
rect 23155 22593 23167 22627
rect 23109 22587 23167 22593
rect 23290 22584 23296 22636
rect 23348 22584 23354 22636
rect 23566 22584 23572 22636
rect 23624 22584 23630 22636
rect 23768 22633 23796 22664
rect 23952 22664 24225 22692
rect 23952 22633 23980 22664
rect 24213 22661 24225 22664
rect 24259 22661 24271 22695
rect 24213 22655 24271 22661
rect 24320 22636 24348 22732
rect 24397 22729 24409 22763
rect 24443 22760 24455 22763
rect 25314 22760 25320 22772
rect 24443 22732 25320 22760
rect 24443 22729 24455 22732
rect 24397 22723 24455 22729
rect 25314 22720 25320 22732
rect 25372 22720 25378 22772
rect 24946 22692 24952 22704
rect 24412 22664 24952 22692
rect 24412 22636 24440 22664
rect 23661 22627 23719 22633
rect 23661 22593 23673 22627
rect 23707 22593 23719 22627
rect 23661 22587 23719 22593
rect 23753 22627 23811 22633
rect 23753 22593 23765 22627
rect 23799 22593 23811 22627
rect 23753 22587 23811 22593
rect 23937 22627 23995 22633
rect 23937 22593 23949 22627
rect 23983 22593 23995 22627
rect 23937 22587 23995 22593
rect 24029 22627 24087 22633
rect 24029 22593 24041 22627
rect 24075 22593 24087 22627
rect 24029 22587 24087 22593
rect 23382 22556 23388 22568
rect 21560 22528 23388 22556
rect 15930 22488 15936 22500
rect 13964 22460 14964 22488
rect 15028 22460 15936 22488
rect 13964 22448 13970 22460
rect 6914 22420 6920 22432
rect 6840 22392 6920 22420
rect 5077 22383 5135 22389
rect 6914 22380 6920 22392
rect 6972 22380 6978 22432
rect 7282 22380 7288 22432
rect 7340 22380 7346 22432
rect 7742 22380 7748 22432
rect 7800 22380 7806 22432
rect 9398 22380 9404 22432
rect 9456 22380 9462 22432
rect 10226 22380 10232 22432
rect 10284 22420 10290 22432
rect 12161 22423 12219 22429
rect 12161 22420 12173 22423
rect 10284 22392 12173 22420
rect 10284 22380 10290 22392
rect 12161 22389 12173 22392
rect 12207 22389 12219 22423
rect 12161 22383 12219 22389
rect 14826 22380 14832 22432
rect 14884 22380 14890 22432
rect 14936 22420 14964 22460
rect 15930 22448 15936 22460
rect 15988 22448 15994 22500
rect 21174 22448 21180 22500
rect 21232 22488 21238 22500
rect 21450 22488 21456 22500
rect 21232 22460 21456 22488
rect 21232 22448 21238 22460
rect 21450 22448 21456 22460
rect 21508 22448 21514 22500
rect 21560 22432 21588 22528
rect 23382 22516 23388 22528
rect 23440 22516 23446 22568
rect 21634 22448 21640 22500
rect 21692 22488 21698 22500
rect 23676 22488 23704 22587
rect 24044 22500 24072 22587
rect 24118 22584 24124 22636
rect 24176 22584 24182 22636
rect 24302 22584 24308 22636
rect 24360 22584 24366 22636
rect 24394 22584 24400 22636
rect 24452 22584 24458 22636
rect 24578 22584 24584 22636
rect 24636 22584 24642 22636
rect 24780 22633 24808 22664
rect 24946 22652 24952 22664
rect 25004 22692 25010 22704
rect 25409 22695 25467 22701
rect 25409 22692 25421 22695
rect 25004 22664 25421 22692
rect 25004 22652 25010 22664
rect 25409 22661 25421 22664
rect 25455 22661 25467 22695
rect 25409 22655 25467 22661
rect 24765 22627 24823 22633
rect 24765 22593 24777 22627
rect 24811 22593 24823 22627
rect 24765 22587 24823 22593
rect 24854 22584 24860 22636
rect 24912 22584 24918 22636
rect 25038 22584 25044 22636
rect 25096 22584 25102 22636
rect 25222 22584 25228 22636
rect 25280 22584 25286 22636
rect 28810 22584 28816 22636
rect 28868 22584 28874 22636
rect 24210 22516 24216 22568
rect 24268 22556 24274 22568
rect 24673 22559 24731 22565
rect 24673 22556 24685 22559
rect 24268 22528 24685 22556
rect 24268 22516 24274 22528
rect 24673 22525 24685 22528
rect 24719 22556 24731 22559
rect 24719 22528 25176 22556
rect 24719 22525 24731 22528
rect 24673 22519 24731 22525
rect 21692 22460 23704 22488
rect 21692 22448 21698 22460
rect 24026 22448 24032 22500
rect 24084 22448 24090 22500
rect 24946 22488 24952 22500
rect 24320 22460 24952 22488
rect 15562 22420 15568 22432
rect 14936 22392 15568 22420
rect 15562 22380 15568 22392
rect 15620 22420 15626 22432
rect 15838 22420 15844 22432
rect 15620 22392 15844 22420
rect 15620 22380 15626 22392
rect 15838 22380 15844 22392
rect 15896 22380 15902 22432
rect 21082 22380 21088 22432
rect 21140 22380 21146 22432
rect 21542 22380 21548 22432
rect 21600 22380 21606 22432
rect 21821 22423 21879 22429
rect 21821 22389 21833 22423
rect 21867 22420 21879 22423
rect 22094 22420 22100 22432
rect 21867 22392 22100 22420
rect 21867 22389 21879 22392
rect 21821 22383 21879 22389
rect 22094 22380 22100 22392
rect 22152 22380 22158 22432
rect 22738 22380 22744 22432
rect 22796 22380 22802 22432
rect 22830 22380 22836 22432
rect 22888 22420 22894 22432
rect 23198 22420 23204 22432
rect 22888 22392 23204 22420
rect 22888 22380 22894 22392
rect 23198 22380 23204 22392
rect 23256 22380 23262 22432
rect 23477 22423 23535 22429
rect 23477 22389 23489 22423
rect 23523 22420 23535 22423
rect 24320 22420 24348 22460
rect 24946 22448 24952 22460
rect 25004 22448 25010 22500
rect 25148 22488 25176 22528
rect 25590 22516 25596 22568
rect 25648 22516 25654 22568
rect 25608 22488 25636 22516
rect 25148 22460 25636 22488
rect 28994 22448 29000 22500
rect 29052 22448 29058 22500
rect 23523 22392 24348 22420
rect 23523 22389 23535 22392
rect 23477 22383 23535 22389
rect 1104 22330 29440 22352
rect 1104 22278 4491 22330
rect 4543 22278 4555 22330
rect 4607 22278 4619 22330
rect 4671 22278 4683 22330
rect 4735 22278 4747 22330
rect 4799 22278 11574 22330
rect 11626 22278 11638 22330
rect 11690 22278 11702 22330
rect 11754 22278 11766 22330
rect 11818 22278 11830 22330
rect 11882 22278 18657 22330
rect 18709 22278 18721 22330
rect 18773 22278 18785 22330
rect 18837 22278 18849 22330
rect 18901 22278 18913 22330
rect 18965 22278 25740 22330
rect 25792 22278 25804 22330
rect 25856 22278 25868 22330
rect 25920 22278 25932 22330
rect 25984 22278 25996 22330
rect 26048 22278 29440 22330
rect 1104 22256 29440 22278
rect 6260 22219 6318 22225
rect 6260 22185 6272 22219
rect 6306 22216 6318 22219
rect 7282 22216 7288 22228
rect 6306 22188 7288 22216
rect 6306 22185 6318 22188
rect 6260 22179 6318 22185
rect 7282 22176 7288 22188
rect 7340 22176 7346 22228
rect 7650 22176 7656 22228
rect 7708 22216 7714 22228
rect 7745 22219 7803 22225
rect 7745 22216 7757 22219
rect 7708 22188 7757 22216
rect 7708 22176 7714 22188
rect 7745 22185 7757 22188
rect 7791 22185 7803 22219
rect 7745 22179 7803 22185
rect 8662 22176 8668 22228
rect 8720 22216 8726 22228
rect 8720 22188 10549 22216
rect 8720 22176 8726 22188
rect 8110 22148 8116 22160
rect 7300 22120 8116 22148
rect 7300 22092 7328 22120
rect 8110 22108 8116 22120
rect 8168 22108 8174 22160
rect 10521 22148 10549 22188
rect 10594 22176 10600 22228
rect 10652 22216 10658 22228
rect 11146 22216 11152 22228
rect 10652 22188 11152 22216
rect 10652 22176 10658 22188
rect 11146 22176 11152 22188
rect 11204 22216 11210 22228
rect 12618 22216 12624 22228
rect 11204 22188 12624 22216
rect 11204 22176 11210 22188
rect 12618 22176 12624 22188
rect 12676 22176 12682 22228
rect 14724 22219 14782 22225
rect 14724 22185 14736 22219
rect 14770 22216 14782 22219
rect 14826 22216 14832 22228
rect 14770 22188 14832 22216
rect 14770 22185 14782 22188
rect 14724 22179 14782 22185
rect 14826 22176 14832 22188
rect 14884 22176 14890 22228
rect 21358 22216 21364 22228
rect 21192 22188 21364 22216
rect 12526 22148 12532 22160
rect 9232 22120 10456 22148
rect 10521 22120 12532 22148
rect 5994 22040 6000 22092
rect 6052 22080 6058 22092
rect 6362 22080 6368 22092
rect 6052 22052 6368 22080
rect 6052 22040 6058 22052
rect 6362 22040 6368 22052
rect 6420 22040 6426 22092
rect 7282 22040 7288 22092
rect 7340 22040 7346 22092
rect 4246 21972 4252 22024
rect 4304 21972 4310 22024
rect 4525 22015 4583 22021
rect 4525 21981 4537 22015
rect 4571 21981 4583 22015
rect 4525 21975 4583 21981
rect 4430 21904 4436 21956
rect 4488 21944 4494 21956
rect 4540 21944 4568 21975
rect 5350 21972 5356 22024
rect 5408 21972 5414 22024
rect 5442 21972 5448 22024
rect 5500 21972 5506 22024
rect 5902 21972 5908 22024
rect 5960 21972 5966 22024
rect 7837 22015 7895 22021
rect 7837 21981 7849 22015
rect 7883 21981 7895 22015
rect 7837 21975 7895 21981
rect 9033 22015 9091 22021
rect 9033 21981 9045 22015
rect 9079 22012 9091 22015
rect 9232 22012 9260 22120
rect 9324 22052 9904 22080
rect 9324 22021 9352 22052
rect 9079 21984 9260 22012
rect 9309 22015 9367 22021
rect 9079 21981 9091 21984
rect 9033 21975 9091 21981
rect 9309 21981 9321 22015
rect 9355 21981 9367 22015
rect 9309 21975 9367 21981
rect 5460 21944 5488 21972
rect 4488 21916 5488 21944
rect 5736 21916 6762 21944
rect 4488 21904 4494 21916
rect 3326 21836 3332 21888
rect 3384 21876 3390 21888
rect 4062 21876 4068 21888
rect 3384 21848 4068 21876
rect 3384 21836 3390 21848
rect 4062 21836 4068 21848
rect 4120 21836 4126 21888
rect 4522 21836 4528 21888
rect 4580 21876 4586 21888
rect 5166 21876 5172 21888
rect 4580 21848 5172 21876
rect 4580 21836 4586 21848
rect 5166 21836 5172 21848
rect 5224 21876 5230 21888
rect 5736 21876 5764 21916
rect 5224 21848 5764 21876
rect 6656 21876 6684 21916
rect 7852 21888 7880 21975
rect 9398 21972 9404 22024
rect 9456 21972 9462 22024
rect 9677 22015 9735 22021
rect 9677 21981 9689 22015
rect 9723 21981 9735 22015
rect 9677 21975 9735 21981
rect 8386 21904 8392 21956
rect 8444 21944 8450 21956
rect 8846 21944 8852 21956
rect 8444 21916 8852 21944
rect 8444 21904 8450 21916
rect 8846 21904 8852 21916
rect 8904 21944 8910 21956
rect 9217 21947 9275 21953
rect 9217 21944 9229 21947
rect 8904 21916 9229 21944
rect 8904 21904 8910 21916
rect 9217 21913 9229 21916
rect 9263 21944 9275 21947
rect 9490 21944 9496 21956
rect 9263 21916 9496 21944
rect 9263 21913 9275 21916
rect 9217 21907 9275 21913
rect 9490 21904 9496 21916
rect 9548 21904 9554 21956
rect 7098 21876 7104 21888
rect 6656 21848 7104 21876
rect 5224 21836 5230 21848
rect 7098 21836 7104 21848
rect 7156 21836 7162 21888
rect 7834 21836 7840 21888
rect 7892 21836 7898 21888
rect 8478 21836 8484 21888
rect 8536 21836 8542 21888
rect 8570 21836 8576 21888
rect 8628 21876 8634 21888
rect 9398 21876 9404 21888
rect 8628 21848 9404 21876
rect 8628 21836 8634 21848
rect 9398 21836 9404 21848
rect 9456 21836 9462 21888
rect 9585 21879 9643 21885
rect 9585 21845 9597 21879
rect 9631 21876 9643 21879
rect 9692 21876 9720 21975
rect 9876 21944 9904 22052
rect 9950 22040 9956 22092
rect 10008 22040 10014 22092
rect 10428 22080 10456 22120
rect 12526 22108 12532 22120
rect 12584 22108 12590 22160
rect 20346 22108 20352 22160
rect 20404 22108 20410 22160
rect 21192 22148 21220 22188
rect 21358 22176 21364 22188
rect 21416 22176 21422 22228
rect 21634 22176 21640 22228
rect 21692 22176 21698 22228
rect 21726 22176 21732 22228
rect 21784 22216 21790 22228
rect 22097 22219 22155 22225
rect 21784 22188 22064 22216
rect 21784 22176 21790 22188
rect 21100 22120 21220 22148
rect 10428 22052 10640 22080
rect 9968 22012 9996 22040
rect 10321 22015 10379 22021
rect 10321 22012 10333 22015
rect 9968 21984 10333 22012
rect 10321 21981 10333 21984
rect 10367 21981 10379 22015
rect 10321 21975 10379 21981
rect 10413 22015 10471 22021
rect 10413 21981 10425 22015
rect 10459 21981 10471 22015
rect 10413 21975 10471 21981
rect 10226 21944 10232 21956
rect 9876 21916 10232 21944
rect 10226 21904 10232 21916
rect 10284 21904 10290 21956
rect 10428 21944 10456 21975
rect 10502 21972 10508 22024
rect 10560 21972 10566 22024
rect 10612 21956 10640 22052
rect 14458 22040 14464 22092
rect 14516 22080 14522 22092
rect 16482 22080 16488 22092
rect 14516 22052 16488 22080
rect 14516 22040 14522 22052
rect 16482 22040 16488 22052
rect 16540 22040 16546 22092
rect 18046 22080 18052 22092
rect 17236 22052 18052 22080
rect 17236 22024 17264 22052
rect 18046 22040 18052 22052
rect 18104 22080 18110 22092
rect 19242 22080 19248 22092
rect 18104 22052 19248 22080
rect 18104 22040 18110 22052
rect 19242 22040 19248 22052
rect 19300 22040 19306 22092
rect 20165 22083 20223 22089
rect 20165 22049 20177 22083
rect 20211 22080 20223 22083
rect 21100 22080 21128 22120
rect 21266 22108 21272 22160
rect 21324 22148 21330 22160
rect 22036 22148 22064 22188
rect 22097 22185 22109 22219
rect 22143 22216 22155 22219
rect 22554 22216 22560 22228
rect 22143 22188 22560 22216
rect 22143 22185 22155 22188
rect 22097 22179 22155 22185
rect 22554 22176 22560 22188
rect 22612 22176 22618 22228
rect 23753 22219 23811 22225
rect 23753 22185 23765 22219
rect 23799 22216 23811 22219
rect 24210 22216 24216 22228
rect 23799 22188 24216 22216
rect 23799 22185 23811 22188
rect 23753 22179 23811 22185
rect 24210 22176 24216 22188
rect 24268 22176 24274 22228
rect 24670 22176 24676 22228
rect 24728 22176 24734 22228
rect 24762 22176 24768 22228
rect 24820 22176 24826 22228
rect 22465 22151 22523 22157
rect 22465 22148 22477 22151
rect 21324 22120 21956 22148
rect 22036 22120 22477 22148
rect 21324 22108 21330 22120
rect 20211 22052 21128 22080
rect 20211 22049 20223 22052
rect 20165 22043 20223 22049
rect 10778 21972 10784 22024
rect 10836 21972 10842 22024
rect 10919 22015 10977 22021
rect 10919 21981 10931 22015
rect 10965 22012 10977 22015
rect 11974 22012 11980 22024
rect 10965 21984 11980 22012
rect 10965 21981 10977 21984
rect 10919 21975 10977 21981
rect 11974 21972 11980 21984
rect 12032 21972 12038 22024
rect 17218 22012 17224 22024
rect 15870 21984 17224 22012
rect 17218 21972 17224 21984
rect 17276 21972 17282 22024
rect 17313 22015 17371 22021
rect 17313 21981 17325 22015
rect 17359 22012 17371 22015
rect 18414 22012 18420 22024
rect 17359 21984 18420 22012
rect 17359 21981 17371 21984
rect 17313 21975 17371 21981
rect 18414 21972 18420 21984
rect 18472 21972 18478 22024
rect 20073 22015 20131 22021
rect 20073 21981 20085 22015
rect 20119 21981 20131 22015
rect 20073 21975 20131 21981
rect 20257 22015 20315 22021
rect 20257 21981 20269 22015
rect 20303 22012 20315 22015
rect 20438 22012 20444 22024
rect 20303 21984 20444 22012
rect 20303 21981 20315 21984
rect 20257 21975 20315 21981
rect 10428 21916 10548 21944
rect 10520 21888 10548 21916
rect 10594 21904 10600 21956
rect 10652 21904 10658 21956
rect 10686 21904 10692 21956
rect 10744 21904 10750 21956
rect 10980 21916 12434 21944
rect 10980 21888 11008 21916
rect 9631 21848 9720 21876
rect 9631 21845 9643 21848
rect 9585 21839 9643 21845
rect 10502 21836 10508 21888
rect 10560 21836 10566 21888
rect 10962 21836 10968 21888
rect 11020 21836 11026 21888
rect 11057 21879 11115 21885
rect 11057 21845 11069 21879
rect 11103 21876 11115 21879
rect 12066 21876 12072 21888
rect 11103 21848 12072 21876
rect 11103 21845 11115 21848
rect 11057 21839 11115 21845
rect 12066 21836 12072 21848
rect 12124 21836 12130 21888
rect 12406 21876 12434 21916
rect 12618 21904 12624 21956
rect 12676 21944 12682 21956
rect 13354 21944 13360 21956
rect 12676 21916 13360 21944
rect 12676 21904 12682 21916
rect 13354 21904 13360 21916
rect 13412 21904 13418 21956
rect 20088 21944 20116 21975
rect 20438 21972 20444 21984
rect 20496 21972 20502 22024
rect 20533 22015 20591 22021
rect 20533 21981 20545 22015
rect 20579 22012 20591 22015
rect 20714 22012 20720 22024
rect 20579 21984 20720 22012
rect 20579 21981 20591 21984
rect 20533 21975 20591 21981
rect 20714 21972 20720 21984
rect 20772 21972 20778 22024
rect 20806 21972 20812 22024
rect 20864 21972 20870 22024
rect 20990 21972 20996 22024
rect 21048 21972 21054 22024
rect 21082 21972 21088 22024
rect 21140 21972 21146 22024
rect 21376 22021 21404 22120
rect 21361 22015 21419 22021
rect 21361 21981 21373 22015
rect 21407 21981 21419 22015
rect 21361 21975 21419 21981
rect 21450 21972 21456 22024
rect 21508 21972 21514 22024
rect 21542 21972 21548 22024
rect 21600 22012 21606 22024
rect 21928 22021 21956 22120
rect 22465 22117 22477 22120
rect 22511 22148 22523 22151
rect 23842 22148 23848 22160
rect 22511 22120 23848 22148
rect 22511 22117 22523 22120
rect 22465 22111 22523 22117
rect 23842 22108 23848 22120
rect 23900 22108 23906 22160
rect 23937 22151 23995 22157
rect 23937 22117 23949 22151
rect 23983 22148 23995 22151
rect 24302 22148 24308 22160
rect 23983 22120 24308 22148
rect 23983 22117 23995 22120
rect 23937 22111 23995 22117
rect 24302 22108 24308 22120
rect 24360 22108 24366 22160
rect 24688 22148 24716 22176
rect 24596 22120 24716 22148
rect 22554 22040 22560 22092
rect 22612 22040 22618 22092
rect 22997 22083 23055 22089
rect 22997 22080 23009 22083
rect 22664 22052 23009 22080
rect 21729 22015 21787 22021
rect 21729 22012 21741 22015
rect 21600 21984 21741 22012
rect 21600 21972 21606 21984
rect 21729 21981 21741 21984
rect 21775 21981 21787 22015
rect 21729 21975 21787 21981
rect 21913 22015 21971 22021
rect 21913 21981 21925 22015
rect 21959 21981 21971 22015
rect 21913 21975 21971 21981
rect 22094 21972 22100 22024
rect 22152 22012 22158 22024
rect 22664 22021 22692 22052
rect 22997 22049 23009 22052
rect 23043 22049 23055 22083
rect 22997 22043 23055 22049
rect 23382 22040 23388 22092
rect 23440 22040 23446 22092
rect 23566 22040 23572 22092
rect 23624 22040 23630 22092
rect 22373 22015 22431 22021
rect 22373 22012 22385 22015
rect 22152 21984 22385 22012
rect 22152 21972 22158 21984
rect 22373 21981 22385 21984
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 22649 22015 22707 22021
rect 22649 21981 22661 22015
rect 22695 21981 22707 22015
rect 22649 21975 22707 21981
rect 22833 22015 22891 22021
rect 22833 21981 22845 22015
rect 22879 22012 22891 22015
rect 22879 21984 23060 22012
rect 22879 21981 22891 21984
rect 22833 21975 22891 21981
rect 20824 21944 20852 21972
rect 20088 21916 20852 21944
rect 21008 21944 21036 21972
rect 21269 21947 21327 21953
rect 21269 21944 21281 21947
rect 21008 21916 21281 21944
rect 21269 21913 21281 21916
rect 21315 21913 21327 21947
rect 21269 21907 21327 21913
rect 21634 21904 21640 21956
rect 21692 21944 21698 21956
rect 21692 21916 22692 21944
rect 21692 21904 21698 21916
rect 12894 21876 12900 21888
rect 12406 21848 12900 21876
rect 12894 21836 12900 21848
rect 12952 21876 12958 21888
rect 13630 21876 13636 21888
rect 12952 21848 13636 21876
rect 12952 21836 12958 21848
rect 13630 21836 13636 21848
rect 13688 21836 13694 21888
rect 16209 21879 16267 21885
rect 16209 21845 16221 21879
rect 16255 21876 16267 21879
rect 16298 21876 16304 21888
rect 16255 21848 16304 21876
rect 16255 21845 16267 21848
rect 16209 21839 16267 21845
rect 16298 21836 16304 21848
rect 16356 21876 16362 21888
rect 16666 21876 16672 21888
rect 16356 21848 16672 21876
rect 16356 21836 16362 21848
rect 16666 21836 16672 21848
rect 16724 21836 16730 21888
rect 17862 21836 17868 21888
rect 17920 21836 17926 21888
rect 20438 21836 20444 21888
rect 20496 21876 20502 21888
rect 20717 21879 20775 21885
rect 20717 21876 20729 21879
rect 20496 21848 20729 21876
rect 20496 21836 20502 21848
rect 20717 21845 20729 21848
rect 20763 21876 20775 21879
rect 21652 21876 21680 21904
rect 20763 21848 21680 21876
rect 22189 21879 22247 21885
rect 20763 21845 20775 21848
rect 20717 21839 20775 21845
rect 22189 21845 22201 21879
rect 22235 21876 22247 21879
rect 22554 21876 22560 21888
rect 22235 21848 22560 21876
rect 22235 21845 22247 21848
rect 22189 21839 22247 21845
rect 22554 21836 22560 21848
rect 22612 21836 22618 21888
rect 22664 21876 22692 21916
rect 22922 21904 22928 21956
rect 22980 21904 22986 21956
rect 23032 21944 23060 21984
rect 23198 21972 23204 22024
rect 23256 22021 23262 22024
rect 23256 22012 23268 22021
rect 23477 22015 23535 22021
rect 23477 22012 23489 22015
rect 23256 21984 23489 22012
rect 23256 21975 23268 21984
rect 23477 21981 23489 21984
rect 23523 21981 23535 22015
rect 23477 21975 23535 21981
rect 23256 21972 23262 21975
rect 23584 21944 23612 22040
rect 23860 22022 23888 22108
rect 24596 22080 24624 22120
rect 24857 22083 24915 22089
rect 24857 22080 24869 22083
rect 24136 22052 24532 22080
rect 24596 22052 24869 22080
rect 23860 22021 23970 22022
rect 23860 22015 23985 22021
rect 23860 21994 23939 22015
rect 23927 21981 23939 21994
rect 23973 21981 23985 22015
rect 23927 21975 23985 21981
rect 23032 21916 23612 21944
rect 23845 21947 23903 21953
rect 23845 21913 23857 21947
rect 23891 21944 23903 21947
rect 24136 21944 24164 22052
rect 24504 22024 24532 22052
rect 24857 22049 24869 22052
rect 24903 22049 24915 22083
rect 25222 22080 25228 22092
rect 24857 22043 24915 22049
rect 24964 22052 25228 22080
rect 24213 22015 24271 22021
rect 24213 21981 24225 22015
rect 24259 21981 24271 22015
rect 24213 21975 24271 21981
rect 23891 21916 24164 21944
rect 24228 21944 24256 21975
rect 24486 21972 24492 22024
rect 24544 22012 24550 22024
rect 24581 22015 24639 22021
rect 24581 22012 24593 22015
rect 24544 21984 24593 22012
rect 24544 21972 24550 21984
rect 24581 21981 24593 21984
rect 24627 21981 24639 22015
rect 24581 21975 24639 21981
rect 24670 21972 24676 22024
rect 24728 22012 24734 22024
rect 24964 22012 24992 22052
rect 25222 22040 25228 22052
rect 25280 22080 25286 22092
rect 25280 22052 25452 22080
rect 25280 22040 25286 22052
rect 24728 21984 24992 22012
rect 24728 21972 24734 21984
rect 25038 21972 25044 22024
rect 25096 21972 25102 22024
rect 25130 21972 25136 22024
rect 25188 21972 25194 22024
rect 25424 22021 25452 22052
rect 25409 22015 25467 22021
rect 25409 21981 25421 22015
rect 25455 21981 25467 22015
rect 25409 21975 25467 21981
rect 25498 21972 25504 22024
rect 25556 22012 25562 22024
rect 25685 22015 25743 22021
rect 25685 22012 25697 22015
rect 25556 21984 25697 22012
rect 25556 21972 25562 21984
rect 25685 21981 25697 21984
rect 25731 21981 25743 22015
rect 25685 21975 25743 21981
rect 25961 22015 26019 22021
rect 25961 21981 25973 22015
rect 26007 21981 26019 22015
rect 25961 21975 26019 21981
rect 25056 21944 25084 21972
rect 25317 21947 25375 21953
rect 25317 21944 25329 21947
rect 24228 21916 24992 21944
rect 25056 21916 25329 21944
rect 23891 21913 23903 21916
rect 23845 21907 23903 21913
rect 23109 21879 23167 21885
rect 23109 21876 23121 21879
rect 22664 21848 23121 21876
rect 23109 21845 23121 21848
rect 23155 21845 23167 21879
rect 23109 21839 23167 21845
rect 23290 21836 23296 21888
rect 23348 21876 23354 21888
rect 23860 21876 23888 21907
rect 23348 21848 23888 21876
rect 24121 21879 24179 21885
rect 23348 21836 23354 21848
rect 24121 21845 24133 21879
rect 24167 21876 24179 21879
rect 24210 21876 24216 21888
rect 24167 21848 24216 21876
rect 24167 21845 24179 21848
rect 24121 21839 24179 21845
rect 24210 21836 24216 21848
rect 24268 21836 24274 21888
rect 24394 21836 24400 21888
rect 24452 21836 24458 21888
rect 24964 21885 24992 21916
rect 25317 21913 25329 21916
rect 25363 21913 25375 21947
rect 25976 21944 26004 21975
rect 28810 21972 28816 22024
rect 28868 21972 28874 22024
rect 25317 21907 25375 21913
rect 25424 21916 26004 21944
rect 24949 21879 25007 21885
rect 24949 21845 24961 21879
rect 24995 21876 25007 21879
rect 25424 21876 25452 21916
rect 24995 21848 25452 21876
rect 25501 21879 25559 21885
rect 24995 21845 25007 21848
rect 24949 21839 25007 21845
rect 25501 21845 25513 21879
rect 25547 21876 25559 21879
rect 25590 21876 25596 21888
rect 25547 21848 25596 21876
rect 25547 21845 25559 21848
rect 25501 21839 25559 21845
rect 25590 21836 25596 21848
rect 25648 21836 25654 21888
rect 25682 21836 25688 21888
rect 25740 21876 25746 21888
rect 25869 21879 25927 21885
rect 25869 21876 25881 21879
rect 25740 21848 25881 21876
rect 25740 21836 25746 21848
rect 25869 21845 25881 21848
rect 25915 21876 25927 21879
rect 28828 21876 28856 21972
rect 25915 21848 28856 21876
rect 25915 21845 25927 21848
rect 25869 21839 25927 21845
rect 1104 21786 29595 21808
rect 1104 21734 8032 21786
rect 8084 21734 8096 21786
rect 8148 21734 8160 21786
rect 8212 21734 8224 21786
rect 8276 21734 8288 21786
rect 8340 21734 15115 21786
rect 15167 21734 15179 21786
rect 15231 21734 15243 21786
rect 15295 21734 15307 21786
rect 15359 21734 15371 21786
rect 15423 21734 22198 21786
rect 22250 21734 22262 21786
rect 22314 21734 22326 21786
rect 22378 21734 22390 21786
rect 22442 21734 22454 21786
rect 22506 21734 29281 21786
rect 29333 21734 29345 21786
rect 29397 21734 29409 21786
rect 29461 21734 29473 21786
rect 29525 21734 29537 21786
rect 29589 21734 29595 21786
rect 1104 21712 29595 21734
rect 4154 21672 4160 21684
rect 3160 21644 4160 21672
rect 3160 21545 3188 21644
rect 4154 21632 4160 21644
rect 4212 21632 4218 21684
rect 4430 21632 4436 21684
rect 4488 21632 4494 21684
rect 5350 21632 5356 21684
rect 5408 21672 5414 21684
rect 5537 21675 5595 21681
rect 5537 21672 5549 21675
rect 5408 21644 5549 21672
rect 5408 21632 5414 21644
rect 5537 21641 5549 21644
rect 5583 21641 5595 21675
rect 5537 21635 5595 21641
rect 5902 21632 5908 21684
rect 5960 21632 5966 21684
rect 6178 21632 6184 21684
rect 6236 21632 6242 21684
rect 7926 21672 7932 21684
rect 6380 21644 7932 21672
rect 3326 21564 3332 21616
rect 3384 21564 3390 21616
rect 4448 21604 4476 21632
rect 3528 21576 4476 21604
rect 3145 21539 3203 21545
rect 3145 21505 3157 21539
rect 3191 21505 3203 21539
rect 3145 21499 3203 21505
rect 3418 21496 3424 21548
rect 3476 21496 3482 21548
rect 3528 21545 3556 21576
rect 4522 21564 4528 21616
rect 4580 21564 4586 21616
rect 3513 21539 3571 21545
rect 3513 21505 3525 21539
rect 3559 21505 3571 21539
rect 3513 21499 3571 21505
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21505 5687 21539
rect 5629 21499 5687 21505
rect 3789 21471 3847 21477
rect 3789 21437 3801 21471
rect 3835 21437 3847 21471
rect 3789 21431 3847 21437
rect 4065 21471 4123 21477
rect 4065 21437 4077 21471
rect 4111 21468 4123 21471
rect 5074 21468 5080 21480
rect 4111 21440 5080 21468
rect 4111 21437 4123 21440
rect 4065 21431 4123 21437
rect 3804 21344 3832 21431
rect 5074 21428 5080 21440
rect 5132 21428 5138 21480
rect 5644 21468 5672 21499
rect 5810 21496 5816 21548
rect 5868 21496 5874 21548
rect 5920 21545 5948 21632
rect 5905 21539 5963 21545
rect 5905 21505 5917 21539
rect 5951 21505 5963 21539
rect 5905 21499 5963 21505
rect 5994 21496 6000 21548
rect 6052 21496 6058 21548
rect 6380 21545 6408 21644
rect 7926 21632 7932 21644
rect 7984 21672 7990 21684
rect 9950 21672 9956 21684
rect 7984 21644 9956 21672
rect 7984 21632 7990 21644
rect 7098 21564 7104 21616
rect 7156 21564 7162 21616
rect 8386 21564 8392 21616
rect 8444 21564 8450 21616
rect 8478 21564 8484 21616
rect 8536 21564 8542 21616
rect 6365 21539 6423 21545
rect 6365 21505 6377 21539
rect 6411 21505 6423 21539
rect 6365 21499 6423 21505
rect 8202 21496 8208 21548
rect 8260 21496 8266 21548
rect 8570 21496 8576 21548
rect 8628 21496 8634 21548
rect 9048 21545 9076 21644
rect 9950 21632 9956 21644
rect 10008 21632 10014 21684
rect 14458 21672 14464 21684
rect 12912 21644 14464 21672
rect 10962 21604 10968 21616
rect 10534 21576 10968 21604
rect 10962 21564 10968 21576
rect 11020 21564 11026 21616
rect 12437 21607 12495 21613
rect 12437 21573 12449 21607
rect 12483 21604 12495 21607
rect 12483 21576 12848 21604
rect 12483 21573 12495 21576
rect 12437 21567 12495 21573
rect 9033 21539 9091 21545
rect 9033 21505 9045 21539
rect 9079 21505 9091 21539
rect 9033 21499 9091 21505
rect 12066 21496 12072 21548
rect 12124 21496 12130 21548
rect 12158 21496 12164 21548
rect 12216 21496 12222 21548
rect 12618 21545 12624 21548
rect 12345 21539 12403 21545
rect 12345 21505 12357 21539
rect 12391 21505 12403 21539
rect 12345 21499 12403 21505
rect 12575 21539 12624 21545
rect 12575 21505 12587 21539
rect 12621 21505 12624 21539
rect 12575 21499 12624 21505
rect 5718 21468 5724 21480
rect 5644 21440 5724 21468
rect 3694 21292 3700 21344
rect 3752 21292 3758 21344
rect 3786 21292 3792 21344
rect 3844 21292 3850 21344
rect 4062 21292 4068 21344
rect 4120 21332 4126 21344
rect 5644 21332 5672 21440
rect 5718 21428 5724 21440
rect 5776 21468 5782 21480
rect 6641 21471 6699 21477
rect 5776 21440 6500 21468
rect 5776 21428 5782 21440
rect 6472 21344 6500 21440
rect 6641 21437 6653 21471
rect 6687 21468 6699 21471
rect 9309 21471 9367 21477
rect 6687 21440 8800 21468
rect 6687 21437 6699 21440
rect 6641 21431 6699 21437
rect 7742 21360 7748 21412
rect 7800 21400 7806 21412
rect 8202 21400 8208 21412
rect 7800 21372 8208 21400
rect 7800 21360 7806 21372
rect 8202 21360 8208 21372
rect 8260 21360 8266 21412
rect 8772 21409 8800 21440
rect 9309 21437 9321 21471
rect 9355 21468 9367 21471
rect 10318 21468 10324 21480
rect 9355 21440 10324 21468
rect 9355 21437 9367 21440
rect 9309 21431 9367 21437
rect 10318 21428 10324 21440
rect 10376 21428 10382 21480
rect 12360 21468 12388 21499
rect 12618 21496 12624 21499
rect 12676 21496 12682 21548
rect 12710 21468 12716 21480
rect 12360 21440 12716 21468
rect 12710 21428 12716 21440
rect 12768 21428 12774 21480
rect 8757 21403 8815 21409
rect 8757 21369 8769 21403
rect 8803 21369 8815 21403
rect 8757 21363 8815 21369
rect 4120 21304 5672 21332
rect 4120 21292 4126 21304
rect 6454 21292 6460 21344
rect 6512 21292 6518 21344
rect 7374 21292 7380 21344
rect 7432 21332 7438 21344
rect 7834 21332 7840 21344
rect 7432 21304 7840 21332
rect 7432 21292 7438 21304
rect 7834 21292 7840 21304
rect 7892 21332 7898 21344
rect 8113 21335 8171 21341
rect 8113 21332 8125 21335
rect 7892 21304 8125 21332
rect 7892 21292 7898 21304
rect 8113 21301 8125 21304
rect 8159 21301 8171 21335
rect 8113 21295 8171 21301
rect 10778 21292 10784 21344
rect 10836 21292 10842 21344
rect 12618 21292 12624 21344
rect 12676 21332 12682 21344
rect 12713 21335 12771 21341
rect 12713 21332 12725 21335
rect 12676 21304 12725 21332
rect 12676 21292 12682 21304
rect 12713 21301 12725 21304
rect 12759 21301 12771 21335
rect 12820 21332 12848 21576
rect 12912 21545 12940 21644
rect 14458 21632 14464 21644
rect 14516 21632 14522 21684
rect 18414 21632 18420 21684
rect 18472 21632 18478 21684
rect 18509 21675 18567 21681
rect 18509 21641 18521 21675
rect 18555 21672 18567 21675
rect 18555 21644 20116 21672
rect 18555 21641 18567 21644
rect 18509 21635 18567 21641
rect 13630 21564 13636 21616
rect 13688 21564 13694 21616
rect 17218 21564 17224 21616
rect 17276 21604 17282 21616
rect 19610 21604 19616 21616
rect 17276 21576 17434 21604
rect 18800 21576 19616 21604
rect 17276 21564 17282 21576
rect 18800 21545 18828 21576
rect 19610 21564 19616 21576
rect 19668 21564 19674 21616
rect 12897 21539 12955 21545
rect 12897 21505 12909 21539
rect 12943 21505 12955 21539
rect 18785 21539 18843 21545
rect 18785 21536 18797 21539
rect 12897 21499 12955 21505
rect 18156 21508 18797 21536
rect 13173 21471 13231 21477
rect 13173 21437 13185 21471
rect 13219 21468 13231 21471
rect 13262 21468 13268 21480
rect 13219 21440 13268 21468
rect 13219 21437 13231 21440
rect 13173 21431 13231 21437
rect 13262 21428 13268 21440
rect 13320 21428 13326 21480
rect 16574 21428 16580 21480
rect 16632 21468 16638 21480
rect 16669 21471 16727 21477
rect 16669 21468 16681 21471
rect 16632 21440 16681 21468
rect 16632 21428 16638 21440
rect 16669 21437 16681 21440
rect 16715 21437 16727 21471
rect 16669 21431 16727 21437
rect 16942 21428 16948 21480
rect 17000 21428 17006 21480
rect 18156 21468 18184 21508
rect 18785 21505 18797 21508
rect 18831 21505 18843 21539
rect 18785 21499 18843 21505
rect 18877 21539 18935 21545
rect 18877 21505 18889 21539
rect 18923 21536 18935 21539
rect 19058 21536 19064 21548
rect 18923 21508 19064 21536
rect 18923 21505 18935 21508
rect 18877 21499 18935 21505
rect 19058 21496 19064 21508
rect 19116 21496 19122 21548
rect 19150 21496 19156 21548
rect 19208 21496 19214 21548
rect 19337 21539 19395 21545
rect 19337 21505 19349 21539
rect 19383 21536 19395 21539
rect 19426 21536 19432 21548
rect 19383 21508 19432 21536
rect 19383 21505 19395 21508
rect 19337 21499 19395 21505
rect 19426 21496 19432 21508
rect 19484 21496 19490 21548
rect 20088 21536 20116 21644
rect 20806 21632 20812 21684
rect 20864 21632 20870 21684
rect 21450 21672 21456 21684
rect 21284 21644 21456 21672
rect 20165 21607 20223 21613
rect 20165 21573 20177 21607
rect 20211 21604 20223 21607
rect 21284 21604 21312 21644
rect 21450 21632 21456 21644
rect 21508 21632 21514 21684
rect 21545 21675 21603 21681
rect 21545 21641 21557 21675
rect 21591 21672 21603 21675
rect 21634 21672 21640 21684
rect 21591 21644 21640 21672
rect 21591 21641 21603 21644
rect 21545 21635 21603 21641
rect 21634 21632 21640 21644
rect 21692 21632 21698 21684
rect 23290 21672 23296 21684
rect 22388 21644 23296 21672
rect 20211 21576 21312 21604
rect 20211 21573 20223 21576
rect 20165 21567 20223 21573
rect 21358 21564 21364 21616
rect 21416 21604 21422 21616
rect 21416 21576 22140 21604
rect 21416 21564 21422 21576
rect 21085 21539 21143 21545
rect 20088 21508 20760 21536
rect 17972 21440 18184 21468
rect 18693 21471 18751 21477
rect 12986 21332 12992 21344
rect 12820 21304 12992 21332
rect 12713 21295 12771 21301
rect 12986 21292 12992 21304
rect 13044 21332 13050 21344
rect 14645 21335 14703 21341
rect 14645 21332 14657 21335
rect 13044 21304 14657 21332
rect 13044 21292 13050 21304
rect 14645 21301 14657 21304
rect 14691 21301 14703 21335
rect 14645 21295 14703 21301
rect 14734 21292 14740 21344
rect 14792 21332 14798 21344
rect 17972 21332 18000 21440
rect 18693 21437 18705 21471
rect 18739 21437 18751 21471
rect 18693 21431 18751 21437
rect 18969 21471 19027 21477
rect 18969 21437 18981 21471
rect 19015 21468 19027 21471
rect 19702 21468 19708 21480
rect 19015 21440 19708 21468
rect 19015 21437 19027 21440
rect 18969 21431 19027 21437
rect 18708 21400 18736 21431
rect 19702 21428 19708 21440
rect 19760 21428 19766 21480
rect 20533 21471 20591 21477
rect 20533 21437 20545 21471
rect 20579 21437 20591 21471
rect 20533 21431 20591 21437
rect 20548 21400 20576 21431
rect 20622 21428 20628 21480
rect 20680 21428 20686 21480
rect 20732 21468 20760 21508
rect 21085 21505 21097 21539
rect 21131 21536 21143 21539
rect 21453 21539 21511 21545
rect 21453 21536 21465 21539
rect 21131 21508 21465 21536
rect 21131 21505 21143 21508
rect 21085 21499 21143 21505
rect 21453 21505 21465 21508
rect 21499 21505 21511 21539
rect 21453 21499 21511 21505
rect 21821 21539 21879 21545
rect 21821 21505 21833 21539
rect 21867 21505 21879 21539
rect 21821 21499 21879 21505
rect 21266 21468 21272 21480
rect 20732 21440 21272 21468
rect 21266 21428 21272 21440
rect 21324 21428 21330 21480
rect 21358 21428 21364 21480
rect 21416 21428 21422 21480
rect 18708 21372 19564 21400
rect 20548 21372 20668 21400
rect 19536 21344 19564 21372
rect 20640 21344 20668 21372
rect 20714 21360 20720 21412
rect 20772 21400 20778 21412
rect 20901 21403 20959 21409
rect 20901 21400 20913 21403
rect 20772 21372 20913 21400
rect 20772 21360 20778 21372
rect 20901 21369 20913 21372
rect 20947 21400 20959 21403
rect 20947 21372 21404 21400
rect 20947 21369 20959 21372
rect 20901 21363 20959 21369
rect 21376 21344 21404 21372
rect 14792 21304 18000 21332
rect 14792 21292 14798 21304
rect 19518 21292 19524 21344
rect 19576 21292 19582 21344
rect 20622 21292 20628 21344
rect 20680 21292 20686 21344
rect 21358 21292 21364 21344
rect 21416 21292 21422 21344
rect 21468 21332 21496 21499
rect 21836 21468 21864 21499
rect 22002 21496 22008 21548
rect 22060 21496 22066 21548
rect 22112 21545 22140 21576
rect 22388 21545 22416 21644
rect 23290 21632 23296 21644
rect 23348 21632 23354 21684
rect 23385 21675 23443 21681
rect 23385 21641 23397 21675
rect 23431 21672 23443 21675
rect 23474 21672 23480 21684
rect 23431 21644 23480 21672
rect 23431 21641 23443 21644
rect 23385 21635 23443 21641
rect 23474 21632 23480 21644
rect 23532 21632 23538 21684
rect 23661 21675 23719 21681
rect 23661 21641 23673 21675
rect 23707 21672 23719 21675
rect 24118 21672 24124 21684
rect 23707 21644 24124 21672
rect 23707 21641 23719 21644
rect 23661 21635 23719 21641
rect 24118 21632 24124 21644
rect 24176 21632 24182 21684
rect 22554 21564 22560 21616
rect 22612 21564 22618 21616
rect 22830 21564 22836 21616
rect 22888 21564 22894 21616
rect 24026 21604 24032 21616
rect 23400 21576 24032 21604
rect 22097 21539 22155 21545
rect 22097 21505 22109 21539
rect 22143 21505 22155 21539
rect 22097 21499 22155 21505
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 22465 21539 22523 21545
rect 22465 21505 22477 21539
rect 22511 21536 22523 21539
rect 22572 21536 22600 21564
rect 22511 21508 22600 21536
rect 22833 21539 22845 21564
rect 22879 21539 22891 21564
rect 22833 21533 22891 21539
rect 22511 21505 22523 21508
rect 22465 21499 22523 21505
rect 23400 21480 23428 21576
rect 23860 21545 23888 21576
rect 24026 21564 24032 21576
rect 24084 21604 24090 21616
rect 24854 21604 24860 21616
rect 24084 21576 24860 21604
rect 24084 21564 24090 21576
rect 24854 21564 24860 21576
rect 24912 21604 24918 21616
rect 25130 21604 25136 21616
rect 24912 21576 25136 21604
rect 24912 21564 24918 21576
rect 25130 21564 25136 21576
rect 25188 21564 25194 21616
rect 23845 21539 23903 21545
rect 23845 21505 23857 21539
rect 23891 21505 23903 21539
rect 23845 21499 23903 21505
rect 24305 21539 24363 21545
rect 24305 21505 24317 21539
rect 24351 21536 24363 21539
rect 24394 21536 24400 21548
rect 24351 21508 24400 21536
rect 24351 21505 24363 21508
rect 24305 21499 24363 21505
rect 24394 21496 24400 21508
rect 24452 21496 24458 21548
rect 24670 21496 24676 21548
rect 24728 21496 24734 21548
rect 24946 21496 24952 21548
rect 25004 21496 25010 21548
rect 25314 21496 25320 21548
rect 25372 21496 25378 21548
rect 25498 21496 25504 21548
rect 25556 21496 25562 21548
rect 26970 21496 26976 21548
rect 27028 21496 27034 21548
rect 27157 21539 27215 21545
rect 27157 21505 27169 21539
rect 27203 21536 27215 21539
rect 27522 21536 27528 21548
rect 27203 21508 27528 21536
rect 27203 21505 27215 21508
rect 27157 21499 27215 21505
rect 22189 21471 22247 21477
rect 22189 21468 22201 21471
rect 21836 21440 22201 21468
rect 22189 21437 22201 21440
rect 22235 21437 22247 21471
rect 22189 21431 22247 21437
rect 22554 21428 22560 21480
rect 22612 21428 22618 21480
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21437 22707 21471
rect 22649 21431 22707 21437
rect 21818 21360 21824 21412
rect 21876 21360 21882 21412
rect 22664 21400 22692 21431
rect 22922 21428 22928 21480
rect 22980 21428 22986 21480
rect 23382 21428 23388 21480
rect 23440 21428 23446 21480
rect 23474 21428 23480 21480
rect 23532 21428 23538 21480
rect 27172 21468 27200 21499
rect 27522 21496 27528 21508
rect 27580 21496 27586 21548
rect 27709 21539 27767 21545
rect 27709 21505 27721 21539
rect 27755 21536 27767 21539
rect 27798 21536 27804 21548
rect 27755 21508 27804 21536
rect 27755 21505 27767 21508
rect 27709 21499 27767 21505
rect 27798 21496 27804 21508
rect 27856 21496 27862 21548
rect 26252 21440 27200 21468
rect 26252 21412 26280 21440
rect 22830 21400 22836 21412
rect 22664 21372 22836 21400
rect 22830 21360 22836 21372
rect 22888 21360 22894 21412
rect 23198 21360 23204 21412
rect 23256 21360 23262 21412
rect 24397 21403 24455 21409
rect 24397 21369 24409 21403
rect 24443 21400 24455 21403
rect 26234 21400 26240 21412
rect 24443 21372 26240 21400
rect 24443 21369 24455 21372
rect 24397 21363 24455 21369
rect 26234 21360 26240 21372
rect 26292 21360 26298 21412
rect 27062 21360 27068 21412
rect 27120 21360 27126 21412
rect 22646 21332 22652 21344
rect 21468 21304 22652 21332
rect 22646 21292 22652 21304
rect 22704 21292 22710 21344
rect 23842 21292 23848 21344
rect 23900 21332 23906 21344
rect 24578 21332 24584 21344
rect 23900 21304 24584 21332
rect 23900 21292 23906 21304
rect 24578 21292 24584 21304
rect 24636 21292 24642 21344
rect 25317 21335 25375 21341
rect 25317 21301 25329 21335
rect 25363 21332 25375 21335
rect 27246 21332 27252 21344
rect 25363 21304 27252 21332
rect 25363 21301 25375 21304
rect 25317 21295 25375 21301
rect 27246 21292 27252 21304
rect 27304 21292 27310 21344
rect 27614 21292 27620 21344
rect 27672 21292 27678 21344
rect 1104 21242 29440 21264
rect 1104 21190 4491 21242
rect 4543 21190 4555 21242
rect 4607 21190 4619 21242
rect 4671 21190 4683 21242
rect 4735 21190 4747 21242
rect 4799 21190 11574 21242
rect 11626 21190 11638 21242
rect 11690 21190 11702 21242
rect 11754 21190 11766 21242
rect 11818 21190 11830 21242
rect 11882 21190 18657 21242
rect 18709 21190 18721 21242
rect 18773 21190 18785 21242
rect 18837 21190 18849 21242
rect 18901 21190 18913 21242
rect 18965 21190 25740 21242
rect 25792 21190 25804 21242
rect 25856 21190 25868 21242
rect 25920 21190 25932 21242
rect 25984 21190 25996 21242
rect 26048 21190 29440 21242
rect 1104 21168 29440 21190
rect 3694 21088 3700 21140
rect 3752 21128 3758 21140
rect 4046 21131 4104 21137
rect 4046 21128 4058 21131
rect 3752 21100 4058 21128
rect 3752 21088 3758 21100
rect 4046 21097 4058 21100
rect 4092 21097 4104 21131
rect 4046 21091 4104 21097
rect 5537 21131 5595 21137
rect 5537 21097 5549 21131
rect 5583 21128 5595 21131
rect 5626 21128 5632 21140
rect 5583 21100 5632 21128
rect 5583 21097 5595 21100
rect 5537 21091 5595 21097
rect 5626 21088 5632 21100
rect 5684 21088 5690 21140
rect 6362 21128 6368 21140
rect 5736 21100 6368 21128
rect 3786 20952 3792 21004
rect 3844 20992 3850 21004
rect 5736 20992 5764 21100
rect 6362 21088 6368 21100
rect 6420 21088 6426 21140
rect 10686 21128 10692 21140
rect 7530 21100 10692 21128
rect 7530 21060 7558 21100
rect 10686 21088 10692 21100
rect 10744 21128 10750 21140
rect 10744 21100 11744 21128
rect 10744 21088 10750 21100
rect 10502 21060 10508 21072
rect 3844 20964 5764 20992
rect 5828 21032 7558 21060
rect 3844 20952 3850 20964
rect 1854 20884 1860 20936
rect 1912 20924 1918 20936
rect 3804 20924 3832 20952
rect 5828 20936 5856 21032
rect 6012 20964 6224 20992
rect 1912 20896 3832 20924
rect 1912 20884 1918 20896
rect 5350 20884 5356 20936
rect 5408 20884 5414 20936
rect 5810 20884 5816 20936
rect 5868 20884 5874 20936
rect 6012 20933 6040 20964
rect 6196 20936 6224 20964
rect 5997 20927 6055 20933
rect 5997 20893 6009 20927
rect 6043 20893 6055 20927
rect 5997 20887 6055 20893
rect 6090 20927 6148 20933
rect 6090 20893 6102 20927
rect 6136 20893 6148 20927
rect 6090 20887 6148 20893
rect 5368 20856 5396 20884
rect 6104 20856 6132 20887
rect 6178 20884 6184 20936
rect 6236 20884 6242 20936
rect 6275 20933 6303 21032
rect 6273 20927 6331 20933
rect 6273 20893 6285 20927
rect 6319 20893 6331 20927
rect 6273 20887 6331 20893
rect 6503 20927 6561 20933
rect 6503 20893 6515 20927
rect 6549 20924 6561 20927
rect 6730 20924 6736 20936
rect 6549 20896 6736 20924
rect 6549 20893 6561 20896
rect 6503 20887 6561 20893
rect 6730 20884 6736 20896
rect 6788 20884 6794 20936
rect 7006 20884 7012 20936
rect 7064 20924 7070 20936
rect 7285 20927 7343 20933
rect 7285 20924 7297 20927
rect 7064 20896 7297 20924
rect 7064 20884 7070 20896
rect 7285 20893 7297 20896
rect 7331 20893 7343 20927
rect 7285 20887 7343 20893
rect 7374 20884 7380 20936
rect 7432 20884 7438 20936
rect 7530 20924 7558 21032
rect 9508 21032 10508 21060
rect 7530 20896 7604 20924
rect 4448 20828 4554 20856
rect 5368 20828 6132 20856
rect 6365 20859 6423 20865
rect 3510 20748 3516 20800
rect 3568 20788 3574 20800
rect 4338 20788 4344 20800
rect 3568 20760 4344 20788
rect 3568 20748 3574 20760
rect 4338 20748 4344 20760
rect 4396 20788 4402 20800
rect 4448 20788 4476 20828
rect 6365 20825 6377 20859
rect 6411 20825 6423 20859
rect 6748 20856 6776 20884
rect 7576 20865 7604 20896
rect 7650 20884 7656 20936
rect 7708 20884 7714 20936
rect 7750 20927 7808 20933
rect 7750 20893 7762 20927
rect 7796 20893 7808 20927
rect 7750 20887 7808 20893
rect 7561 20859 7619 20865
rect 6748 20828 7420 20856
rect 6365 20819 6423 20825
rect 4396 20760 4476 20788
rect 4396 20748 4402 20760
rect 5626 20748 5632 20800
rect 5684 20788 5690 20800
rect 6380 20788 6408 20819
rect 5684 20760 6408 20788
rect 6641 20791 6699 20797
rect 5684 20748 5690 20760
rect 6641 20757 6653 20791
rect 6687 20788 6699 20791
rect 6914 20788 6920 20800
rect 6687 20760 6920 20788
rect 6687 20757 6699 20760
rect 6641 20751 6699 20757
rect 6914 20748 6920 20760
rect 6972 20748 6978 20800
rect 7392 20788 7420 20828
rect 7561 20825 7573 20859
rect 7607 20825 7619 20859
rect 7561 20819 7619 20825
rect 7760 20788 7788 20887
rect 8478 20884 8484 20936
rect 8536 20924 8542 20936
rect 9508 20924 9536 21032
rect 10502 21020 10508 21032
rect 10560 21060 10566 21072
rect 10560 21032 11008 21060
rect 10560 21020 10566 21032
rect 9585 20995 9643 21001
rect 9585 20961 9597 20995
rect 9631 20992 9643 20995
rect 10778 20992 10784 21004
rect 9631 20964 10784 20992
rect 9631 20961 9643 20964
rect 9585 20955 9643 20961
rect 10778 20952 10784 20964
rect 10836 20952 10842 21004
rect 10042 20924 10048 20936
rect 8536 20896 10048 20924
rect 8536 20884 8542 20896
rect 10042 20884 10048 20896
rect 10100 20884 10106 20936
rect 10413 20927 10471 20933
rect 10413 20893 10425 20927
rect 10459 20924 10471 20927
rect 10870 20924 10876 20936
rect 10459 20896 10876 20924
rect 10459 20893 10471 20896
rect 10413 20887 10471 20893
rect 10870 20884 10876 20896
rect 10928 20884 10934 20936
rect 10980 20924 11008 21032
rect 11422 20924 11428 20936
rect 10980 20896 11428 20924
rect 11422 20884 11428 20896
rect 11480 20884 11486 20936
rect 11514 20884 11520 20936
rect 11572 20884 11578 20936
rect 11716 20933 11744 21100
rect 12618 21088 12624 21140
rect 12676 21128 12682 21140
rect 12676 21100 14688 21128
rect 12676 21088 12682 21100
rect 13446 21020 13452 21072
rect 13504 21060 13510 21072
rect 14660 21060 14688 21100
rect 14734 21088 14740 21140
rect 14792 21088 14798 21140
rect 16485 21131 16543 21137
rect 16485 21097 16497 21131
rect 16531 21128 16543 21131
rect 16942 21128 16948 21140
rect 16531 21100 16948 21128
rect 16531 21097 16543 21100
rect 16485 21091 16543 21097
rect 16942 21088 16948 21100
rect 17000 21088 17006 21140
rect 17862 21088 17868 21140
rect 17920 21088 17926 21140
rect 19150 21088 19156 21140
rect 19208 21088 19214 21140
rect 19518 21088 19524 21140
rect 19576 21088 19582 21140
rect 19610 21088 19616 21140
rect 19668 21088 19674 21140
rect 21192 21100 23060 21128
rect 13504 21032 14504 21060
rect 14660 21032 15884 21060
rect 13504 21020 13510 21032
rect 11790 20952 11796 21004
rect 11848 20992 11854 21004
rect 12161 20995 12219 21001
rect 12161 20992 12173 20995
rect 11848 20964 12173 20992
rect 11848 20952 11854 20964
rect 12161 20961 12173 20964
rect 12207 20961 12219 20995
rect 12161 20955 12219 20961
rect 12437 20995 12495 21001
rect 12437 20961 12449 20995
rect 12483 20992 12495 20995
rect 14274 20992 14280 21004
rect 12483 20964 14280 20992
rect 12483 20961 12495 20964
rect 12437 20955 12495 20961
rect 14274 20952 14280 20964
rect 14332 20952 14338 21004
rect 11701 20927 11759 20933
rect 11701 20893 11713 20927
rect 11747 20893 11759 20927
rect 11701 20887 11759 20893
rect 11890 20927 11948 20933
rect 11890 20893 11902 20927
rect 11936 20924 11948 20927
rect 14093 20927 14151 20933
rect 14093 20924 14105 20927
rect 11936 20896 12020 20924
rect 11936 20893 11948 20896
rect 11890 20887 11948 20893
rect 9950 20816 9956 20868
rect 10008 20856 10014 20868
rect 11146 20856 11152 20868
rect 10008 20828 11152 20856
rect 10008 20816 10014 20828
rect 11146 20816 11152 20828
rect 11204 20816 11210 20868
rect 11793 20859 11851 20865
rect 11793 20825 11805 20859
rect 11839 20825 11851 20859
rect 11793 20819 11851 20825
rect 7392 20760 7788 20788
rect 7929 20791 7987 20797
rect 7929 20757 7941 20791
rect 7975 20788 7987 20791
rect 8570 20788 8576 20800
rect 7975 20760 8576 20788
rect 7975 20757 7987 20760
rect 7929 20751 7987 20757
rect 8570 20748 8576 20760
rect 8628 20748 8634 20800
rect 10134 20748 10140 20800
rect 10192 20748 10198 20800
rect 10778 20748 10784 20800
rect 10836 20788 10842 20800
rect 11808 20788 11836 20819
rect 11992 20800 12020 20896
rect 13740 20896 14105 20924
rect 12894 20816 12900 20868
rect 12952 20816 12958 20868
rect 10836 20760 11836 20788
rect 10836 20748 10842 20760
rect 11974 20748 11980 20800
rect 12032 20748 12038 20800
rect 12069 20791 12127 20797
rect 12069 20757 12081 20791
rect 12115 20788 12127 20791
rect 13740 20788 13768 20896
rect 14093 20893 14105 20896
rect 14139 20893 14151 20927
rect 14093 20887 14151 20893
rect 14182 20884 14188 20936
rect 14240 20884 14246 20936
rect 14476 20924 14504 21032
rect 14558 20927 14616 20933
rect 14558 20924 14570 20927
rect 14476 20896 14570 20924
rect 14558 20893 14570 20896
rect 14604 20893 14616 20927
rect 14558 20887 14616 20893
rect 14829 20927 14887 20933
rect 14829 20893 14841 20927
rect 14875 20893 14887 20927
rect 14829 20887 14887 20893
rect 13814 20816 13820 20868
rect 13872 20856 13878 20868
rect 14369 20859 14427 20865
rect 14369 20856 14381 20859
rect 13872 20828 14381 20856
rect 13872 20816 13878 20828
rect 14369 20825 14381 20828
rect 14415 20825 14427 20859
rect 14369 20819 14427 20825
rect 14461 20859 14519 20865
rect 14461 20825 14473 20859
rect 14507 20856 14519 20859
rect 14844 20856 14872 20887
rect 14507 20828 14872 20856
rect 14507 20825 14519 20828
rect 14461 20819 14519 20825
rect 12115 20760 13768 20788
rect 13909 20791 13967 20797
rect 12115 20757 12127 20760
rect 12069 20751 12127 20757
rect 13909 20757 13921 20791
rect 13955 20788 13967 20791
rect 14476 20788 14504 20819
rect 13955 20760 14504 20788
rect 13955 20757 13967 20760
rect 13909 20751 13967 20757
rect 15470 20748 15476 20800
rect 15528 20748 15534 20800
rect 15856 20788 15884 21032
rect 17880 20992 17908 21088
rect 15948 20964 17908 20992
rect 18325 20995 18383 21001
rect 15948 20933 15976 20964
rect 18325 20961 18337 20995
rect 18371 20992 18383 20995
rect 18509 20995 18567 21001
rect 18509 20992 18521 20995
rect 18371 20964 18521 20992
rect 18371 20961 18383 20964
rect 18325 20955 18383 20961
rect 18509 20961 18521 20964
rect 18555 20992 18567 20995
rect 19168 20992 19196 21088
rect 18555 20964 19196 20992
rect 18555 20961 18567 20964
rect 18509 20955 18567 20961
rect 15933 20927 15991 20933
rect 15933 20893 15945 20927
rect 15979 20893 15991 20927
rect 15933 20887 15991 20893
rect 16022 20884 16028 20936
rect 16080 20924 16086 20936
rect 16209 20927 16267 20933
rect 16209 20924 16221 20927
rect 16080 20896 16221 20924
rect 16080 20884 16086 20896
rect 16209 20893 16221 20896
rect 16255 20893 16267 20927
rect 16209 20887 16267 20893
rect 16301 20927 16359 20933
rect 16301 20893 16313 20927
rect 16347 20924 16359 20927
rect 16482 20924 16488 20936
rect 16347 20896 16488 20924
rect 16347 20893 16359 20896
rect 16301 20887 16359 20893
rect 16482 20884 16488 20896
rect 16540 20884 16546 20936
rect 16574 20884 16580 20936
rect 16632 20884 16638 20936
rect 19334 20924 19340 20936
rect 17986 20896 19340 20924
rect 19334 20884 19340 20896
rect 19392 20884 19398 20936
rect 19536 20933 19564 21088
rect 19628 20933 19656 21088
rect 20530 21020 20536 21072
rect 20588 21060 20594 21072
rect 21192 21060 21220 21100
rect 20588 21032 21220 21060
rect 20588 21020 20594 21032
rect 19702 20952 19708 21004
rect 19760 20992 19766 21004
rect 19886 20992 19892 21004
rect 19760 20964 19892 20992
rect 19760 20952 19766 20964
rect 19886 20952 19892 20964
rect 19944 20992 19950 21004
rect 20349 20995 20407 21001
rect 20349 20992 20361 20995
rect 19944 20964 20361 20992
rect 19944 20952 19950 20964
rect 20349 20961 20361 20964
rect 20395 20961 20407 20995
rect 20349 20955 20407 20961
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20893 19579 20927
rect 19521 20887 19579 20893
rect 19613 20927 19671 20933
rect 19613 20893 19625 20927
rect 19659 20893 19671 20927
rect 19613 20887 19671 20893
rect 19794 20884 19800 20936
rect 19852 20924 19858 20936
rect 19981 20927 20039 20933
rect 19981 20924 19993 20927
rect 19852 20896 19993 20924
rect 19852 20884 19858 20896
rect 19981 20893 19993 20896
rect 20027 20893 20039 20927
rect 19981 20887 20039 20893
rect 16114 20816 16120 20868
rect 16172 20816 16178 20868
rect 16853 20859 16911 20865
rect 16853 20825 16865 20859
rect 16899 20856 16911 20859
rect 17126 20856 17132 20868
rect 16899 20828 17132 20856
rect 16899 20825 16911 20828
rect 16853 20819 16911 20825
rect 17126 20816 17132 20828
rect 17184 20816 17190 20868
rect 18138 20816 18144 20868
rect 18196 20856 18202 20868
rect 18966 20856 18972 20868
rect 18196 20828 18972 20856
rect 18196 20816 18202 20828
rect 18966 20816 18972 20828
rect 19024 20856 19030 20868
rect 19024 20828 19196 20856
rect 19024 20816 19030 20828
rect 18874 20788 18880 20800
rect 15856 20760 18880 20788
rect 18874 20748 18880 20760
rect 18932 20748 18938 20800
rect 19058 20748 19064 20800
rect 19116 20748 19122 20800
rect 19168 20788 19196 20828
rect 19242 20816 19248 20868
rect 19300 20856 19306 20868
rect 20548 20856 20576 21020
rect 20622 20884 20628 20936
rect 20680 20924 20686 20936
rect 21100 20933 21128 21032
rect 21450 21020 21456 21072
rect 21508 21060 21514 21072
rect 21508 21032 22416 21060
rect 21508 21020 21514 21032
rect 21177 20995 21235 21001
rect 21177 20961 21189 20995
rect 21223 20992 21235 20995
rect 21542 20992 21548 21004
rect 21223 20964 21548 20992
rect 21223 20961 21235 20964
rect 21177 20955 21235 20961
rect 21542 20952 21548 20964
rect 21600 20992 21606 21004
rect 22388 20992 22416 21032
rect 23032 21004 23060 21100
rect 23382 21088 23388 21140
rect 23440 21128 23446 21140
rect 23477 21131 23535 21137
rect 23477 21128 23489 21131
rect 23440 21100 23489 21128
rect 23440 21088 23446 21100
rect 23477 21097 23489 21100
rect 23523 21097 23535 21131
rect 23477 21091 23535 21097
rect 23934 21088 23940 21140
rect 23992 21128 23998 21140
rect 24210 21128 24216 21140
rect 23992 21100 24216 21128
rect 23992 21088 23998 21100
rect 24210 21088 24216 21100
rect 24268 21088 24274 21140
rect 25869 21131 25927 21137
rect 25869 21097 25881 21131
rect 25915 21128 25927 21131
rect 26142 21128 26148 21140
rect 25915 21100 26148 21128
rect 25915 21097 25927 21100
rect 25869 21091 25927 21097
rect 26142 21088 26148 21100
rect 26200 21088 26206 21140
rect 26970 21088 26976 21140
rect 27028 21128 27034 21140
rect 27065 21131 27123 21137
rect 27065 21128 27077 21131
rect 27028 21100 27077 21128
rect 27028 21088 27034 21100
rect 27065 21097 27077 21100
rect 27111 21128 27123 21131
rect 27801 21131 27859 21137
rect 27801 21128 27813 21131
rect 27111 21100 27813 21128
rect 27111 21097 27123 21100
rect 27065 21091 27123 21097
rect 27801 21097 27813 21100
rect 27847 21097 27859 21131
rect 27801 21091 27859 21097
rect 23293 21063 23351 21069
rect 23293 21029 23305 21063
rect 23339 21060 23351 21063
rect 23566 21060 23572 21072
rect 23339 21032 23572 21060
rect 23339 21029 23351 21032
rect 23293 21023 23351 21029
rect 23566 21020 23572 21032
rect 23624 21020 23630 21072
rect 27982 21060 27988 21072
rect 23676 21032 24992 21060
rect 21600 20964 22140 20992
rect 21600 20952 21606 20964
rect 22112 20936 22140 20964
rect 22388 20964 22784 20992
rect 20901 20927 20959 20933
rect 20901 20924 20913 20927
rect 20680 20896 20913 20924
rect 20680 20884 20686 20896
rect 20901 20893 20913 20896
rect 20947 20893 20959 20927
rect 20901 20887 20959 20893
rect 21085 20927 21143 20933
rect 21085 20893 21097 20927
rect 21131 20893 21143 20927
rect 21085 20887 21143 20893
rect 19300 20828 20576 20856
rect 20916 20856 20944 20887
rect 21266 20884 21272 20936
rect 21324 20884 21330 20936
rect 21358 20884 21364 20936
rect 21416 20924 21422 20936
rect 21453 20927 21511 20933
rect 21453 20924 21465 20927
rect 21416 20896 21465 20924
rect 21416 20884 21422 20896
rect 21453 20893 21465 20896
rect 21499 20893 21511 20927
rect 21453 20887 21511 20893
rect 21637 20927 21695 20933
rect 21637 20893 21649 20927
rect 21683 20924 21695 20927
rect 21726 20924 21732 20936
rect 21683 20896 21732 20924
rect 21683 20893 21695 20896
rect 21637 20887 21695 20893
rect 21726 20884 21732 20896
rect 21784 20884 21790 20936
rect 22094 20884 22100 20936
rect 22152 20884 22158 20936
rect 22388 20933 22416 20964
rect 22373 20927 22431 20933
rect 22373 20893 22385 20927
rect 22419 20893 22431 20927
rect 22373 20887 22431 20893
rect 22646 20884 22652 20936
rect 22704 20884 22710 20936
rect 22756 20924 22784 20964
rect 23014 20952 23020 21004
rect 23072 20992 23078 21004
rect 23676 20992 23704 21032
rect 23072 20964 23704 20992
rect 23860 20964 24164 20992
rect 23072 20952 23078 20964
rect 23201 20927 23259 20933
rect 22756 20896 23152 20924
rect 23014 20856 23020 20868
rect 20916 20828 23020 20856
rect 19300 20816 19306 20828
rect 23014 20816 23020 20828
rect 23072 20816 23078 20868
rect 23124 20856 23152 20896
rect 23201 20893 23213 20927
rect 23247 20924 23259 20927
rect 23661 20927 23719 20933
rect 23661 20924 23673 20927
rect 23247 20896 23673 20924
rect 23247 20893 23259 20896
rect 23201 20887 23259 20893
rect 23661 20893 23673 20896
rect 23707 20924 23719 20927
rect 23750 20924 23756 20936
rect 23707 20896 23756 20924
rect 23707 20893 23719 20896
rect 23661 20887 23719 20893
rect 23750 20884 23756 20896
rect 23808 20884 23814 20936
rect 23860 20933 23888 20964
rect 24136 20936 24164 20964
rect 23845 20927 23903 20933
rect 23845 20893 23857 20927
rect 23891 20893 23903 20927
rect 23845 20887 23903 20893
rect 23937 20927 23995 20933
rect 23937 20893 23949 20927
rect 23983 20893 23995 20927
rect 23937 20887 23995 20893
rect 23860 20856 23888 20887
rect 23124 20828 23888 20856
rect 19518 20788 19524 20800
rect 19168 20760 19524 20788
rect 19518 20748 19524 20760
rect 19576 20748 19582 20800
rect 22646 20748 22652 20800
rect 22704 20788 22710 20800
rect 23952 20788 23980 20887
rect 24118 20884 24124 20936
rect 24176 20884 24182 20936
rect 24964 20933 24992 21032
rect 27448 21032 27988 21060
rect 25225 20995 25283 21001
rect 25225 20961 25237 20995
rect 25271 20992 25283 20995
rect 25590 20992 25596 21004
rect 25271 20964 25596 20992
rect 25271 20961 25283 20964
rect 25225 20955 25283 20961
rect 25590 20952 25596 20964
rect 25648 20952 25654 21004
rect 26697 20995 26755 21001
rect 26697 20992 26709 20995
rect 26068 20964 26709 20992
rect 24949 20927 25007 20933
rect 24949 20893 24961 20927
rect 24995 20893 25007 20927
rect 24949 20887 25007 20893
rect 25314 20816 25320 20868
rect 25372 20856 25378 20868
rect 25869 20859 25927 20865
rect 25869 20856 25881 20859
rect 25372 20828 25881 20856
rect 25372 20816 25378 20828
rect 25869 20825 25881 20828
rect 25915 20825 25927 20859
rect 25869 20819 25927 20825
rect 24026 20788 24032 20800
rect 22704 20760 24032 20788
rect 22704 20748 22710 20760
rect 24026 20748 24032 20760
rect 24084 20748 24090 20800
rect 26068 20797 26096 20964
rect 26697 20961 26709 20964
rect 26743 20992 26755 20995
rect 27062 20992 27068 21004
rect 26743 20964 27068 20992
rect 26743 20961 26755 20964
rect 26697 20955 26755 20961
rect 27062 20952 27068 20964
rect 27120 20992 27126 21004
rect 27448 20992 27476 21032
rect 27982 21020 27988 21032
rect 28040 21020 28046 21072
rect 27120 20964 27476 20992
rect 27120 20952 27126 20964
rect 26145 20927 26203 20933
rect 26145 20893 26157 20927
rect 26191 20924 26203 20927
rect 26234 20924 26240 20936
rect 26191 20896 26240 20924
rect 26191 20893 26203 20896
rect 26145 20887 26203 20893
rect 26234 20884 26240 20896
rect 26292 20884 26298 20936
rect 26602 20884 26608 20936
rect 26660 20924 26666 20936
rect 27448 20933 27476 20964
rect 27522 20952 27528 21004
rect 27580 20952 27586 21004
rect 27617 20995 27675 21001
rect 27617 20961 27629 20995
rect 27663 20992 27675 20995
rect 27798 20992 27804 21004
rect 27663 20964 27804 20992
rect 27663 20961 27675 20964
rect 27617 20955 27675 20961
rect 27798 20952 27804 20964
rect 27856 20992 27862 21004
rect 28902 20992 28908 21004
rect 27856 20964 28908 20992
rect 27856 20952 27862 20964
rect 28902 20952 28908 20964
rect 28960 20952 28966 21004
rect 26789 20927 26847 20933
rect 26789 20924 26801 20927
rect 26660 20896 26801 20924
rect 26660 20884 26666 20896
rect 26789 20893 26801 20896
rect 26835 20893 26847 20927
rect 26789 20887 26847 20893
rect 27341 20927 27399 20933
rect 27341 20893 27353 20927
rect 27387 20893 27399 20927
rect 27341 20887 27399 20893
rect 27433 20927 27491 20933
rect 27433 20893 27445 20927
rect 27479 20893 27491 20927
rect 27540 20924 27568 20952
rect 27709 20927 27767 20933
rect 27709 20924 27721 20927
rect 27540 20896 27721 20924
rect 27433 20887 27491 20893
rect 27709 20893 27721 20896
rect 27755 20893 27767 20927
rect 28445 20927 28503 20933
rect 28445 20924 28457 20927
rect 27709 20887 27767 20893
rect 27816 20896 28457 20924
rect 27356 20856 27384 20887
rect 27816 20856 27844 20896
rect 28445 20893 28457 20896
rect 28491 20893 28503 20927
rect 28445 20887 28503 20893
rect 27356 20828 27844 20856
rect 27448 20800 27476 20828
rect 27982 20816 27988 20868
rect 28040 20856 28046 20868
rect 28261 20859 28319 20865
rect 28261 20856 28273 20859
rect 28040 20828 28273 20856
rect 28040 20816 28046 20828
rect 28261 20825 28273 20828
rect 28307 20825 28319 20859
rect 28261 20819 28319 20825
rect 25777 20791 25835 20797
rect 25777 20757 25789 20791
rect 25823 20788 25835 20791
rect 26053 20791 26111 20797
rect 26053 20788 26065 20791
rect 25823 20760 26065 20788
rect 25823 20757 25835 20760
rect 25777 20751 25835 20757
rect 26053 20757 26065 20760
rect 26099 20757 26111 20791
rect 26053 20751 26111 20757
rect 27430 20748 27436 20800
rect 27488 20748 27494 20800
rect 28166 20748 28172 20800
rect 28224 20748 28230 20800
rect 28534 20748 28540 20800
rect 28592 20788 28598 20800
rect 28629 20791 28687 20797
rect 28629 20788 28641 20791
rect 28592 20760 28641 20788
rect 28592 20748 28598 20760
rect 28629 20757 28641 20760
rect 28675 20757 28687 20791
rect 28629 20751 28687 20757
rect 1104 20698 29595 20720
rect 1104 20646 8032 20698
rect 8084 20646 8096 20698
rect 8148 20646 8160 20698
rect 8212 20646 8224 20698
rect 8276 20646 8288 20698
rect 8340 20646 15115 20698
rect 15167 20646 15179 20698
rect 15231 20646 15243 20698
rect 15295 20646 15307 20698
rect 15359 20646 15371 20698
rect 15423 20646 22198 20698
rect 22250 20646 22262 20698
rect 22314 20646 22326 20698
rect 22378 20646 22390 20698
rect 22442 20646 22454 20698
rect 22506 20646 29281 20698
rect 29333 20646 29345 20698
rect 29397 20646 29409 20698
rect 29461 20646 29473 20698
rect 29525 20646 29537 20698
rect 29589 20646 29595 20698
rect 1104 20624 29595 20646
rect 3970 20584 3976 20596
rect 3344 20556 3976 20584
rect 3344 20457 3372 20556
rect 3970 20544 3976 20556
rect 4028 20544 4034 20596
rect 6178 20544 6184 20596
rect 6236 20584 6242 20596
rect 7006 20584 7012 20596
rect 6236 20556 7012 20584
rect 6236 20544 6242 20556
rect 7006 20544 7012 20556
rect 7064 20584 7070 20596
rect 7064 20556 8340 20584
rect 7064 20544 7070 20556
rect 3418 20476 3424 20528
rect 3476 20516 3482 20528
rect 3605 20519 3663 20525
rect 3605 20516 3617 20519
rect 3476 20488 3617 20516
rect 3476 20476 3482 20488
rect 3605 20485 3617 20488
rect 3651 20516 3663 20519
rect 4062 20516 4068 20528
rect 3651 20488 4068 20516
rect 3651 20485 3663 20488
rect 3605 20479 3663 20485
rect 4062 20476 4068 20488
rect 4120 20476 4126 20528
rect 4246 20516 4252 20528
rect 4172 20488 4252 20516
rect 4172 20457 4200 20488
rect 4246 20476 4252 20488
rect 4304 20516 4310 20528
rect 4304 20488 5488 20516
rect 4304 20476 4310 20488
rect 3329 20451 3387 20457
rect 3329 20417 3341 20451
rect 3375 20417 3387 20451
rect 3329 20411 3387 20417
rect 3513 20451 3571 20457
rect 3513 20417 3525 20451
rect 3559 20417 3571 20451
rect 3513 20411 3571 20417
rect 3697 20451 3755 20457
rect 3697 20417 3709 20451
rect 3743 20417 3755 20451
rect 3697 20411 3755 20417
rect 4157 20451 4215 20457
rect 4157 20417 4169 20451
rect 4203 20417 4215 20451
rect 4157 20411 4215 20417
rect 4525 20451 4583 20457
rect 4525 20417 4537 20451
rect 4571 20448 4583 20451
rect 5350 20448 5356 20460
rect 4571 20420 5356 20448
rect 4571 20417 4583 20420
rect 4525 20411 4583 20417
rect 3528 20312 3556 20411
rect 3712 20380 3740 20411
rect 4540 20380 4568 20411
rect 5350 20408 5356 20420
rect 5408 20408 5414 20460
rect 3712 20352 4568 20380
rect 4709 20383 4767 20389
rect 4709 20349 4721 20383
rect 4755 20380 4767 20383
rect 4890 20380 4896 20392
rect 4755 20352 4896 20380
rect 4755 20349 4767 20352
rect 4709 20343 4767 20349
rect 4724 20312 4752 20343
rect 4890 20340 4896 20352
rect 4948 20340 4954 20392
rect 3528 20284 4752 20312
rect 3878 20204 3884 20256
rect 3936 20204 3942 20256
rect 5460 20244 5488 20488
rect 7098 20476 7104 20528
rect 7156 20476 7162 20528
rect 8312 20516 8340 20556
rect 8386 20544 8392 20596
rect 8444 20584 8450 20596
rect 11238 20584 11244 20596
rect 8444 20556 11244 20584
rect 8444 20544 8450 20556
rect 8478 20516 8484 20528
rect 8312 20488 8484 20516
rect 8478 20476 8484 20488
rect 8536 20476 8542 20528
rect 9968 20525 9996 20556
rect 11238 20544 11244 20556
rect 11296 20544 11302 20596
rect 14274 20544 14280 20596
rect 14332 20584 14338 20596
rect 14921 20587 14979 20593
rect 14921 20584 14933 20587
rect 14332 20556 14933 20584
rect 14332 20544 14338 20556
rect 14921 20553 14933 20556
rect 14967 20553 14979 20587
rect 14921 20547 14979 20553
rect 16942 20544 16948 20596
rect 17000 20544 17006 20596
rect 17037 20587 17095 20593
rect 17037 20553 17049 20587
rect 17083 20553 17095 20587
rect 19058 20584 19064 20596
rect 17037 20547 17095 20553
rect 17328 20556 19064 20584
rect 9953 20519 10011 20525
rect 9953 20485 9965 20519
rect 9999 20485 10011 20519
rect 9953 20479 10011 20485
rect 10226 20476 10232 20528
rect 10284 20516 10290 20528
rect 10505 20519 10563 20525
rect 10505 20516 10517 20519
rect 10284 20488 10517 20516
rect 10284 20476 10290 20488
rect 10505 20485 10517 20488
rect 10551 20485 10563 20519
rect 10505 20479 10563 20485
rect 10594 20476 10600 20528
rect 10652 20516 10658 20528
rect 12342 20516 12348 20528
rect 10652 20488 12348 20516
rect 10652 20476 10658 20488
rect 12342 20476 12348 20488
rect 12400 20476 12406 20528
rect 12802 20476 12808 20528
rect 12860 20476 12866 20528
rect 17052 20460 17080 20547
rect 9674 20408 9680 20460
rect 9732 20408 9738 20460
rect 9858 20408 9864 20460
rect 9916 20408 9922 20460
rect 10045 20451 10103 20457
rect 10045 20417 10057 20451
rect 10091 20417 10103 20451
rect 10045 20411 10103 20417
rect 6362 20340 6368 20392
rect 6420 20340 6426 20392
rect 6638 20340 6644 20392
rect 6696 20340 6702 20392
rect 8205 20383 8263 20389
rect 8205 20380 8217 20383
rect 8128 20352 8217 20380
rect 7098 20244 7104 20256
rect 5460 20216 7104 20244
rect 7098 20204 7104 20216
rect 7156 20204 7162 20256
rect 7190 20204 7196 20256
rect 7248 20244 7254 20256
rect 8128 20253 8156 20352
rect 8205 20349 8217 20352
rect 8251 20349 8263 20383
rect 10060 20380 10088 20411
rect 10134 20408 10140 20460
rect 10192 20448 10198 20460
rect 10321 20451 10379 20457
rect 10321 20448 10333 20451
rect 10192 20420 10333 20448
rect 10192 20408 10198 20420
rect 10321 20417 10333 20420
rect 10367 20417 10379 20451
rect 10321 20411 10379 20417
rect 10410 20408 10416 20460
rect 10468 20448 10474 20460
rect 10689 20451 10747 20457
rect 10689 20448 10701 20451
rect 10468 20420 10701 20448
rect 10468 20408 10474 20420
rect 10689 20417 10701 20420
rect 10735 20448 10747 20451
rect 10962 20448 10968 20460
rect 10735 20420 10968 20448
rect 10735 20417 10747 20420
rect 10689 20411 10747 20417
rect 10962 20408 10968 20420
rect 11020 20408 11026 20460
rect 11146 20408 11152 20460
rect 11204 20448 11210 20460
rect 11790 20448 11796 20460
rect 11204 20420 11796 20448
rect 11204 20408 11210 20420
rect 11790 20408 11796 20420
rect 11848 20408 11854 20460
rect 13725 20451 13783 20457
rect 13725 20417 13737 20451
rect 13771 20448 13783 20451
rect 14182 20448 14188 20460
rect 13771 20420 14188 20448
rect 13771 20417 13783 20420
rect 13725 20411 13783 20417
rect 10060 20352 11008 20380
rect 8205 20343 8263 20349
rect 8478 20272 8484 20324
rect 8536 20312 8542 20324
rect 10229 20315 10287 20321
rect 10229 20312 10241 20315
rect 8536 20284 10241 20312
rect 8536 20272 8542 20284
rect 10229 20281 10241 20284
rect 10275 20281 10287 20315
rect 10229 20275 10287 20281
rect 10318 20272 10324 20324
rect 10376 20312 10382 20324
rect 10873 20315 10931 20321
rect 10873 20312 10885 20315
rect 10376 20284 10885 20312
rect 10376 20272 10382 20284
rect 10873 20281 10885 20284
rect 10919 20281 10931 20315
rect 10873 20275 10931 20281
rect 8113 20247 8171 20253
rect 8113 20244 8125 20247
rect 7248 20216 8125 20244
rect 7248 20204 7254 20216
rect 8113 20213 8125 20216
rect 8159 20213 8171 20247
rect 8113 20207 8171 20213
rect 8202 20204 8208 20256
rect 8260 20244 8266 20256
rect 8849 20247 8907 20253
rect 8849 20244 8861 20247
rect 8260 20216 8861 20244
rect 8260 20204 8266 20216
rect 8849 20213 8861 20216
rect 8895 20213 8907 20247
rect 10980 20244 11008 20352
rect 12066 20340 12072 20392
rect 12124 20340 12130 20392
rect 12434 20340 12440 20392
rect 12492 20380 12498 20392
rect 13541 20383 13599 20389
rect 12492 20352 13124 20380
rect 12492 20340 12498 20352
rect 13096 20312 13124 20352
rect 13541 20349 13553 20383
rect 13587 20380 13599 20383
rect 13740 20380 13768 20411
rect 14182 20408 14188 20420
rect 14240 20408 14246 20460
rect 14369 20451 14427 20457
rect 14369 20417 14381 20451
rect 14415 20417 14427 20451
rect 14369 20411 14427 20417
rect 13587 20352 13768 20380
rect 14384 20380 14412 20411
rect 14550 20408 14556 20460
rect 14608 20408 14614 20460
rect 14642 20408 14648 20460
rect 14700 20408 14706 20460
rect 14734 20408 14740 20460
rect 14792 20408 14798 20460
rect 15470 20408 15476 20460
rect 15528 20408 15534 20460
rect 16482 20408 16488 20460
rect 16540 20408 16546 20460
rect 16850 20408 16856 20460
rect 16908 20408 16914 20460
rect 17034 20408 17040 20460
rect 17092 20408 17098 20460
rect 17218 20408 17224 20460
rect 17276 20408 17282 20460
rect 17328 20457 17356 20556
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 21361 20587 21419 20593
rect 21361 20553 21373 20587
rect 21407 20584 21419 20587
rect 22021 20587 22079 20593
rect 22021 20584 22033 20587
rect 21407 20556 22033 20584
rect 21407 20553 21419 20556
rect 21361 20547 21419 20553
rect 22021 20553 22033 20556
rect 22067 20553 22079 20587
rect 22021 20547 22079 20553
rect 22189 20587 22247 20593
rect 22189 20553 22201 20587
rect 22235 20584 22247 20587
rect 22554 20584 22560 20596
rect 22235 20556 22560 20584
rect 22235 20553 22247 20556
rect 22189 20547 22247 20553
rect 22554 20544 22560 20556
rect 22612 20544 22618 20596
rect 22646 20544 22652 20596
rect 22704 20544 22710 20596
rect 22830 20544 22836 20596
rect 22888 20544 22894 20596
rect 23109 20587 23167 20593
rect 23109 20553 23121 20587
rect 23155 20584 23167 20587
rect 23290 20584 23296 20596
rect 23155 20556 23296 20584
rect 23155 20553 23167 20556
rect 23109 20547 23167 20553
rect 23290 20544 23296 20556
rect 23348 20544 23354 20596
rect 23477 20587 23535 20593
rect 23477 20553 23489 20587
rect 23523 20584 23535 20587
rect 24670 20584 24676 20596
rect 23523 20556 24676 20584
rect 23523 20553 23535 20556
rect 23477 20547 23535 20553
rect 24670 20544 24676 20556
rect 24728 20544 24734 20596
rect 27062 20544 27068 20596
rect 27120 20544 27126 20596
rect 27540 20556 28764 20584
rect 17957 20519 18015 20525
rect 17957 20485 17969 20519
rect 18003 20516 18015 20519
rect 20993 20519 21051 20525
rect 18003 20488 19472 20516
rect 18003 20485 18015 20488
rect 17957 20479 18015 20485
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 17494 20408 17500 20460
rect 17552 20408 17558 20460
rect 17586 20408 17592 20460
rect 17644 20408 17650 20460
rect 17681 20451 17739 20457
rect 17681 20417 17693 20451
rect 17727 20417 17739 20451
rect 17681 20411 17739 20417
rect 15488 20380 15516 20408
rect 14384 20352 15516 20380
rect 16500 20380 16528 20408
rect 17696 20380 17724 20411
rect 18138 20408 18144 20460
rect 18196 20408 18202 20460
rect 18322 20408 18328 20460
rect 18380 20408 18386 20460
rect 18785 20451 18843 20457
rect 18785 20417 18797 20451
rect 18831 20417 18843 20451
rect 18785 20411 18843 20417
rect 16500 20352 17724 20380
rect 13587 20349 13599 20352
rect 13541 20343 13599 20349
rect 17954 20340 17960 20392
rect 18012 20380 18018 20392
rect 18417 20383 18475 20389
rect 18417 20380 18429 20383
rect 18012 20352 18429 20380
rect 18012 20340 18018 20352
rect 18417 20349 18429 20352
rect 18463 20380 18475 20383
rect 18800 20380 18828 20411
rect 18874 20408 18880 20460
rect 18932 20448 18938 20460
rect 19444 20457 19472 20488
rect 20993 20485 21005 20519
rect 21039 20516 21051 20519
rect 21542 20516 21548 20528
rect 21039 20488 21548 20516
rect 21039 20485 21051 20488
rect 20993 20479 21051 20485
rect 21542 20476 21548 20488
rect 21600 20476 21606 20528
rect 21821 20519 21879 20525
rect 21821 20485 21833 20519
rect 21867 20485 21879 20519
rect 21821 20479 21879 20485
rect 19153 20451 19211 20457
rect 19153 20448 19165 20451
rect 18932 20420 19165 20448
rect 18932 20408 18938 20420
rect 19153 20417 19165 20420
rect 19199 20417 19211 20451
rect 19153 20411 19211 20417
rect 19429 20451 19487 20457
rect 19429 20417 19441 20451
rect 19475 20417 19487 20451
rect 19429 20411 19487 20417
rect 21082 20408 21088 20460
rect 21140 20448 21146 20460
rect 21177 20451 21235 20457
rect 21177 20448 21189 20451
rect 21140 20420 21189 20448
rect 21140 20408 21146 20420
rect 21177 20417 21189 20420
rect 21223 20417 21235 20451
rect 21177 20411 21235 20417
rect 21453 20451 21511 20457
rect 21453 20417 21465 20451
rect 21499 20448 21511 20451
rect 21560 20448 21588 20476
rect 21499 20420 21588 20448
rect 21637 20451 21695 20457
rect 21499 20417 21511 20420
rect 21453 20411 21511 20417
rect 21637 20417 21649 20451
rect 21683 20417 21695 20451
rect 21637 20411 21695 20417
rect 20530 20380 20536 20392
rect 18463 20352 18736 20380
rect 18800 20352 20536 20380
rect 18463 20349 18475 20352
rect 18417 20343 18475 20349
rect 16669 20315 16727 20321
rect 13096 20284 14688 20312
rect 14660 20256 14688 20284
rect 16669 20281 16681 20315
rect 16715 20312 16727 20315
rect 18506 20312 18512 20324
rect 16715 20284 18512 20312
rect 16715 20281 16727 20284
rect 16669 20275 16727 20281
rect 18506 20272 18512 20284
rect 18564 20272 18570 20324
rect 13170 20244 13176 20256
rect 10980 20216 13176 20244
rect 8849 20207 8907 20213
rect 13170 20204 13176 20216
rect 13228 20204 13234 20256
rect 14274 20204 14280 20256
rect 14332 20204 14338 20256
rect 14642 20204 14648 20256
rect 14700 20204 14706 20256
rect 17126 20204 17132 20256
rect 17184 20244 17190 20256
rect 17865 20247 17923 20253
rect 17865 20244 17877 20247
rect 17184 20216 17877 20244
rect 17184 20204 17190 20216
rect 17865 20213 17877 20216
rect 17911 20213 17923 20247
rect 18708 20244 18736 20352
rect 20530 20340 20536 20352
rect 20588 20340 20594 20392
rect 21192 20380 21220 20411
rect 21542 20380 21548 20392
rect 21192 20352 21548 20380
rect 21542 20340 21548 20352
rect 21600 20380 21606 20392
rect 21652 20380 21680 20411
rect 21600 20352 21680 20380
rect 21600 20340 21606 20352
rect 18877 20315 18935 20321
rect 18877 20281 18889 20315
rect 18923 20312 18935 20315
rect 19242 20312 19248 20324
rect 18923 20284 19248 20312
rect 18923 20281 18935 20284
rect 18877 20275 18935 20281
rect 19242 20272 19248 20284
rect 19300 20272 19306 20324
rect 21266 20272 21272 20324
rect 21324 20312 21330 20324
rect 21836 20312 21864 20479
rect 22664 20448 22692 20544
rect 22848 20516 22876 20544
rect 24305 20519 24363 20525
rect 24305 20516 24317 20519
rect 22848 20488 24317 20516
rect 23676 20457 23704 20488
rect 24305 20485 24317 20488
rect 24351 20485 24363 20519
rect 24305 20479 24363 20485
rect 22925 20451 22983 20457
rect 22925 20448 22937 20451
rect 22664 20420 22937 20448
rect 22925 20417 22937 20420
rect 22971 20417 22983 20451
rect 22925 20411 22983 20417
rect 23661 20451 23719 20457
rect 23661 20417 23673 20451
rect 23707 20417 23719 20451
rect 23661 20411 23719 20417
rect 23750 20408 23756 20460
rect 23808 20408 23814 20460
rect 23845 20451 23903 20457
rect 23845 20417 23857 20451
rect 23891 20417 23903 20451
rect 23845 20411 23903 20417
rect 22002 20340 22008 20392
rect 22060 20380 22066 20392
rect 22741 20383 22799 20389
rect 22741 20380 22753 20383
rect 22060 20352 22753 20380
rect 22060 20340 22094 20352
rect 22741 20349 22753 20352
rect 22787 20380 22799 20383
rect 23768 20380 23796 20408
rect 22787 20352 23796 20380
rect 22787 20349 22799 20352
rect 22741 20343 22799 20349
rect 22066 20312 22094 20340
rect 21324 20284 22094 20312
rect 21324 20272 21330 20284
rect 23106 20272 23112 20324
rect 23164 20312 23170 20324
rect 23860 20312 23888 20411
rect 23934 20408 23940 20460
rect 23992 20408 23998 20460
rect 24026 20408 24032 20460
rect 24084 20408 24090 20460
rect 24118 20408 24124 20460
rect 24176 20408 24182 20460
rect 25314 20408 25320 20460
rect 25372 20448 25378 20460
rect 26602 20448 26608 20460
rect 25372 20420 26608 20448
rect 25372 20408 25378 20420
rect 26602 20408 26608 20420
rect 26660 20408 26666 20460
rect 27080 20457 27108 20544
rect 27540 20516 27568 20556
rect 28534 20516 28540 20528
rect 27356 20488 27568 20516
rect 27356 20460 27384 20488
rect 27065 20451 27123 20457
rect 27065 20417 27077 20451
rect 27111 20417 27123 20451
rect 27065 20411 27123 20417
rect 27338 20408 27344 20460
rect 27396 20408 27402 20460
rect 27430 20408 27436 20460
rect 27488 20408 27494 20460
rect 24305 20383 24363 20389
rect 24305 20349 24317 20383
rect 24351 20349 24363 20383
rect 24305 20343 24363 20349
rect 26697 20383 26755 20389
rect 26697 20349 26709 20383
rect 26743 20380 26755 20383
rect 27448 20380 27476 20408
rect 26743 20352 27476 20380
rect 27540 20380 27568 20488
rect 27908 20488 28540 20516
rect 27908 20457 27936 20488
rect 28534 20476 28540 20488
rect 28592 20476 28598 20528
rect 28540 20473 28598 20476
rect 27893 20451 27951 20457
rect 27893 20417 27905 20451
rect 27939 20417 27951 20451
rect 27893 20411 27951 20417
rect 27985 20451 28043 20457
rect 27985 20417 27997 20451
rect 28031 20417 28043 20451
rect 27985 20411 28043 20417
rect 28000 20380 28028 20411
rect 28074 20408 28080 20460
rect 28132 20448 28138 20460
rect 28169 20451 28227 20457
rect 28169 20448 28181 20451
rect 28132 20420 28181 20448
rect 28132 20408 28138 20420
rect 28169 20417 28181 20420
rect 28215 20417 28227 20451
rect 28169 20411 28227 20417
rect 28261 20451 28319 20457
rect 28261 20417 28273 20451
rect 28307 20417 28319 20451
rect 28540 20439 28552 20473
rect 28586 20439 28598 20473
rect 28540 20433 28598 20439
rect 28629 20451 28687 20457
rect 28261 20411 28319 20417
rect 28629 20417 28641 20451
rect 28675 20448 28687 20451
rect 28736 20448 28764 20556
rect 28675 20420 28764 20448
rect 28813 20451 28871 20457
rect 28675 20417 28687 20420
rect 28629 20411 28687 20417
rect 28813 20417 28825 20451
rect 28859 20417 28871 20451
rect 28813 20411 28871 20417
rect 27540 20352 28028 20380
rect 28276 20380 28304 20411
rect 28828 20380 28856 20411
rect 28902 20408 28908 20460
rect 28960 20408 28966 20460
rect 28276 20352 28856 20380
rect 26743 20349 26755 20352
rect 26697 20343 26755 20349
rect 23164 20284 23888 20312
rect 23164 20272 23170 20284
rect 19426 20244 19432 20256
rect 18708 20216 19432 20244
rect 17865 20207 17923 20213
rect 19426 20204 19432 20216
rect 19484 20204 19490 20256
rect 21545 20247 21603 20253
rect 21545 20213 21557 20247
rect 21591 20244 21603 20247
rect 22005 20247 22063 20253
rect 22005 20244 22017 20247
rect 21591 20216 22017 20244
rect 21591 20213 21603 20216
rect 21545 20207 21603 20213
rect 22005 20213 22017 20216
rect 22051 20213 22063 20247
rect 22005 20207 22063 20213
rect 23750 20204 23756 20256
rect 23808 20244 23814 20256
rect 24320 20244 24348 20343
rect 27246 20272 27252 20324
rect 27304 20312 27310 20324
rect 28276 20312 28304 20352
rect 27304 20284 28304 20312
rect 27304 20272 27310 20284
rect 23808 20216 24348 20244
rect 23808 20204 23814 20216
rect 27338 20204 27344 20256
rect 27396 20204 27402 20256
rect 27522 20204 27528 20256
rect 27580 20244 27586 20256
rect 27617 20247 27675 20253
rect 27617 20244 27629 20247
rect 27580 20216 27629 20244
rect 27580 20204 27586 20216
rect 27617 20213 27629 20216
rect 27663 20213 27675 20247
rect 27617 20207 27675 20213
rect 27706 20204 27712 20256
rect 27764 20204 27770 20256
rect 28350 20204 28356 20256
rect 28408 20204 28414 20256
rect 1104 20154 29440 20176
rect 1104 20102 4491 20154
rect 4543 20102 4555 20154
rect 4607 20102 4619 20154
rect 4671 20102 4683 20154
rect 4735 20102 4747 20154
rect 4799 20102 11574 20154
rect 11626 20102 11638 20154
rect 11690 20102 11702 20154
rect 11754 20102 11766 20154
rect 11818 20102 11830 20154
rect 11882 20102 18657 20154
rect 18709 20102 18721 20154
rect 18773 20102 18785 20154
rect 18837 20102 18849 20154
rect 18901 20102 18913 20154
rect 18965 20102 25740 20154
rect 25792 20102 25804 20154
rect 25856 20102 25868 20154
rect 25920 20102 25932 20154
rect 25984 20102 25996 20154
rect 26048 20102 29440 20154
rect 1104 20080 29440 20102
rect 3878 20000 3884 20052
rect 3936 20000 3942 20052
rect 3970 20000 3976 20052
rect 4028 20040 4034 20052
rect 4433 20043 4491 20049
rect 4433 20040 4445 20043
rect 4028 20012 4445 20040
rect 4028 20000 4034 20012
rect 4433 20009 4445 20012
rect 4479 20009 4491 20043
rect 4433 20003 4491 20009
rect 6638 20000 6644 20052
rect 6696 20040 6702 20052
rect 6917 20043 6975 20049
rect 6917 20040 6929 20043
rect 6696 20012 6929 20040
rect 6696 20000 6702 20012
rect 6917 20009 6929 20012
rect 6963 20009 6975 20043
rect 8202 20040 8208 20052
rect 6917 20003 6975 20009
rect 7024 20012 8208 20040
rect 2133 19907 2191 19913
rect 2133 19873 2145 19907
rect 2179 19904 2191 19907
rect 3896 19904 3924 20000
rect 7024 19904 7052 20012
rect 8202 20000 8208 20012
rect 8260 20000 8266 20052
rect 8757 20043 8815 20049
rect 8757 20009 8769 20043
rect 8803 20040 8815 20043
rect 9674 20040 9680 20052
rect 8803 20012 9680 20040
rect 8803 20009 8815 20012
rect 8757 20003 8815 20009
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 12066 20000 12072 20052
rect 12124 20040 12130 20052
rect 12621 20043 12679 20049
rect 12621 20040 12633 20043
rect 12124 20012 12633 20040
rect 12124 20000 12130 20012
rect 12621 20009 12633 20012
rect 12667 20009 12679 20043
rect 12621 20003 12679 20009
rect 16117 20043 16175 20049
rect 16117 20009 16129 20043
rect 16163 20040 16175 20043
rect 16850 20040 16856 20052
rect 16163 20012 16856 20040
rect 16163 20009 16175 20012
rect 16117 20003 16175 20009
rect 16850 20000 16856 20012
rect 16908 20000 16914 20052
rect 17034 20000 17040 20052
rect 17092 20040 17098 20052
rect 18138 20040 18144 20052
rect 17092 20012 18144 20040
rect 17092 20000 17098 20012
rect 18138 20000 18144 20012
rect 18196 20000 18202 20052
rect 18506 20000 18512 20052
rect 18564 20040 18570 20052
rect 22646 20040 22652 20052
rect 18564 20012 22652 20040
rect 18564 20000 18570 20012
rect 22646 20000 22652 20012
rect 22704 20000 22710 20052
rect 27617 20043 27675 20049
rect 27617 20009 27629 20043
rect 27663 20040 27675 20043
rect 28074 20040 28080 20052
rect 27663 20012 28080 20040
rect 27663 20009 27675 20012
rect 27617 20003 27675 20009
rect 28074 20000 28080 20012
rect 28132 20000 28138 20052
rect 9398 19972 9404 19984
rect 2179 19876 3924 19904
rect 6380 19876 7052 19904
rect 7760 19944 9404 19972
rect 2179 19873 2191 19876
rect 2133 19867 2191 19873
rect 1854 19796 1860 19848
rect 1912 19796 1918 19848
rect 6380 19845 6408 19876
rect 3881 19839 3939 19845
rect 3881 19805 3893 19839
rect 3927 19805 3939 19839
rect 3881 19799 3939 19805
rect 6365 19839 6423 19845
rect 6365 19805 6377 19839
rect 6411 19805 6423 19839
rect 6365 19799 6423 19805
rect 3418 19768 3424 19780
rect 3358 19740 3424 19768
rect 3418 19728 3424 19740
rect 3476 19728 3482 19780
rect 3605 19703 3663 19709
rect 3605 19669 3617 19703
rect 3651 19700 3663 19703
rect 3896 19700 3924 19799
rect 6454 19796 6460 19848
rect 6512 19836 6518 19848
rect 6641 19839 6699 19845
rect 6641 19836 6653 19839
rect 6512 19808 6653 19836
rect 6512 19796 6518 19808
rect 6641 19805 6653 19808
rect 6687 19805 6699 19839
rect 6641 19799 6699 19805
rect 6733 19839 6791 19845
rect 6733 19805 6745 19839
rect 6779 19836 6791 19839
rect 6822 19836 6828 19848
rect 6779 19808 6828 19836
rect 6779 19805 6791 19808
rect 6733 19799 6791 19805
rect 6822 19796 6828 19808
rect 6880 19796 6886 19848
rect 6914 19796 6920 19848
rect 6972 19836 6978 19848
rect 7190 19845 7196 19848
rect 7009 19839 7067 19845
rect 7009 19836 7021 19839
rect 6972 19808 7021 19836
rect 6972 19796 6978 19808
rect 7009 19805 7021 19808
rect 7055 19805 7067 19839
rect 7009 19799 7067 19805
rect 7157 19839 7196 19845
rect 7157 19805 7169 19839
rect 7157 19799 7196 19805
rect 7190 19796 7196 19799
rect 7248 19796 7254 19848
rect 7515 19839 7573 19845
rect 7515 19805 7527 19839
rect 7561 19836 7573 19839
rect 7760 19836 7788 19944
rect 9398 19932 9404 19944
rect 9456 19932 9462 19984
rect 12434 19972 12440 19984
rect 10796 19944 12440 19972
rect 10796 19904 10824 19944
rect 7852 19876 10824 19904
rect 7852 19848 7880 19876
rect 7561 19808 7788 19836
rect 7561 19805 7573 19808
rect 7515 19799 7573 19805
rect 7834 19796 7840 19848
rect 7892 19796 7898 19848
rect 8205 19839 8263 19845
rect 8205 19805 8217 19839
rect 8251 19836 8263 19839
rect 8846 19836 8852 19848
rect 8251 19808 8852 19836
rect 8251 19805 8263 19808
rect 8205 19799 8263 19805
rect 8846 19796 8852 19808
rect 8904 19796 8910 19848
rect 8938 19796 8944 19848
rect 8996 19796 9002 19848
rect 10042 19796 10048 19848
rect 10100 19796 10106 19848
rect 10796 19845 10824 19876
rect 10597 19839 10655 19845
rect 10597 19805 10609 19839
rect 10643 19805 10655 19839
rect 10597 19799 10655 19805
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19805 10839 19839
rect 10781 19799 10839 19805
rect 11011 19839 11069 19845
rect 11011 19805 11023 19839
rect 11057 19836 11069 19839
rect 11057 19808 11376 19836
rect 11057 19805 11069 19808
rect 11011 19799 11069 19805
rect 6546 19728 6552 19780
rect 6604 19728 6610 19780
rect 7282 19728 7288 19780
rect 7340 19728 7346 19780
rect 7377 19771 7435 19777
rect 7377 19737 7389 19771
rect 7423 19737 7435 19771
rect 10410 19768 10416 19780
rect 7377 19731 7435 19737
rect 7668 19740 10416 19768
rect 7392 19700 7420 19731
rect 7668 19709 7696 19740
rect 10410 19728 10416 19740
rect 10468 19728 10474 19780
rect 3651 19672 7420 19700
rect 7653 19703 7711 19709
rect 3651 19669 3663 19672
rect 3605 19663 3663 19669
rect 7653 19669 7665 19703
rect 7699 19669 7711 19703
rect 7653 19663 7711 19669
rect 9582 19660 9588 19712
rect 9640 19660 9646 19712
rect 10134 19660 10140 19712
rect 10192 19660 10198 19712
rect 10612 19700 10640 19799
rect 10870 19728 10876 19780
rect 10928 19728 10934 19780
rect 11054 19700 11060 19712
rect 10612 19672 11060 19700
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 11146 19660 11152 19712
rect 11204 19660 11210 19712
rect 11348 19700 11376 19808
rect 12066 19796 12072 19848
rect 12124 19796 12130 19848
rect 12268 19845 12296 19944
rect 12434 19932 12440 19944
rect 12492 19932 12498 19984
rect 27264 19944 28028 19972
rect 27264 19848 27292 19944
rect 28000 19904 28028 19944
rect 27356 19876 27660 19904
rect 28000 19876 28120 19904
rect 27356 19848 27384 19876
rect 12253 19839 12311 19845
rect 12253 19805 12265 19839
rect 12299 19805 12311 19839
rect 12253 19799 12311 19805
rect 12342 19796 12348 19848
rect 12400 19796 12406 19848
rect 12526 19845 12532 19848
rect 12483 19839 12532 19845
rect 12483 19805 12495 19839
rect 12529 19805 12532 19839
rect 12483 19799 12532 19805
rect 12526 19796 12532 19799
rect 12584 19796 12590 19848
rect 12986 19796 12992 19848
rect 13044 19796 13050 19848
rect 13170 19796 13176 19848
rect 13228 19836 13234 19848
rect 13998 19836 14004 19848
rect 13228 19808 14004 19836
rect 13228 19796 13234 19808
rect 13998 19796 14004 19808
rect 14056 19836 14062 19848
rect 14734 19836 14740 19848
rect 14056 19808 14740 19836
rect 14056 19796 14062 19808
rect 14734 19796 14740 19808
rect 14792 19796 14798 19848
rect 15933 19839 15991 19845
rect 15933 19836 15945 19839
rect 14936 19808 15945 19836
rect 14936 19780 14964 19808
rect 15933 19805 15945 19808
rect 15979 19836 15991 19839
rect 17954 19836 17960 19848
rect 15979 19808 17960 19836
rect 15979 19805 15991 19808
rect 15933 19799 15991 19805
rect 17954 19796 17960 19808
rect 18012 19796 18018 19848
rect 27246 19796 27252 19848
rect 27304 19796 27310 19848
rect 27338 19796 27344 19848
rect 27396 19796 27402 19848
rect 27522 19846 27528 19848
rect 27448 19818 27528 19846
rect 14918 19728 14924 19780
rect 14976 19728 14982 19780
rect 15749 19771 15807 19777
rect 15749 19737 15761 19771
rect 15795 19768 15807 19771
rect 15838 19768 15844 19780
rect 15795 19740 15844 19768
rect 15795 19737 15807 19740
rect 15749 19731 15807 19737
rect 15838 19728 15844 19740
rect 15896 19728 15902 19780
rect 16850 19728 16856 19780
rect 16908 19768 16914 19780
rect 23382 19768 23388 19780
rect 16908 19740 19564 19768
rect 16908 19728 16914 19740
rect 19536 19712 19564 19740
rect 19628 19740 23388 19768
rect 19628 19712 19656 19740
rect 23382 19728 23388 19740
rect 23440 19728 23446 19780
rect 27448 19768 27476 19818
rect 27522 19796 27528 19818
rect 27580 19796 27586 19848
rect 27632 19845 27660 19876
rect 27617 19839 27675 19845
rect 27617 19805 27629 19839
rect 27663 19805 27675 19839
rect 27617 19799 27675 19805
rect 27801 19839 27859 19845
rect 27801 19805 27813 19839
rect 27847 19836 27859 19839
rect 27982 19836 27988 19848
rect 27847 19808 27988 19836
rect 27847 19805 27859 19808
rect 27801 19799 27859 19805
rect 27982 19796 27988 19808
rect 28040 19796 28046 19848
rect 28092 19845 28120 19876
rect 28077 19839 28135 19845
rect 28077 19805 28089 19839
rect 28123 19805 28135 19839
rect 28077 19799 28135 19805
rect 28166 19796 28172 19848
rect 28224 19836 28230 19848
rect 28353 19839 28411 19845
rect 28353 19836 28365 19839
rect 28224 19808 28365 19836
rect 28224 19796 28230 19808
rect 28353 19805 28365 19808
rect 28399 19805 28411 19839
rect 28353 19799 28411 19805
rect 28261 19771 28319 19777
rect 28261 19768 28273 19771
rect 27448 19740 28273 19768
rect 28261 19737 28273 19740
rect 28307 19737 28319 19771
rect 28261 19731 28319 19737
rect 12250 19700 12256 19712
rect 11348 19672 12256 19700
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 12894 19660 12900 19712
rect 12952 19700 12958 19712
rect 13541 19703 13599 19709
rect 13541 19700 13553 19703
rect 12952 19672 13553 19700
rect 12952 19660 12958 19672
rect 13541 19669 13553 19672
rect 13587 19669 13599 19703
rect 13541 19663 13599 19669
rect 14642 19660 14648 19712
rect 14700 19700 14706 19712
rect 17586 19700 17592 19712
rect 14700 19672 17592 19700
rect 14700 19660 14706 19672
rect 17586 19660 17592 19672
rect 17644 19700 17650 19712
rect 19334 19700 19340 19712
rect 17644 19672 19340 19700
rect 17644 19660 17650 19672
rect 19334 19660 19340 19672
rect 19392 19660 19398 19712
rect 19518 19660 19524 19712
rect 19576 19660 19582 19712
rect 19610 19660 19616 19712
rect 19668 19660 19674 19712
rect 19702 19660 19708 19712
rect 19760 19700 19766 19712
rect 26970 19700 26976 19712
rect 19760 19672 26976 19700
rect 19760 19660 19766 19672
rect 26970 19660 26976 19672
rect 27028 19660 27034 19712
rect 27062 19660 27068 19712
rect 27120 19660 27126 19712
rect 27433 19703 27491 19709
rect 27433 19669 27445 19703
rect 27479 19700 27491 19703
rect 27614 19700 27620 19712
rect 27479 19672 27620 19700
rect 27479 19669 27491 19672
rect 27433 19663 27491 19669
rect 27614 19660 27620 19672
rect 27672 19660 27678 19712
rect 27893 19703 27951 19709
rect 27893 19669 27905 19703
rect 27939 19700 27951 19703
rect 28718 19700 28724 19712
rect 27939 19672 28724 19700
rect 27939 19669 27951 19672
rect 27893 19663 27951 19669
rect 28718 19660 28724 19672
rect 28776 19660 28782 19712
rect 1104 19610 29595 19632
rect 1104 19558 8032 19610
rect 8084 19558 8096 19610
rect 8148 19558 8160 19610
rect 8212 19558 8224 19610
rect 8276 19558 8288 19610
rect 8340 19558 15115 19610
rect 15167 19558 15179 19610
rect 15231 19558 15243 19610
rect 15295 19558 15307 19610
rect 15359 19558 15371 19610
rect 15423 19558 22198 19610
rect 22250 19558 22262 19610
rect 22314 19558 22326 19610
rect 22378 19558 22390 19610
rect 22442 19558 22454 19610
rect 22506 19558 29281 19610
rect 29333 19558 29345 19610
rect 29397 19558 29409 19610
rect 29461 19558 29473 19610
rect 29525 19558 29537 19610
rect 29589 19558 29595 19610
rect 1104 19536 29595 19558
rect 1578 19456 1584 19508
rect 1636 19456 1642 19508
rect 9582 19496 9588 19508
rect 7300 19468 9588 19496
rect 1486 19320 1492 19372
rect 1544 19320 1550 19372
rect 6546 19320 6552 19372
rect 6604 19360 6610 19372
rect 7006 19360 7012 19372
rect 6604 19332 7012 19360
rect 6604 19320 6610 19332
rect 7006 19320 7012 19332
rect 7064 19320 7070 19372
rect 7300 19369 7328 19468
rect 9582 19456 9588 19468
rect 9640 19456 9646 19508
rect 11054 19456 11060 19508
rect 11112 19496 11118 19508
rect 12161 19499 12219 19505
rect 12161 19496 12173 19499
rect 11112 19468 12173 19496
rect 11112 19456 11118 19468
rect 12161 19465 12173 19468
rect 12207 19465 12219 19499
rect 12161 19459 12219 19465
rect 12250 19456 12256 19508
rect 12308 19496 12314 19508
rect 12526 19496 12532 19508
rect 12308 19468 12532 19496
rect 12308 19456 12314 19468
rect 12526 19456 12532 19468
rect 12584 19456 12590 19508
rect 12728 19468 13124 19496
rect 7561 19431 7619 19437
rect 7561 19397 7573 19431
rect 7607 19428 7619 19431
rect 7742 19428 7748 19440
rect 7607 19400 7748 19428
rect 7607 19397 7619 19400
rect 7561 19391 7619 19397
rect 7742 19388 7748 19400
rect 7800 19388 7806 19440
rect 8205 19431 8263 19437
rect 8205 19397 8217 19431
rect 8251 19428 8263 19431
rect 8478 19428 8484 19440
rect 8251 19400 8484 19428
rect 8251 19397 8263 19400
rect 8205 19391 8263 19397
rect 8478 19388 8484 19400
rect 8536 19388 8542 19440
rect 9766 19428 9772 19440
rect 9430 19400 9772 19428
rect 9766 19388 9772 19400
rect 9824 19388 9830 19440
rect 10870 19388 10876 19440
rect 10928 19428 10934 19440
rect 12618 19428 12624 19440
rect 10928 19400 12624 19428
rect 10928 19388 10934 19400
rect 12618 19388 12624 19400
rect 12676 19428 12682 19440
rect 12728 19428 12756 19468
rect 12676 19400 12756 19428
rect 12676 19388 12682 19400
rect 7285 19363 7343 19369
rect 7285 19329 7297 19363
rect 7331 19329 7343 19363
rect 7285 19323 7343 19329
rect 7469 19363 7527 19369
rect 7469 19329 7481 19363
rect 7515 19329 7527 19363
rect 7469 19323 7527 19329
rect 7024 19292 7052 19320
rect 7484 19292 7512 19323
rect 7650 19320 7656 19372
rect 7708 19320 7714 19372
rect 7926 19320 7932 19372
rect 7984 19320 7990 19372
rect 9858 19320 9864 19372
rect 9916 19360 9922 19372
rect 12805 19363 12863 19369
rect 9916 19332 12756 19360
rect 9916 19320 9922 19332
rect 7834 19292 7840 19304
rect 7024 19264 7840 19292
rect 7834 19252 7840 19264
rect 7892 19252 7898 19304
rect 8846 19252 8852 19304
rect 8904 19292 8910 19304
rect 9214 19292 9220 19304
rect 8904 19264 9220 19292
rect 8904 19252 8910 19264
rect 9214 19252 9220 19264
rect 9272 19292 9278 19304
rect 9677 19295 9735 19301
rect 9677 19292 9689 19295
rect 9272 19264 9689 19292
rect 9272 19252 9278 19264
rect 9677 19261 9689 19264
rect 9723 19261 9735 19295
rect 9677 19255 9735 19261
rect 11609 19295 11667 19301
rect 11609 19261 11621 19295
rect 11655 19292 11667 19295
rect 12158 19292 12164 19304
rect 11655 19264 12164 19292
rect 11655 19261 11667 19264
rect 11609 19255 11667 19261
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 12728 19292 12756 19332
rect 12805 19329 12817 19363
rect 12851 19360 12863 19363
rect 12894 19360 12900 19372
rect 12851 19332 12900 19360
rect 12851 19329 12863 19332
rect 12805 19323 12863 19329
rect 12894 19320 12900 19332
rect 12952 19320 12958 19372
rect 13096 19369 13124 19468
rect 13262 19456 13268 19508
rect 13320 19496 13326 19508
rect 13357 19499 13415 19505
rect 13357 19496 13369 19499
rect 13320 19468 13369 19496
rect 13320 19456 13326 19468
rect 13357 19465 13369 19468
rect 13403 19465 13415 19499
rect 13357 19459 13415 19465
rect 14550 19456 14556 19508
rect 14608 19456 14614 19508
rect 15194 19456 15200 19508
rect 15252 19496 15258 19508
rect 16114 19496 16120 19508
rect 15252 19468 16120 19496
rect 15252 19456 15258 19468
rect 16114 19456 16120 19468
rect 16172 19456 16178 19508
rect 16850 19456 16856 19508
rect 16908 19456 16914 19508
rect 17218 19456 17224 19508
rect 17276 19456 17282 19508
rect 17954 19456 17960 19508
rect 18012 19496 18018 19508
rect 18969 19499 19027 19505
rect 18969 19496 18981 19499
rect 18012 19468 18981 19496
rect 18012 19456 18018 19468
rect 18969 19465 18981 19468
rect 19015 19465 19027 19499
rect 18969 19459 19027 19465
rect 19058 19456 19064 19508
rect 19116 19456 19122 19508
rect 19702 19496 19708 19508
rect 19168 19468 19708 19496
rect 12989 19363 13047 19369
rect 12989 19329 13001 19363
rect 13035 19329 13047 19363
rect 12989 19323 13047 19329
rect 13081 19363 13139 19369
rect 13081 19329 13093 19363
rect 13127 19329 13139 19363
rect 13081 19323 13139 19329
rect 13004 19292 13032 19323
rect 13170 19320 13176 19372
rect 13228 19320 13234 19372
rect 14568 19360 14596 19456
rect 16393 19431 16451 19437
rect 16393 19428 16405 19431
rect 14936 19400 16405 19428
rect 14936 19369 14964 19400
rect 16393 19397 16405 19400
rect 16439 19397 16451 19431
rect 16393 19391 16451 19397
rect 13280 19332 14596 19360
rect 14921 19363 14979 19369
rect 13280 19292 13308 19332
rect 14921 19329 14933 19363
rect 14967 19329 14979 19363
rect 14921 19323 14979 19329
rect 15102 19320 15108 19372
rect 15160 19320 15166 19372
rect 15197 19363 15255 19369
rect 15197 19329 15209 19363
rect 15243 19329 15255 19363
rect 15197 19323 15255 19329
rect 12728 19264 13308 19292
rect 15212 19292 15240 19323
rect 15286 19320 15292 19372
rect 15344 19320 15350 19372
rect 15562 19360 15568 19372
rect 15396 19332 15568 19360
rect 15396 19292 15424 19332
rect 15562 19320 15568 19332
rect 15620 19360 15626 19372
rect 16868 19369 16896 19456
rect 16945 19431 17003 19437
rect 16945 19397 16957 19431
rect 16991 19428 17003 19431
rect 19168 19428 19196 19468
rect 19702 19456 19708 19468
rect 19760 19456 19766 19508
rect 19886 19456 19892 19508
rect 19944 19456 19950 19508
rect 20530 19456 20536 19508
rect 20588 19456 20594 19508
rect 28074 19456 28080 19508
rect 28132 19456 28138 19508
rect 16991 19400 19196 19428
rect 19245 19431 19303 19437
rect 16991 19397 17003 19400
rect 16945 19391 17003 19397
rect 19245 19397 19257 19431
rect 19291 19428 19303 19431
rect 19426 19428 19432 19440
rect 19291 19400 19432 19428
rect 19291 19397 19303 19400
rect 19245 19391 19303 19397
rect 19426 19388 19432 19400
rect 19484 19388 19490 19440
rect 19610 19388 19616 19440
rect 19668 19388 19674 19440
rect 20257 19431 20315 19437
rect 20257 19397 20269 19431
rect 20303 19428 20315 19431
rect 22554 19428 22560 19440
rect 20303 19400 22560 19428
rect 20303 19397 20315 19400
rect 20257 19391 20315 19397
rect 22554 19388 22560 19400
rect 22612 19388 22618 19440
rect 28092 19428 28120 19456
rect 27540 19400 28120 19428
rect 16669 19363 16727 19369
rect 16669 19360 16681 19363
rect 15620 19332 16681 19360
rect 15620 19320 15626 19332
rect 16669 19329 16681 19332
rect 16715 19329 16727 19363
rect 16669 19323 16727 19329
rect 16853 19363 16911 19369
rect 16853 19329 16865 19363
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 17037 19363 17095 19369
rect 17037 19329 17049 19363
rect 17083 19360 17095 19363
rect 18877 19363 18935 19369
rect 17083 19332 18828 19360
rect 17083 19329 17095 19332
rect 17037 19323 17095 19329
rect 15212 19264 15424 19292
rect 15841 19295 15899 19301
rect 15841 19261 15853 19295
rect 15887 19292 15899 19295
rect 15930 19292 15936 19304
rect 15887 19264 15936 19292
rect 15887 19261 15899 19264
rect 15841 19255 15899 19261
rect 15930 19252 15936 19264
rect 15988 19252 15994 19304
rect 6454 19184 6460 19236
rect 6512 19224 6518 19236
rect 6512 19196 7972 19224
rect 6512 19184 6518 19196
rect 7834 19116 7840 19168
rect 7892 19116 7898 19168
rect 7944 19156 7972 19196
rect 9582 19184 9588 19236
rect 9640 19224 9646 19236
rect 17954 19224 17960 19236
rect 9640 19196 17960 19224
rect 9640 19184 9646 19196
rect 17954 19184 17960 19196
rect 18012 19184 18018 19236
rect 18693 19227 18751 19233
rect 18693 19193 18705 19227
rect 18739 19193 18751 19227
rect 18800 19224 18828 19332
rect 18877 19329 18889 19363
rect 18923 19360 18935 19363
rect 18923 19332 19288 19360
rect 18923 19329 18935 19332
rect 18877 19323 18935 19329
rect 19260 19292 19288 19332
rect 19334 19320 19340 19372
rect 19392 19320 19398 19372
rect 19518 19320 19524 19372
rect 19576 19320 19582 19372
rect 19705 19363 19763 19369
rect 19705 19329 19717 19363
rect 19751 19360 19763 19363
rect 19981 19363 20039 19369
rect 19751 19332 19932 19360
rect 19751 19329 19763 19332
rect 19705 19323 19763 19329
rect 19610 19292 19616 19304
rect 19260 19264 19616 19292
rect 19610 19252 19616 19264
rect 19668 19252 19674 19304
rect 19904 19292 19932 19332
rect 19981 19329 19993 19363
rect 20027 19360 20039 19363
rect 20070 19360 20076 19372
rect 20027 19332 20076 19360
rect 20027 19329 20039 19332
rect 19981 19323 20039 19329
rect 20070 19320 20076 19332
rect 20128 19320 20134 19372
rect 20162 19320 20168 19372
rect 20220 19320 20226 19372
rect 20349 19363 20407 19369
rect 20349 19329 20361 19363
rect 20395 19329 20407 19363
rect 20349 19323 20407 19329
rect 20364 19292 20392 19323
rect 27430 19320 27436 19372
rect 27488 19320 27494 19372
rect 27540 19369 27568 19400
rect 27525 19363 27583 19369
rect 27525 19329 27537 19363
rect 27571 19329 27583 19363
rect 27525 19323 27583 19329
rect 27617 19363 27675 19369
rect 27617 19329 27629 19363
rect 27663 19329 27675 19363
rect 27617 19323 27675 19329
rect 19904 19264 20392 19292
rect 27448 19292 27476 19320
rect 27632 19292 27660 19323
rect 27448 19264 27660 19292
rect 19794 19224 19800 19236
rect 18800 19196 19800 19224
rect 18693 19187 18751 19193
rect 12618 19156 12624 19168
rect 7944 19128 12624 19156
rect 12618 19116 12624 19128
rect 12676 19116 12682 19168
rect 12710 19116 12716 19168
rect 12768 19156 12774 19168
rect 12894 19156 12900 19168
rect 12768 19128 12900 19156
rect 12768 19116 12774 19128
rect 12894 19116 12900 19128
rect 12952 19156 12958 19168
rect 13722 19156 13728 19168
rect 12952 19128 13728 19156
rect 12952 19116 12958 19128
rect 13722 19116 13728 19128
rect 13780 19116 13786 19168
rect 13814 19116 13820 19168
rect 13872 19156 13878 19168
rect 15010 19156 15016 19168
rect 13872 19128 15016 19156
rect 13872 19116 13878 19128
rect 15010 19116 15016 19128
rect 15068 19116 15074 19168
rect 15470 19116 15476 19168
rect 15528 19116 15534 19168
rect 18708 19156 18736 19187
rect 19794 19184 19800 19196
rect 19852 19224 19858 19236
rect 19904 19224 19932 19264
rect 27798 19252 27804 19304
rect 27856 19252 27862 19304
rect 19852 19196 19932 19224
rect 19852 19184 19858 19196
rect 21266 19156 21272 19168
rect 18708 19128 21272 19156
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 1104 19066 29440 19088
rect 1104 19014 4491 19066
rect 4543 19014 4555 19066
rect 4607 19014 4619 19066
rect 4671 19014 4683 19066
rect 4735 19014 4747 19066
rect 4799 19014 11574 19066
rect 11626 19014 11638 19066
rect 11690 19014 11702 19066
rect 11754 19014 11766 19066
rect 11818 19014 11830 19066
rect 11882 19014 18657 19066
rect 18709 19014 18721 19066
rect 18773 19014 18785 19066
rect 18837 19014 18849 19066
rect 18901 19014 18913 19066
rect 18965 19014 25740 19066
rect 25792 19014 25804 19066
rect 25856 19014 25868 19066
rect 25920 19014 25932 19066
rect 25984 19014 25996 19066
rect 26048 19014 29440 19066
rect 1104 18992 29440 19014
rect 8757 18955 8815 18961
rect 8757 18921 8769 18955
rect 8803 18952 8815 18955
rect 8938 18952 8944 18964
rect 8803 18924 8944 18952
rect 8803 18921 8815 18924
rect 8757 18915 8815 18921
rect 8938 18912 8944 18924
rect 8996 18912 9002 18964
rect 9582 18912 9588 18964
rect 9640 18912 9646 18964
rect 11885 18955 11943 18961
rect 11885 18921 11897 18955
rect 11931 18952 11943 18955
rect 12158 18952 12164 18964
rect 11931 18924 12164 18952
rect 11931 18921 11943 18924
rect 11885 18915 11943 18921
rect 12158 18912 12164 18924
rect 12216 18912 12222 18964
rect 12802 18952 12808 18964
rect 12268 18924 12808 18952
rect 6362 18776 6368 18828
rect 6420 18816 6426 18828
rect 7009 18819 7067 18825
rect 7009 18816 7021 18819
rect 6420 18788 7021 18816
rect 6420 18776 6426 18788
rect 7009 18785 7021 18788
rect 7055 18785 7067 18819
rect 7009 18779 7067 18785
rect 7285 18819 7343 18825
rect 7285 18785 7297 18819
rect 7331 18816 7343 18819
rect 7834 18816 7840 18828
rect 7331 18788 7840 18816
rect 7331 18785 7343 18788
rect 7285 18779 7343 18785
rect 7834 18776 7840 18788
rect 7892 18776 7898 18828
rect 8956 18816 8984 18912
rect 8956 18788 9076 18816
rect 3510 18708 3516 18760
rect 3568 18748 3574 18760
rect 4065 18751 4123 18757
rect 4065 18748 4077 18751
rect 3568 18720 4077 18748
rect 3568 18708 3574 18720
rect 4065 18717 4077 18720
rect 4111 18748 4123 18751
rect 6181 18751 6239 18757
rect 4111 18720 5304 18748
rect 4111 18717 4123 18720
rect 4065 18711 4123 18717
rect 5276 18624 5304 18720
rect 6181 18717 6193 18751
rect 6227 18748 6239 18751
rect 6227 18720 6316 18748
rect 6227 18717 6239 18720
rect 6181 18711 6239 18717
rect 6288 18692 6316 18720
rect 6454 18708 6460 18760
rect 6512 18708 6518 18760
rect 6549 18751 6607 18757
rect 6549 18717 6561 18751
rect 6595 18748 6607 18751
rect 6914 18748 6920 18760
rect 6595 18720 6920 18748
rect 6595 18717 6607 18720
rect 6549 18711 6607 18717
rect 6914 18708 6920 18720
rect 6972 18708 6978 18760
rect 8570 18708 8576 18760
rect 8628 18748 8634 18760
rect 9048 18757 9076 18788
rect 9214 18776 9220 18828
rect 9272 18776 9278 18828
rect 9950 18776 9956 18828
rect 10008 18816 10014 18828
rect 10137 18819 10195 18825
rect 10137 18816 10149 18819
rect 10008 18788 10149 18816
rect 10008 18776 10014 18788
rect 10137 18785 10149 18788
rect 10183 18785 10195 18819
rect 10137 18779 10195 18785
rect 10413 18819 10471 18825
rect 10413 18785 10425 18819
rect 10459 18816 10471 18819
rect 11146 18816 11152 18828
rect 10459 18788 11152 18816
rect 10459 18785 10471 18788
rect 10413 18779 10471 18785
rect 11146 18776 11152 18788
rect 11204 18776 11210 18828
rect 12268 18816 12296 18924
rect 12802 18912 12808 18924
rect 12860 18952 12866 18964
rect 13170 18952 13176 18964
rect 12860 18924 13176 18952
rect 12860 18912 12866 18924
rect 13170 18912 13176 18924
rect 13228 18912 13234 18964
rect 13814 18912 13820 18964
rect 13872 18912 13878 18964
rect 13906 18912 13912 18964
rect 13964 18952 13970 18964
rect 13964 18924 15700 18952
rect 13964 18912 13970 18924
rect 12618 18844 12624 18896
rect 12676 18884 12682 18896
rect 13832 18884 13860 18912
rect 12676 18856 13860 18884
rect 12676 18844 12682 18856
rect 15470 18844 15476 18896
rect 15528 18844 15534 18896
rect 15562 18844 15568 18896
rect 15620 18844 15626 18896
rect 15672 18884 15700 18924
rect 15930 18912 15936 18964
rect 15988 18912 15994 18964
rect 19426 18912 19432 18964
rect 19484 18952 19490 18964
rect 19797 18955 19855 18961
rect 19797 18952 19809 18955
rect 19484 18924 19809 18952
rect 19484 18912 19490 18924
rect 19797 18921 19809 18924
rect 19843 18921 19855 18955
rect 19797 18915 19855 18921
rect 19886 18912 19892 18964
rect 19944 18952 19950 18964
rect 20257 18955 20315 18961
rect 20257 18952 20269 18955
rect 19944 18924 20269 18952
rect 19944 18912 19950 18924
rect 20257 18921 20269 18924
rect 20303 18921 20315 18955
rect 20257 18915 20315 18921
rect 28997 18955 29055 18961
rect 28997 18921 29009 18955
rect 29043 18952 29055 18955
rect 29043 18924 29500 18952
rect 29043 18921 29055 18924
rect 28997 18915 29055 18921
rect 29472 18896 29500 18924
rect 17678 18884 17684 18896
rect 15672 18856 17684 18884
rect 17678 18844 17684 18856
rect 17736 18844 17742 18896
rect 19150 18844 19156 18896
rect 19208 18884 19214 18896
rect 19208 18856 20116 18884
rect 19208 18844 19214 18856
rect 11532 18788 12296 18816
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8628 18720 8953 18748
rect 8628 18708 8634 18720
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 9034 18751 9092 18757
rect 9034 18717 9046 18751
rect 9080 18717 9092 18751
rect 9232 18748 9260 18776
rect 9309 18751 9367 18757
rect 9309 18748 9321 18751
rect 9232 18720 9321 18748
rect 9034 18711 9092 18717
rect 9309 18717 9321 18720
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 9398 18708 9404 18760
rect 9456 18757 9462 18760
rect 9456 18748 9464 18757
rect 9456 18720 9501 18748
rect 9456 18711 9464 18720
rect 9456 18708 9462 18711
rect 6270 18640 6276 18692
rect 6328 18640 6334 18692
rect 6365 18683 6423 18689
rect 6365 18649 6377 18683
rect 6411 18680 6423 18683
rect 7006 18680 7012 18692
rect 6411 18652 7012 18680
rect 6411 18649 6423 18652
rect 6365 18643 6423 18649
rect 7006 18640 7012 18652
rect 7064 18640 7070 18692
rect 7282 18640 7288 18692
rect 7340 18640 7346 18692
rect 7742 18640 7748 18692
rect 7800 18640 7806 18692
rect 9217 18683 9275 18689
rect 9217 18649 9229 18683
rect 9263 18649 9275 18683
rect 9217 18643 9275 18649
rect 3970 18572 3976 18624
rect 4028 18612 4034 18624
rect 4709 18615 4767 18621
rect 4709 18612 4721 18615
rect 4028 18584 4721 18612
rect 4028 18572 4034 18584
rect 4709 18581 4721 18584
rect 4755 18581 4767 18615
rect 4709 18575 4767 18581
rect 5258 18572 5264 18624
rect 5316 18572 5322 18624
rect 5810 18572 5816 18624
rect 5868 18612 5874 18624
rect 6733 18615 6791 18621
rect 6733 18612 6745 18615
rect 5868 18584 6745 18612
rect 5868 18572 5874 18584
rect 6733 18581 6745 18584
rect 6779 18581 6791 18615
rect 7300 18612 7328 18640
rect 9232 18612 9260 18643
rect 7300 18584 9260 18612
rect 6733 18575 6791 18581
rect 9306 18572 9312 18624
rect 9364 18612 9370 18624
rect 10686 18612 10692 18624
rect 9364 18584 10692 18612
rect 9364 18572 9370 18584
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 11054 18572 11060 18624
rect 11112 18612 11118 18624
rect 11532 18612 11560 18788
rect 12526 18776 12532 18828
rect 12584 18776 12590 18828
rect 14461 18819 14519 18825
rect 14461 18785 14473 18819
rect 14507 18816 14519 18819
rect 15488 18816 15516 18844
rect 14507 18788 15516 18816
rect 15580 18816 15608 18844
rect 19061 18819 19119 18825
rect 19061 18816 19073 18819
rect 15580 18788 16896 18816
rect 14507 18785 14519 18788
rect 14461 18779 14519 18785
rect 12253 18751 12311 18757
rect 12253 18717 12265 18751
rect 12299 18717 12311 18751
rect 12544 18748 12572 18776
rect 16500 18760 16528 18788
rect 12621 18751 12679 18757
rect 12621 18748 12633 18751
rect 12544 18720 12633 18748
rect 12253 18711 12311 18717
rect 12621 18717 12633 18720
rect 12667 18717 12679 18751
rect 12621 18711 12679 18717
rect 11112 18584 11560 18612
rect 12268 18612 12296 18711
rect 12710 18708 12716 18760
rect 12768 18708 12774 18760
rect 14185 18751 14243 18757
rect 14185 18717 14197 18751
rect 14231 18717 14243 18751
rect 14185 18711 14243 18717
rect 16301 18751 16359 18757
rect 16301 18717 16313 18751
rect 16347 18748 16359 18751
rect 16482 18748 16488 18760
rect 16347 18720 16488 18748
rect 16347 18717 16359 18720
rect 16301 18711 16359 18717
rect 12342 18640 12348 18692
rect 12400 18680 12406 18692
rect 12437 18683 12495 18689
rect 12437 18680 12449 18683
rect 12400 18652 12449 18680
rect 12400 18640 12406 18652
rect 12437 18649 12449 18652
rect 12483 18649 12495 18683
rect 12437 18643 12495 18649
rect 12529 18683 12587 18689
rect 12529 18649 12541 18683
rect 12575 18680 12587 18683
rect 12728 18680 12756 18708
rect 14200 18680 14228 18711
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 16577 18751 16635 18757
rect 16577 18717 16589 18751
rect 16623 18748 16635 18751
rect 16758 18748 16764 18760
rect 16623 18720 16764 18748
rect 16623 18717 16635 18720
rect 16577 18711 16635 18717
rect 14366 18680 14372 18692
rect 12575 18652 14136 18680
rect 14200 18652 14372 18680
rect 12575 18649 12587 18652
rect 12529 18643 12587 18649
rect 12710 18612 12716 18624
rect 12268 18584 12716 18612
rect 11112 18572 11118 18584
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 12802 18572 12808 18624
rect 12860 18572 12866 18624
rect 14108 18612 14136 18652
rect 14366 18640 14372 18652
rect 14424 18640 14430 18692
rect 14550 18640 14556 18692
rect 14608 18640 14614 18692
rect 15470 18640 15476 18692
rect 15528 18640 15534 18692
rect 16592 18680 16620 18711
rect 16758 18708 16764 18720
rect 16816 18708 16822 18760
rect 16040 18652 16620 18680
rect 16868 18680 16896 18788
rect 17420 18788 19073 18816
rect 17420 18757 17448 18788
rect 19061 18785 19073 18788
rect 19107 18785 19119 18819
rect 19061 18779 19119 18785
rect 19168 18788 19932 18816
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18717 17463 18751
rect 17773 18751 17831 18757
rect 17773 18748 17785 18751
rect 17405 18711 17463 18717
rect 17512 18720 17785 18748
rect 17512 18680 17540 18720
rect 17773 18717 17785 18720
rect 17819 18717 17831 18751
rect 17773 18711 17831 18717
rect 18509 18751 18567 18757
rect 18509 18717 18521 18751
rect 18555 18748 18567 18751
rect 18782 18748 18788 18760
rect 18555 18720 18788 18748
rect 18555 18717 18567 18720
rect 18509 18711 18567 18717
rect 18782 18708 18788 18720
rect 18840 18748 18846 18760
rect 19168 18748 19196 18788
rect 18840 18720 19196 18748
rect 19245 18751 19303 18757
rect 18840 18708 18846 18720
rect 19245 18717 19257 18751
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18748 19671 18751
rect 19794 18748 19800 18760
rect 19659 18720 19800 18748
rect 19659 18717 19671 18720
rect 19613 18711 19671 18717
rect 16868 18652 17540 18680
rect 17589 18683 17647 18689
rect 14568 18612 14596 18640
rect 14108 18584 14596 18612
rect 14734 18572 14740 18624
rect 14792 18612 14798 18624
rect 16040 18612 16068 18652
rect 17589 18649 17601 18683
rect 17635 18649 17647 18683
rect 17589 18643 17647 18649
rect 14792 18584 16068 18612
rect 14792 18572 14798 18584
rect 16114 18572 16120 18624
rect 16172 18612 16178 18624
rect 17494 18612 17500 18624
rect 16172 18584 17500 18612
rect 16172 18572 16178 18584
rect 17494 18572 17500 18584
rect 17552 18612 17558 18624
rect 17604 18612 17632 18643
rect 17678 18640 17684 18692
rect 17736 18680 17742 18692
rect 19260 18680 19288 18711
rect 19794 18708 19800 18720
rect 19852 18708 19858 18760
rect 19904 18757 19932 18788
rect 20088 18757 20116 18856
rect 29454 18844 29460 18896
rect 29512 18844 29518 18896
rect 19889 18751 19947 18757
rect 19889 18717 19901 18751
rect 19935 18717 19947 18751
rect 19889 18711 19947 18717
rect 20073 18751 20131 18757
rect 20073 18717 20085 18751
rect 20119 18717 20131 18751
rect 20073 18711 20131 18717
rect 27706 18708 27712 18760
rect 27764 18748 27770 18760
rect 28813 18751 28871 18757
rect 28813 18748 28825 18751
rect 27764 18720 28825 18748
rect 27764 18708 27770 18720
rect 28813 18717 28825 18720
rect 28859 18717 28871 18751
rect 28813 18711 28871 18717
rect 17736 18652 19288 18680
rect 17736 18640 17742 18652
rect 19426 18640 19432 18692
rect 19484 18640 19490 18692
rect 19521 18683 19579 18689
rect 19521 18649 19533 18683
rect 19567 18680 19579 18683
rect 23290 18680 23296 18692
rect 19567 18652 23296 18680
rect 19567 18649 19579 18652
rect 19521 18643 19579 18649
rect 23290 18640 23296 18652
rect 23348 18640 23354 18692
rect 17552 18584 17632 18612
rect 17552 18572 17558 18584
rect 17954 18572 17960 18624
rect 18012 18572 18018 18624
rect 23934 18572 23940 18624
rect 23992 18612 23998 18624
rect 24486 18612 24492 18624
rect 23992 18584 24492 18612
rect 23992 18572 23998 18584
rect 24486 18572 24492 18584
rect 24544 18572 24550 18624
rect 1104 18522 29595 18544
rect 1104 18470 8032 18522
rect 8084 18470 8096 18522
rect 8148 18470 8160 18522
rect 8212 18470 8224 18522
rect 8276 18470 8288 18522
rect 8340 18470 15115 18522
rect 15167 18470 15179 18522
rect 15231 18470 15243 18522
rect 15295 18470 15307 18522
rect 15359 18470 15371 18522
rect 15423 18470 22198 18522
rect 22250 18470 22262 18522
rect 22314 18470 22326 18522
rect 22378 18470 22390 18522
rect 22442 18470 22454 18522
rect 22506 18470 29281 18522
rect 29333 18470 29345 18522
rect 29397 18470 29409 18522
rect 29461 18470 29473 18522
rect 29525 18470 29537 18522
rect 29589 18470 29595 18522
rect 1104 18448 29595 18470
rect 1854 18368 1860 18420
rect 1912 18408 1918 18420
rect 3694 18408 3700 18420
rect 1912 18380 3700 18408
rect 1912 18368 1918 18380
rect 3694 18368 3700 18380
rect 3752 18368 3758 18420
rect 6270 18368 6276 18420
rect 6328 18408 6334 18420
rect 8205 18411 8263 18417
rect 8205 18408 8217 18411
rect 6328 18380 8217 18408
rect 6328 18368 6334 18380
rect 8205 18377 8217 18380
rect 8251 18377 8263 18411
rect 8205 18371 8263 18377
rect 9306 18368 9312 18420
rect 9364 18368 9370 18420
rect 9674 18368 9680 18420
rect 9732 18408 9738 18420
rect 11333 18411 11391 18417
rect 11333 18408 11345 18411
rect 9732 18380 11345 18408
rect 9732 18368 9738 18380
rect 11333 18377 11345 18380
rect 11379 18377 11391 18411
rect 12618 18408 12624 18420
rect 11333 18371 11391 18377
rect 12406 18380 12624 18408
rect 1872 18281 1900 18368
rect 5258 18300 5264 18352
rect 5316 18340 5322 18352
rect 5905 18343 5963 18349
rect 5905 18340 5917 18343
rect 5316 18312 5917 18340
rect 5316 18300 5322 18312
rect 5905 18309 5917 18312
rect 5951 18309 5963 18343
rect 5905 18303 5963 18309
rect 1857 18275 1915 18281
rect 1857 18241 1869 18275
rect 1903 18241 1915 18275
rect 1857 18235 1915 18241
rect 3234 18232 3240 18284
rect 3292 18232 3298 18284
rect 3694 18232 3700 18284
rect 3752 18232 3758 18284
rect 5629 18275 5687 18281
rect 5629 18272 5641 18275
rect 5106 18244 5304 18272
rect 5276 18216 5304 18244
rect 5460 18244 5641 18272
rect 2133 18207 2191 18213
rect 2133 18173 2145 18207
rect 2179 18204 2191 18207
rect 3418 18204 3424 18216
rect 2179 18176 3424 18204
rect 2179 18173 2191 18176
rect 2133 18167 2191 18173
rect 3418 18164 3424 18176
rect 3476 18164 3482 18216
rect 3510 18164 3516 18216
rect 3568 18204 3574 18216
rect 3605 18207 3663 18213
rect 3605 18204 3617 18207
rect 3568 18176 3617 18204
rect 3568 18164 3574 18176
rect 3605 18173 3617 18176
rect 3651 18173 3663 18207
rect 3605 18167 3663 18173
rect 3973 18207 4031 18213
rect 3973 18173 3985 18207
rect 4019 18204 4031 18207
rect 4019 18176 5120 18204
rect 4019 18173 4031 18176
rect 3973 18167 4031 18173
rect 5092 18148 5120 18176
rect 5258 18164 5264 18216
rect 5316 18164 5322 18216
rect 5074 18096 5080 18148
rect 5132 18096 5138 18148
rect 5166 18028 5172 18080
rect 5224 18068 5230 18080
rect 5460 18077 5488 18244
rect 5629 18241 5641 18244
rect 5675 18241 5687 18275
rect 5629 18235 5687 18241
rect 5718 18232 5724 18284
rect 5776 18272 5782 18284
rect 5813 18275 5871 18281
rect 5813 18272 5825 18275
rect 5776 18244 5825 18272
rect 5776 18232 5782 18244
rect 5813 18241 5825 18244
rect 5859 18241 5871 18275
rect 5813 18235 5871 18241
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18272 6055 18275
rect 6270 18272 6276 18284
rect 6043 18244 6276 18272
rect 6043 18241 6055 18244
rect 5997 18235 6055 18241
rect 5828 18204 5856 18235
rect 6270 18232 6276 18244
rect 6328 18272 6334 18284
rect 6730 18272 6736 18284
rect 6328 18244 6736 18272
rect 6328 18232 6334 18244
rect 6730 18232 6736 18244
rect 6788 18232 6794 18284
rect 6825 18275 6883 18281
rect 6825 18241 6837 18275
rect 6871 18241 6883 18275
rect 6825 18235 6883 18241
rect 6546 18204 6552 18216
rect 5828 18176 6552 18204
rect 6546 18164 6552 18176
rect 6604 18164 6610 18216
rect 6840 18204 6868 18235
rect 6914 18232 6920 18284
rect 6972 18272 6978 18284
rect 7193 18275 7251 18281
rect 7193 18272 7205 18275
rect 6972 18244 7205 18272
rect 6972 18232 6978 18244
rect 7193 18241 7205 18244
rect 7239 18272 7251 18275
rect 7650 18272 7656 18284
rect 7239 18244 7656 18272
rect 7239 18241 7251 18244
rect 7193 18235 7251 18241
rect 7650 18232 7656 18244
rect 7708 18272 7714 18284
rect 7834 18272 7840 18284
rect 7708 18244 7840 18272
rect 7708 18232 7714 18244
rect 7834 18232 7840 18244
rect 7892 18232 7898 18284
rect 6840 18176 6960 18204
rect 6932 18136 6960 18176
rect 7006 18164 7012 18216
rect 7064 18204 7070 18216
rect 7285 18207 7343 18213
rect 7285 18204 7297 18207
rect 7064 18176 7297 18204
rect 7064 18164 7070 18176
rect 7285 18173 7297 18176
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 7558 18164 7564 18216
rect 7616 18164 7622 18216
rect 7098 18136 7104 18148
rect 6932 18108 7104 18136
rect 7098 18096 7104 18108
rect 7156 18136 7162 18148
rect 9324 18136 9352 18368
rect 10321 18343 10379 18349
rect 10321 18340 10333 18343
rect 9416 18312 10333 18340
rect 9416 18281 9444 18312
rect 10321 18309 10333 18312
rect 10367 18340 10379 18343
rect 12406 18340 12434 18380
rect 12618 18368 12624 18380
rect 12676 18368 12682 18420
rect 12710 18368 12716 18420
rect 12768 18408 12774 18420
rect 14001 18411 14059 18417
rect 14001 18408 14013 18411
rect 12768 18380 14013 18408
rect 12768 18368 12774 18380
rect 14001 18377 14013 18380
rect 14047 18377 14059 18411
rect 14001 18371 14059 18377
rect 14366 18368 14372 18420
rect 14424 18408 14430 18420
rect 16574 18408 16580 18420
rect 14424 18380 16580 18408
rect 14424 18368 14430 18380
rect 10367 18312 12434 18340
rect 12989 18343 13047 18349
rect 10367 18309 10379 18312
rect 10321 18303 10379 18309
rect 12989 18309 13001 18343
rect 13035 18340 13047 18343
rect 13906 18340 13912 18352
rect 13035 18312 13912 18340
rect 13035 18309 13047 18312
rect 12989 18303 13047 18309
rect 13906 18300 13912 18312
rect 13964 18300 13970 18352
rect 9401 18275 9459 18281
rect 9401 18241 9413 18275
rect 9447 18241 9459 18275
rect 9401 18235 9459 18241
rect 9585 18275 9643 18281
rect 9585 18241 9597 18275
rect 9631 18241 9643 18275
rect 9585 18235 9643 18241
rect 9600 18204 9628 18235
rect 9674 18232 9680 18284
rect 9732 18232 9738 18284
rect 9766 18232 9772 18284
rect 9824 18232 9830 18284
rect 10045 18275 10103 18281
rect 10045 18241 10057 18275
rect 10091 18272 10103 18275
rect 10091 18244 10180 18272
rect 10091 18241 10103 18244
rect 10045 18235 10103 18241
rect 9600 18176 10088 18204
rect 7156 18108 9352 18136
rect 7156 18096 7162 18108
rect 9490 18096 9496 18148
rect 9548 18136 9554 18148
rect 9646 18136 9674 18176
rect 9548 18108 9674 18136
rect 9548 18096 9554 18108
rect 10060 18080 10088 18176
rect 10152 18136 10180 18244
rect 10226 18232 10232 18284
rect 10284 18232 10290 18284
rect 10413 18275 10471 18281
rect 10413 18272 10425 18275
rect 10336 18244 10425 18272
rect 10336 18216 10364 18244
rect 10413 18241 10425 18244
rect 10459 18241 10471 18275
rect 10413 18235 10471 18241
rect 12618 18232 12624 18284
rect 12676 18232 12682 18284
rect 12769 18275 12827 18281
rect 12769 18241 12781 18275
rect 12815 18272 12827 18275
rect 12815 18241 12848 18272
rect 12769 18235 12848 18241
rect 10318 18164 10324 18216
rect 10376 18164 10382 18216
rect 10781 18207 10839 18213
rect 10781 18173 10793 18207
rect 10827 18204 10839 18207
rect 11238 18204 11244 18216
rect 10827 18176 11244 18204
rect 10827 18173 10839 18176
rect 10781 18167 10839 18173
rect 11238 18164 11244 18176
rect 11296 18164 11302 18216
rect 11330 18164 11336 18216
rect 11388 18204 11394 18216
rect 11517 18207 11575 18213
rect 11517 18204 11529 18207
rect 11388 18176 11529 18204
rect 11388 18164 11394 18176
rect 11517 18173 11529 18176
rect 11563 18173 11575 18207
rect 12820 18204 12848 18235
rect 12894 18232 12900 18284
rect 12952 18232 12958 18284
rect 13127 18275 13185 18281
rect 13127 18241 13139 18275
rect 13173 18272 13185 18275
rect 13354 18272 13360 18284
rect 13173 18244 13360 18272
rect 13173 18241 13185 18244
rect 13127 18235 13185 18241
rect 13354 18232 13360 18244
rect 13412 18232 13418 18284
rect 14752 18281 14780 18380
rect 16574 18368 16580 18380
rect 16632 18408 16638 18420
rect 17954 18408 17960 18420
rect 16632 18380 17080 18408
rect 16632 18368 16638 18380
rect 15470 18300 15476 18352
rect 15528 18300 15534 18352
rect 17052 18281 17080 18380
rect 17328 18380 17960 18408
rect 17328 18349 17356 18380
rect 17954 18368 17960 18380
rect 18012 18368 18018 18420
rect 18138 18368 18144 18420
rect 18196 18408 18202 18420
rect 18196 18380 18644 18408
rect 18196 18368 18202 18380
rect 17313 18343 17371 18349
rect 17313 18309 17325 18343
rect 17359 18309 17371 18343
rect 17313 18303 17371 18309
rect 14737 18275 14795 18281
rect 14737 18241 14749 18275
rect 14783 18241 14795 18275
rect 14737 18235 14795 18241
rect 17037 18275 17095 18281
rect 17037 18241 17049 18275
rect 17083 18241 17095 18275
rect 18616 18272 18644 18380
rect 18782 18368 18788 18420
rect 18840 18368 18846 18420
rect 19978 18368 19984 18420
rect 20036 18408 20042 18420
rect 20993 18411 21051 18417
rect 20036 18380 20852 18408
rect 20036 18368 20042 18380
rect 20162 18340 20168 18352
rect 19536 18312 20168 18340
rect 19536 18284 19564 18312
rect 20162 18300 20168 18312
rect 20220 18340 20226 18352
rect 20220 18312 20668 18340
rect 20220 18300 20226 18312
rect 19058 18272 19064 18284
rect 17037 18235 17095 18241
rect 13449 18207 13507 18213
rect 13449 18204 13461 18207
rect 12820 18176 13461 18204
rect 11517 18167 11575 18173
rect 13449 18173 13461 18176
rect 13495 18204 13507 18207
rect 13814 18204 13820 18216
rect 13495 18176 13820 18204
rect 13495 18173 13507 18176
rect 13449 18167 13507 18173
rect 13814 18164 13820 18176
rect 13872 18164 13878 18216
rect 15013 18207 15071 18213
rect 15013 18173 15025 18207
rect 15059 18204 15071 18207
rect 15470 18204 15476 18216
rect 15059 18176 15476 18204
rect 15059 18173 15071 18176
rect 15013 18167 15071 18173
rect 15470 18164 15476 18176
rect 15528 18164 15534 18216
rect 15562 18164 15568 18216
rect 15620 18204 15626 18216
rect 18046 18204 18052 18216
rect 15620 18176 18052 18204
rect 15620 18164 15626 18176
rect 18046 18164 18052 18176
rect 18104 18204 18110 18216
rect 18432 18204 18460 18258
rect 18616 18244 19064 18272
rect 19058 18232 19064 18244
rect 19116 18272 19122 18284
rect 19337 18275 19395 18281
rect 19337 18272 19349 18275
rect 19116 18244 19349 18272
rect 19116 18232 19122 18244
rect 19337 18241 19349 18244
rect 19383 18241 19395 18275
rect 19337 18235 19395 18241
rect 19426 18232 19432 18284
rect 19484 18232 19490 18284
rect 19518 18232 19524 18284
rect 19576 18232 19582 18284
rect 19794 18232 19800 18284
rect 19852 18232 19858 18284
rect 20349 18275 20407 18281
rect 20349 18241 20361 18275
rect 20395 18241 20407 18275
rect 20349 18235 20407 18241
rect 18506 18204 18512 18216
rect 18104 18176 18512 18204
rect 18104 18164 18110 18176
rect 18506 18164 18512 18176
rect 18564 18164 18570 18216
rect 19242 18164 19248 18216
rect 19300 18164 19306 18216
rect 20364 18204 20392 18235
rect 20438 18232 20444 18284
rect 20496 18272 20502 18284
rect 20640 18281 20668 18312
rect 20625 18275 20683 18281
rect 20496 18244 20541 18272
rect 20496 18232 20502 18244
rect 20625 18241 20637 18275
rect 20671 18241 20683 18275
rect 20625 18235 20683 18241
rect 20714 18232 20720 18284
rect 20772 18232 20778 18284
rect 20824 18281 20852 18380
rect 20993 18377 21005 18411
rect 21039 18408 21051 18411
rect 25314 18408 25320 18420
rect 21039 18380 25320 18408
rect 21039 18377 21051 18380
rect 20993 18371 21051 18377
rect 25314 18368 25320 18380
rect 25372 18368 25378 18420
rect 25424 18380 28396 18408
rect 23474 18340 23480 18352
rect 22940 18312 23480 18340
rect 22940 18281 22968 18312
rect 23474 18300 23480 18312
rect 23532 18300 23538 18352
rect 24486 18340 24492 18352
rect 24426 18312 24492 18340
rect 24486 18300 24492 18312
rect 24544 18340 24550 18352
rect 24946 18340 24952 18352
rect 24544 18312 24952 18340
rect 24544 18300 24550 18312
rect 24946 18300 24952 18312
rect 25004 18340 25010 18352
rect 25424 18340 25452 18380
rect 25004 18312 25452 18340
rect 25004 18300 25010 18312
rect 20814 18275 20872 18281
rect 20814 18241 20826 18275
rect 20860 18241 20872 18275
rect 20814 18235 20872 18241
rect 22925 18275 22983 18281
rect 22925 18241 22937 18275
rect 22971 18241 22983 18275
rect 28368 18272 28396 18380
rect 28626 18272 28632 18284
rect 28368 18258 28632 18272
rect 28382 18244 28632 18258
rect 22925 18235 22983 18241
rect 28626 18232 28632 18244
rect 28684 18232 28690 18284
rect 19352 18176 20392 18204
rect 12161 18139 12219 18145
rect 12161 18136 12173 18139
rect 10152 18108 12173 18136
rect 12161 18105 12173 18108
rect 12207 18105 12219 18139
rect 14734 18136 14740 18148
rect 12161 18099 12219 18105
rect 12406 18108 14740 18136
rect 5445 18071 5503 18077
rect 5445 18068 5457 18071
rect 5224 18040 5457 18068
rect 5224 18028 5230 18040
rect 5445 18037 5457 18040
rect 5491 18037 5503 18071
rect 5445 18031 5503 18037
rect 6181 18071 6239 18077
rect 6181 18037 6193 18071
rect 6227 18068 6239 18071
rect 7650 18068 7656 18080
rect 6227 18040 7656 18068
rect 6227 18037 6239 18040
rect 6181 18031 6239 18037
rect 7650 18028 7656 18040
rect 7708 18028 7714 18080
rect 9858 18028 9864 18080
rect 9916 18068 9922 18080
rect 9953 18071 10011 18077
rect 9953 18068 9965 18071
rect 9916 18040 9965 18068
rect 9916 18028 9922 18040
rect 9953 18037 9965 18040
rect 9999 18037 10011 18071
rect 9953 18031 10011 18037
rect 10042 18028 10048 18080
rect 10100 18028 10106 18080
rect 10134 18028 10140 18080
rect 10192 18068 10198 18080
rect 10597 18071 10655 18077
rect 10597 18068 10609 18071
rect 10192 18040 10609 18068
rect 10192 18028 10198 18040
rect 10597 18037 10609 18040
rect 10643 18037 10655 18071
rect 10597 18031 10655 18037
rect 10686 18028 10692 18080
rect 10744 18068 10750 18080
rect 12066 18068 12072 18080
rect 10744 18040 12072 18068
rect 10744 18028 10750 18040
rect 12066 18028 12072 18040
rect 12124 18068 12130 18080
rect 12406 18068 12434 18108
rect 14734 18096 14740 18108
rect 14792 18096 14798 18148
rect 16758 18136 16764 18148
rect 16040 18108 16764 18136
rect 12124 18040 12434 18068
rect 13265 18071 13323 18077
rect 12124 18028 12130 18040
rect 13265 18037 13277 18071
rect 13311 18068 13323 18071
rect 16040 18068 16068 18108
rect 16758 18096 16764 18108
rect 16816 18096 16822 18148
rect 18322 18096 18328 18148
rect 18380 18136 18386 18148
rect 19352 18136 19380 18176
rect 23198 18164 23204 18216
rect 23256 18164 23262 18216
rect 23658 18164 23664 18216
rect 23716 18204 23722 18216
rect 24949 18207 25007 18213
rect 24949 18204 24961 18207
rect 23716 18176 24961 18204
rect 23716 18164 23722 18176
rect 24949 18173 24961 18176
rect 24995 18204 25007 18207
rect 25041 18207 25099 18213
rect 25041 18204 25053 18207
rect 24995 18176 25053 18204
rect 24995 18173 25007 18176
rect 24949 18167 25007 18173
rect 25041 18173 25053 18176
rect 25087 18204 25099 18207
rect 25498 18204 25504 18216
rect 25087 18176 25504 18204
rect 25087 18173 25099 18176
rect 25041 18167 25099 18173
rect 25498 18164 25504 18176
rect 25556 18164 25562 18216
rect 26878 18164 26884 18216
rect 26936 18204 26942 18216
rect 26973 18207 27031 18213
rect 26973 18204 26985 18207
rect 26936 18176 26985 18204
rect 26936 18164 26942 18176
rect 26973 18173 26985 18176
rect 27019 18173 27031 18207
rect 26973 18167 27031 18173
rect 27246 18164 27252 18216
rect 27304 18164 27310 18216
rect 28994 18164 29000 18216
rect 29052 18164 29058 18216
rect 18380 18108 19380 18136
rect 20257 18139 20315 18145
rect 18380 18096 18386 18108
rect 20257 18105 20269 18139
rect 20303 18136 20315 18139
rect 21082 18136 21088 18148
rect 20303 18108 21088 18136
rect 20303 18105 20315 18108
rect 20257 18099 20315 18105
rect 21082 18096 21088 18108
rect 21140 18096 21146 18148
rect 25222 18096 25228 18148
rect 25280 18136 25286 18148
rect 26418 18136 26424 18148
rect 25280 18108 26424 18136
rect 25280 18096 25286 18108
rect 26418 18096 26424 18108
rect 26476 18096 26482 18148
rect 13311 18040 16068 18068
rect 13311 18037 13323 18040
rect 13265 18031 13323 18037
rect 16114 18028 16120 18080
rect 16172 18068 16178 18080
rect 16485 18071 16543 18077
rect 16485 18068 16497 18071
rect 16172 18040 16497 18068
rect 16172 18028 16178 18040
rect 16485 18037 16497 18040
rect 16531 18037 16543 18071
rect 16485 18031 16543 18037
rect 24854 18028 24860 18080
rect 24912 18068 24918 18080
rect 25685 18071 25743 18077
rect 25685 18068 25697 18071
rect 24912 18040 25697 18068
rect 24912 18028 24918 18040
rect 25685 18037 25697 18040
rect 25731 18037 25743 18071
rect 25685 18031 25743 18037
rect 1104 17978 29440 18000
rect 1104 17926 4491 17978
rect 4543 17926 4555 17978
rect 4607 17926 4619 17978
rect 4671 17926 4683 17978
rect 4735 17926 4747 17978
rect 4799 17926 11574 17978
rect 11626 17926 11638 17978
rect 11690 17926 11702 17978
rect 11754 17926 11766 17978
rect 11818 17926 11830 17978
rect 11882 17926 18657 17978
rect 18709 17926 18721 17978
rect 18773 17926 18785 17978
rect 18837 17926 18849 17978
rect 18901 17926 18913 17978
rect 18965 17926 25740 17978
rect 25792 17926 25804 17978
rect 25856 17926 25868 17978
rect 25920 17926 25932 17978
rect 25984 17926 25996 17978
rect 26048 17926 29440 17978
rect 1104 17904 29440 17926
rect 3234 17824 3240 17876
rect 3292 17864 3298 17876
rect 5258 17864 5264 17876
rect 3292 17836 5264 17864
rect 3292 17824 3298 17836
rect 5258 17824 5264 17836
rect 5316 17864 5322 17876
rect 7742 17864 7748 17876
rect 5316 17836 7748 17864
rect 5316 17824 5322 17836
rect 3694 17688 3700 17740
rect 3752 17728 3758 17740
rect 5261 17731 5319 17737
rect 5261 17728 5273 17731
rect 3752 17700 5273 17728
rect 3752 17688 3758 17700
rect 5261 17697 5273 17700
rect 5307 17697 5319 17731
rect 5261 17691 5319 17697
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17660 4491 17663
rect 5166 17660 5172 17672
rect 4479 17632 5172 17660
rect 4479 17629 4491 17632
rect 4433 17623 4491 17629
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 6656 17646 6684 17836
rect 7742 17824 7748 17836
rect 7800 17824 7806 17876
rect 11054 17824 11060 17876
rect 11112 17824 11118 17876
rect 11330 17824 11336 17876
rect 11388 17824 11394 17876
rect 12069 17867 12127 17873
rect 12069 17833 12081 17867
rect 12115 17864 12127 17867
rect 12618 17864 12624 17876
rect 12115 17836 12624 17864
rect 12115 17833 12127 17836
rect 12069 17827 12127 17833
rect 12618 17824 12624 17836
rect 12676 17824 12682 17876
rect 13906 17824 13912 17876
rect 13964 17824 13970 17876
rect 19794 17824 19800 17876
rect 19852 17824 19858 17876
rect 20714 17824 20720 17876
rect 20772 17864 20778 17876
rect 21818 17864 21824 17876
rect 20772 17836 21824 17864
rect 20772 17824 20778 17836
rect 21818 17824 21824 17836
rect 21876 17824 21882 17876
rect 22462 17824 22468 17876
rect 22520 17864 22526 17876
rect 22646 17864 22652 17876
rect 22520 17836 22652 17864
rect 22520 17824 22526 17836
rect 22646 17824 22652 17836
rect 22704 17864 22710 17876
rect 22830 17864 22836 17876
rect 22704 17836 22836 17864
rect 22704 17824 22710 17836
rect 22830 17824 22836 17836
rect 22888 17824 22894 17876
rect 23198 17824 23204 17876
rect 23256 17864 23262 17876
rect 23293 17867 23351 17873
rect 23293 17864 23305 17867
rect 23256 17836 23305 17864
rect 23256 17824 23262 17836
rect 23293 17833 23305 17836
rect 23339 17833 23351 17867
rect 23293 17827 23351 17833
rect 23382 17824 23388 17876
rect 23440 17864 23446 17876
rect 25130 17864 25136 17876
rect 23440 17836 25136 17864
rect 23440 17824 23446 17836
rect 25130 17824 25136 17836
rect 25188 17824 25194 17876
rect 25866 17824 25872 17876
rect 25924 17864 25930 17876
rect 26786 17864 26792 17876
rect 25924 17836 26792 17864
rect 25924 17824 25930 17836
rect 26786 17824 26792 17836
rect 26844 17824 26850 17876
rect 27157 17867 27215 17873
rect 27157 17833 27169 17867
rect 27203 17864 27215 17867
rect 27246 17864 27252 17876
rect 27203 17836 27252 17864
rect 27203 17833 27215 17836
rect 27157 17827 27215 17833
rect 27246 17824 27252 17836
rect 27304 17824 27310 17876
rect 7558 17756 7564 17808
rect 7616 17756 7622 17808
rect 7009 17731 7067 17737
rect 7009 17697 7021 17731
rect 7055 17728 7067 17731
rect 7576 17728 7604 17756
rect 7055 17700 7604 17728
rect 9585 17731 9643 17737
rect 7055 17697 7067 17700
rect 7009 17691 7067 17697
rect 7282 17620 7288 17672
rect 7340 17620 7346 17672
rect 7392 17669 7420 17700
rect 9585 17697 9597 17731
rect 9631 17728 9643 17731
rect 9950 17728 9956 17740
rect 9631 17700 9956 17728
rect 9631 17697 9643 17700
rect 9585 17691 9643 17697
rect 9950 17688 9956 17700
rect 10008 17688 10014 17740
rect 7377 17663 7435 17669
rect 7377 17629 7389 17663
rect 7423 17629 7435 17663
rect 7377 17623 7435 17629
rect 7561 17663 7619 17669
rect 7561 17629 7573 17663
rect 7607 17629 7619 17663
rect 7561 17623 7619 17629
rect 3418 17552 3424 17604
rect 3476 17592 3482 17604
rect 4522 17592 4528 17604
rect 3476 17564 4528 17592
rect 3476 17552 3482 17564
rect 4522 17552 4528 17564
rect 4580 17552 4586 17604
rect 4798 17552 4804 17604
rect 4856 17592 4862 17604
rect 5537 17595 5595 17601
rect 4856 17564 5488 17592
rect 4856 17552 4862 17564
rect 5460 17536 5488 17564
rect 5537 17561 5549 17595
rect 5583 17592 5595 17595
rect 5810 17592 5816 17604
rect 5583 17564 5816 17592
rect 5583 17561 5595 17564
rect 5537 17555 5595 17561
rect 5810 17552 5816 17564
rect 5868 17552 5874 17604
rect 7098 17552 7104 17604
rect 7156 17552 7162 17604
rect 4985 17527 5043 17533
rect 4985 17493 4997 17527
rect 5031 17524 5043 17527
rect 5166 17524 5172 17536
rect 5031 17496 5172 17524
rect 5031 17493 5043 17496
rect 4985 17487 5043 17493
rect 5166 17484 5172 17496
rect 5224 17484 5230 17536
rect 5442 17484 5448 17536
rect 5500 17484 5506 17536
rect 6362 17484 6368 17536
rect 6420 17524 6426 17536
rect 7576 17524 7604 17623
rect 7650 17620 7656 17672
rect 7708 17620 7714 17672
rect 11072 17660 11100 17824
rect 11348 17728 11376 17824
rect 18598 17756 18604 17808
rect 18656 17796 18662 17808
rect 18656 17768 20208 17796
rect 18656 17756 18662 17768
rect 12161 17731 12219 17737
rect 11348 17700 11836 17728
rect 10994 17632 11100 17660
rect 11238 17620 11244 17672
rect 11296 17620 11302 17672
rect 11422 17620 11428 17672
rect 11480 17620 11486 17672
rect 11808 17669 11836 17700
rect 12161 17697 12173 17731
rect 12207 17728 12219 17731
rect 17313 17731 17371 17737
rect 17313 17728 17325 17731
rect 12207 17700 17325 17728
rect 12207 17697 12219 17700
rect 12161 17691 12219 17697
rect 17313 17697 17325 17700
rect 17359 17728 17371 17731
rect 19334 17728 19340 17740
rect 17359 17700 19340 17728
rect 17359 17697 17371 17700
rect 17313 17691 17371 17697
rect 19334 17688 19340 17700
rect 19392 17728 19398 17740
rect 20073 17731 20131 17737
rect 20073 17728 20085 17731
rect 19392 17700 20085 17728
rect 19392 17688 19398 17700
rect 20073 17697 20085 17700
rect 20119 17697 20131 17731
rect 20180 17728 20208 17768
rect 23308 17768 23888 17796
rect 22373 17731 22431 17737
rect 20180 17700 21496 17728
rect 20073 17691 20131 17697
rect 11974 17669 11980 17672
rect 11518 17663 11576 17669
rect 11518 17629 11530 17663
rect 11564 17629 11576 17663
rect 11518 17623 11576 17629
rect 11793 17663 11851 17669
rect 11793 17629 11805 17663
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 11931 17663 11980 17669
rect 11931 17629 11943 17663
rect 11977 17629 11980 17663
rect 11931 17623 11980 17629
rect 9861 17595 9919 17601
rect 9861 17561 9873 17595
rect 9907 17592 9919 17595
rect 10134 17592 10140 17604
rect 9907 17564 10140 17592
rect 9907 17561 9919 17564
rect 9861 17555 9919 17561
rect 10134 17552 10140 17564
rect 10192 17552 10198 17604
rect 11146 17552 11152 17604
rect 11204 17552 11210 17604
rect 11256 17592 11284 17620
rect 11532 17592 11560 17623
rect 11974 17620 11980 17623
rect 12032 17620 12038 17672
rect 16114 17620 16120 17672
rect 16172 17620 16178 17672
rect 18598 17620 18604 17672
rect 18656 17660 18662 17672
rect 19245 17663 19303 17669
rect 19245 17660 19257 17663
rect 18656 17632 18722 17660
rect 18892 17632 19257 17660
rect 18656 17620 18662 17632
rect 11256 17564 11560 17592
rect 11701 17595 11759 17601
rect 11701 17561 11713 17595
rect 11747 17561 11759 17595
rect 11701 17555 11759 17561
rect 12437 17595 12495 17601
rect 12437 17561 12449 17595
rect 12483 17561 12495 17595
rect 12437 17555 12495 17561
rect 6420 17496 7604 17524
rect 11164 17524 11192 17552
rect 11716 17524 11744 17555
rect 11164 17496 11744 17524
rect 12452 17524 12480 17555
rect 13170 17552 13176 17604
rect 13228 17552 13234 17604
rect 14182 17552 14188 17604
rect 14240 17552 14246 17604
rect 15933 17595 15991 17601
rect 15933 17561 15945 17595
rect 15979 17592 15991 17595
rect 15979 17564 16436 17592
rect 15979 17561 15991 17564
rect 15933 17555 15991 17561
rect 16408 17536 16436 17564
rect 17586 17552 17592 17604
rect 17644 17552 17650 17604
rect 14642 17524 14648 17536
rect 12452 17496 14648 17524
rect 6420 17484 6426 17496
rect 14642 17484 14648 17496
rect 14700 17484 14706 17536
rect 16390 17484 16396 17536
rect 16448 17484 16454 17536
rect 16666 17484 16672 17536
rect 16724 17484 16730 17536
rect 17126 17484 17132 17536
rect 17184 17524 17190 17536
rect 17862 17524 17868 17536
rect 17184 17496 17868 17524
rect 17184 17484 17190 17496
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 18414 17484 18420 17536
rect 18472 17524 18478 17536
rect 18892 17524 18920 17632
rect 19245 17629 19257 17632
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17629 19487 17663
rect 19429 17623 19487 17629
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17660 19671 17663
rect 19978 17660 19984 17672
rect 19659 17632 19984 17660
rect 19659 17629 19671 17632
rect 19613 17623 19671 17629
rect 19444 17536 19472 17623
rect 19978 17620 19984 17632
rect 20036 17620 20042 17672
rect 21468 17646 21496 17700
rect 22373 17697 22385 17731
rect 22419 17728 22431 17731
rect 22646 17728 22652 17740
rect 22419 17700 22652 17728
rect 22419 17697 22431 17700
rect 22373 17691 22431 17697
rect 22646 17688 22652 17700
rect 22704 17728 22710 17740
rect 22925 17731 22983 17737
rect 22925 17728 22937 17731
rect 22704 17700 22937 17728
rect 22704 17688 22710 17700
rect 22925 17697 22937 17700
rect 22971 17697 22983 17731
rect 22925 17691 22983 17697
rect 23308 17672 23336 17768
rect 23750 17728 23756 17740
rect 23492 17700 23756 17728
rect 22281 17663 22339 17669
rect 22281 17629 22293 17663
rect 22327 17660 22339 17663
rect 22462 17660 22468 17672
rect 22327 17632 22468 17660
rect 22327 17629 22339 17632
rect 22281 17623 22339 17629
rect 22462 17620 22468 17632
rect 22520 17620 22526 17672
rect 22554 17620 22560 17672
rect 22612 17660 22618 17672
rect 22741 17663 22799 17669
rect 22741 17660 22753 17663
rect 22612 17632 22753 17660
rect 22612 17620 22618 17632
rect 22741 17629 22753 17632
rect 22787 17629 22799 17663
rect 22741 17623 22799 17629
rect 23017 17663 23075 17669
rect 23017 17629 23029 17663
rect 23063 17629 23075 17663
rect 23017 17623 23075 17629
rect 19521 17595 19579 17601
rect 19521 17561 19533 17595
rect 19567 17592 19579 17595
rect 20254 17592 20260 17604
rect 19567 17564 20260 17592
rect 19567 17561 19579 17564
rect 19521 17555 19579 17561
rect 20254 17552 20260 17564
rect 20312 17552 20318 17604
rect 20346 17552 20352 17604
rect 20404 17552 20410 17604
rect 21818 17552 21824 17604
rect 21876 17592 21882 17604
rect 23032 17592 23060 17623
rect 23290 17620 23296 17672
rect 23348 17620 23354 17672
rect 23492 17669 23520 17700
rect 23750 17688 23756 17700
rect 23808 17688 23814 17740
rect 23477 17663 23535 17669
rect 23477 17629 23489 17663
rect 23523 17629 23535 17663
rect 23860 17660 23888 17768
rect 25498 17756 25504 17808
rect 25556 17796 25562 17808
rect 25556 17768 26188 17796
rect 25556 17756 25562 17768
rect 23937 17731 23995 17737
rect 23937 17697 23949 17731
rect 23983 17728 23995 17731
rect 24854 17728 24860 17740
rect 23983 17700 24860 17728
rect 23983 17697 23995 17700
rect 23937 17691 23995 17697
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 26160 17737 26188 17768
rect 26234 17756 26240 17808
rect 26292 17796 26298 17808
rect 26694 17796 26700 17808
rect 26292 17768 26700 17796
rect 26292 17756 26298 17768
rect 26694 17756 26700 17768
rect 26752 17756 26758 17808
rect 26970 17756 26976 17808
rect 27028 17796 27034 17808
rect 27890 17796 27896 17808
rect 27028 17768 27896 17796
rect 27028 17756 27034 17768
rect 25041 17731 25099 17737
rect 25041 17697 25053 17731
rect 25087 17728 25099 17731
rect 25777 17731 25835 17737
rect 25777 17728 25789 17731
rect 25087 17700 25789 17728
rect 25087 17697 25099 17700
rect 25041 17691 25099 17697
rect 25777 17697 25789 17700
rect 25823 17697 25835 17731
rect 25777 17691 25835 17697
rect 26145 17731 26203 17737
rect 26145 17697 26157 17731
rect 26191 17697 26203 17731
rect 26145 17691 26203 17697
rect 26418 17688 26424 17740
rect 26476 17688 26482 17740
rect 26510 17688 26516 17740
rect 26568 17728 26574 17740
rect 27080 17728 27108 17768
rect 27890 17756 27896 17768
rect 27948 17796 27954 17808
rect 27948 17768 28396 17796
rect 27948 17756 27954 17768
rect 26568 17700 27108 17728
rect 26568 17688 26574 17700
rect 24397 17663 24455 17669
rect 24397 17660 24409 17663
rect 23860 17632 24409 17660
rect 23477 17623 23535 17629
rect 24397 17629 24409 17632
rect 24443 17660 24455 17663
rect 24762 17660 24768 17672
rect 24443 17632 24768 17660
rect 24443 17629 24455 17632
rect 24397 17623 24455 17629
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 25130 17620 25136 17672
rect 25188 17620 25194 17672
rect 25314 17620 25320 17672
rect 25372 17620 25378 17672
rect 25501 17663 25559 17669
rect 25501 17629 25513 17663
rect 25547 17660 25559 17663
rect 25866 17660 25872 17672
rect 25547 17632 25872 17660
rect 25547 17629 25559 17632
rect 25501 17623 25559 17629
rect 25866 17620 25872 17632
rect 25924 17620 25930 17672
rect 25958 17620 25964 17672
rect 26016 17660 26022 17672
rect 26053 17663 26111 17669
rect 26053 17660 26065 17663
rect 26016 17632 26065 17660
rect 26016 17620 26022 17632
rect 26053 17629 26065 17632
rect 26099 17629 26111 17663
rect 26053 17623 26111 17629
rect 26602 17620 26608 17672
rect 26660 17620 26666 17672
rect 26973 17663 27031 17669
rect 26973 17660 26985 17663
rect 26712 17632 26985 17660
rect 21876 17564 23060 17592
rect 21876 17552 21882 17564
rect 23566 17552 23572 17604
rect 23624 17552 23630 17604
rect 23661 17595 23719 17601
rect 23661 17561 23673 17595
rect 23707 17561 23719 17595
rect 23661 17555 23719 17561
rect 23799 17595 23857 17601
rect 23799 17561 23811 17595
rect 23845 17592 23857 17595
rect 24026 17592 24032 17604
rect 23845 17564 24032 17592
rect 23845 17561 23857 17564
rect 23799 17555 23857 17561
rect 18472 17496 18920 17524
rect 18472 17484 18478 17496
rect 19058 17484 19064 17536
rect 19116 17484 19122 17536
rect 19426 17484 19432 17536
rect 19484 17484 19490 17536
rect 22557 17527 22615 17533
rect 22557 17493 22569 17527
rect 22603 17524 22615 17527
rect 23106 17524 23112 17536
rect 22603 17496 23112 17524
rect 22603 17493 22615 17496
rect 22557 17487 22615 17493
rect 23106 17484 23112 17496
rect 23164 17484 23170 17536
rect 23676 17524 23704 17555
rect 24026 17552 24032 17564
rect 24084 17592 24090 17604
rect 24084 17564 24992 17592
rect 24084 17552 24090 17564
rect 24854 17524 24860 17536
rect 23676 17496 24860 17524
rect 24854 17484 24860 17496
rect 24912 17484 24918 17536
rect 24964 17524 24992 17564
rect 25406 17552 25412 17604
rect 25464 17552 25470 17604
rect 25639 17595 25697 17601
rect 25639 17592 25651 17595
rect 25516 17564 25651 17592
rect 25516 17524 25544 17564
rect 25639 17561 25651 17564
rect 25685 17592 25697 17595
rect 26712 17592 26740 17632
rect 26973 17629 26985 17632
rect 27019 17629 27031 17663
rect 26973 17623 27031 17629
rect 25685 17564 26740 17592
rect 25685 17561 25697 17564
rect 25639 17555 25697 17561
rect 26786 17552 26792 17604
rect 26844 17552 26850 17604
rect 26881 17595 26939 17601
rect 26881 17561 26893 17595
rect 26927 17592 26939 17595
rect 27080 17592 27108 17700
rect 28368 17728 28396 17768
rect 28442 17728 28448 17740
rect 28368 17700 28448 17728
rect 27154 17620 27160 17672
rect 27212 17660 27218 17672
rect 28368 17669 28396 17700
rect 28442 17688 28448 17700
rect 28500 17728 28506 17740
rect 28994 17728 29000 17740
rect 28500 17700 29000 17728
rect 28500 17688 28506 17700
rect 28994 17688 29000 17700
rect 29052 17688 29058 17740
rect 27893 17663 27951 17669
rect 27893 17660 27905 17663
rect 27212 17632 27905 17660
rect 27212 17620 27218 17632
rect 27893 17629 27905 17632
rect 27939 17629 27951 17663
rect 27893 17623 27951 17629
rect 28169 17663 28227 17669
rect 28169 17629 28181 17663
rect 28215 17629 28227 17663
rect 28169 17623 28227 17629
rect 28353 17663 28411 17669
rect 28353 17629 28365 17663
rect 28399 17629 28411 17663
rect 28353 17623 28411 17629
rect 26927 17564 27108 17592
rect 27433 17595 27491 17601
rect 26927 17561 26939 17564
rect 26881 17555 26939 17561
rect 27433 17561 27445 17595
rect 27479 17561 27491 17595
rect 27433 17555 27491 17561
rect 24964 17496 25544 17524
rect 25869 17527 25927 17533
rect 25869 17493 25881 17527
rect 25915 17524 25927 17527
rect 26142 17524 26148 17536
rect 25915 17496 26148 17524
rect 25915 17493 25927 17496
rect 25869 17487 25927 17493
rect 26142 17484 26148 17496
rect 26200 17484 26206 17536
rect 26234 17484 26240 17536
rect 26292 17484 26298 17536
rect 26418 17484 26424 17536
rect 26476 17524 26482 17536
rect 27448 17524 27476 17555
rect 27522 17552 27528 17604
rect 27580 17592 27586 17604
rect 27617 17595 27675 17601
rect 27617 17592 27629 17595
rect 27580 17564 27629 17592
rect 27580 17552 27586 17564
rect 27617 17561 27629 17564
rect 27663 17561 27675 17595
rect 28184 17592 28212 17623
rect 27617 17555 27675 17561
rect 27816 17564 28396 17592
rect 26476 17496 27476 17524
rect 26476 17484 26482 17496
rect 27706 17484 27712 17536
rect 27764 17524 27770 17536
rect 27816 17533 27844 17564
rect 28368 17536 28396 17564
rect 27801 17527 27859 17533
rect 27801 17524 27813 17527
rect 27764 17496 27813 17524
rect 27764 17484 27770 17496
rect 27801 17493 27813 17496
rect 27847 17493 27859 17527
rect 27801 17487 27859 17493
rect 27982 17484 27988 17536
rect 28040 17484 28046 17536
rect 28074 17484 28080 17536
rect 28132 17524 28138 17536
rect 28261 17527 28319 17533
rect 28261 17524 28273 17527
rect 28132 17496 28273 17524
rect 28132 17484 28138 17496
rect 28261 17493 28273 17496
rect 28307 17493 28319 17527
rect 28261 17487 28319 17493
rect 28350 17484 28356 17536
rect 28408 17484 28414 17536
rect 1104 17434 29595 17456
rect 1104 17382 8032 17434
rect 8084 17382 8096 17434
rect 8148 17382 8160 17434
rect 8212 17382 8224 17434
rect 8276 17382 8288 17434
rect 8340 17382 15115 17434
rect 15167 17382 15179 17434
rect 15231 17382 15243 17434
rect 15295 17382 15307 17434
rect 15359 17382 15371 17434
rect 15423 17382 22198 17434
rect 22250 17382 22262 17434
rect 22314 17382 22326 17434
rect 22378 17382 22390 17434
rect 22442 17382 22454 17434
rect 22506 17382 29281 17434
rect 29333 17382 29345 17434
rect 29397 17382 29409 17434
rect 29461 17382 29473 17434
rect 29525 17382 29537 17434
rect 29589 17382 29595 17434
rect 1104 17360 29595 17382
rect 3694 17320 3700 17332
rect 3528 17292 3700 17320
rect 3528 17261 3556 17292
rect 3694 17280 3700 17292
rect 3752 17280 3758 17332
rect 4338 17320 4344 17332
rect 3804 17292 4344 17320
rect 3513 17255 3571 17261
rect 3513 17221 3525 17255
rect 3559 17221 3571 17255
rect 3513 17215 3571 17221
rect 3804 17196 3832 17292
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 4522 17280 4528 17332
rect 4580 17280 4586 17332
rect 5074 17280 5080 17332
rect 5132 17320 5138 17332
rect 5169 17323 5227 17329
rect 5169 17320 5181 17323
rect 5132 17292 5181 17320
rect 5132 17280 5138 17292
rect 5169 17289 5181 17292
rect 5215 17289 5227 17323
rect 5169 17283 5227 17289
rect 5276 17292 6040 17320
rect 4798 17212 4804 17264
rect 4856 17212 4862 17264
rect 5276 17252 5304 17292
rect 5092 17224 5304 17252
rect 3329 17187 3387 17193
rect 3329 17153 3341 17187
rect 3375 17153 3387 17187
rect 3329 17147 3387 17153
rect 3605 17187 3663 17193
rect 3605 17153 3617 17187
rect 3651 17153 3663 17187
rect 3605 17147 3663 17153
rect 3697 17187 3755 17193
rect 3697 17153 3709 17187
rect 3743 17184 3755 17187
rect 3786 17184 3792 17196
rect 3743 17156 3792 17184
rect 3743 17153 3755 17156
rect 3697 17147 3755 17153
rect 3344 17048 3372 17147
rect 3510 17076 3516 17128
rect 3568 17116 3574 17128
rect 3620 17116 3648 17147
rect 3786 17144 3792 17156
rect 3844 17144 3850 17196
rect 3970 17144 3976 17196
rect 4028 17144 4034 17196
rect 4062 17144 4068 17196
rect 4120 17184 4126 17196
rect 4157 17187 4215 17193
rect 4157 17184 4169 17187
rect 4120 17156 4169 17184
rect 4120 17144 4126 17156
rect 4157 17153 4169 17156
rect 4203 17153 4215 17187
rect 4157 17147 4215 17153
rect 4246 17144 4252 17196
rect 4304 17144 4310 17196
rect 4338 17144 4344 17196
rect 4396 17193 4402 17196
rect 4396 17187 4423 17193
rect 4411 17153 4423 17187
rect 4396 17147 4423 17153
rect 4396 17144 4402 17147
rect 4522 17144 4528 17196
rect 4580 17144 4586 17196
rect 4617 17187 4675 17193
rect 4617 17153 4629 17187
rect 4663 17153 4675 17187
rect 4617 17147 4675 17153
rect 4893 17187 4951 17193
rect 4893 17153 4905 17187
rect 4939 17153 4951 17187
rect 4893 17147 4951 17153
rect 4985 17187 5043 17193
rect 4985 17153 4997 17187
rect 5031 17184 5043 17187
rect 5092 17184 5120 17224
rect 5442 17212 5448 17264
rect 5500 17252 5506 17264
rect 5500 17224 5948 17252
rect 5500 17212 5506 17224
rect 5920 17196 5948 17224
rect 6012 17196 6040 17292
rect 9950 17280 9956 17332
rect 10008 17320 10014 17332
rect 12802 17320 12808 17332
rect 10008 17292 12204 17320
rect 10008 17280 10014 17292
rect 9968 17252 9996 17280
rect 9600 17224 9996 17252
rect 5031 17156 5120 17184
rect 5031 17153 5043 17156
rect 4985 17147 5043 17153
rect 4540 17116 4568 17144
rect 3568 17088 4568 17116
rect 4632 17116 4660 17147
rect 4798 17116 4804 17128
rect 4632 17088 4804 17116
rect 3568 17076 3574 17088
rect 4798 17076 4804 17088
rect 4856 17076 4862 17128
rect 4908 17116 4936 17147
rect 5258 17144 5264 17196
rect 5316 17144 5322 17196
rect 5534 17144 5540 17196
rect 5592 17144 5598 17196
rect 5629 17187 5687 17193
rect 5629 17153 5641 17187
rect 5675 17153 5687 17187
rect 5629 17147 5687 17153
rect 5644 17116 5672 17147
rect 5902 17144 5908 17196
rect 5960 17144 5966 17196
rect 5994 17144 6000 17196
rect 6052 17144 6058 17196
rect 9600 17193 9628 17224
rect 11330 17212 11336 17264
rect 11388 17252 11394 17264
rect 11882 17252 11888 17264
rect 11388 17224 11888 17252
rect 11388 17212 11394 17224
rect 11882 17212 11888 17224
rect 11940 17212 11946 17264
rect 12176 17193 12204 17292
rect 12452 17292 12808 17320
rect 12452 17261 12480 17292
rect 12802 17280 12808 17292
rect 12860 17280 12866 17332
rect 13814 17280 13820 17332
rect 13872 17320 13878 17332
rect 13909 17323 13967 17329
rect 13909 17320 13921 17323
rect 13872 17292 13921 17320
rect 13872 17280 13878 17292
rect 13909 17289 13921 17292
rect 13955 17289 13967 17323
rect 16666 17320 16672 17332
rect 13909 17283 13967 17289
rect 15028 17292 16672 17320
rect 12437 17255 12495 17261
rect 12437 17221 12449 17255
rect 12483 17221 12495 17255
rect 12437 17215 12495 17221
rect 13170 17212 13176 17264
rect 13228 17212 13234 17264
rect 9585 17187 9643 17193
rect 9585 17153 9597 17187
rect 9631 17153 9643 17187
rect 12161 17187 12219 17193
rect 9585 17147 9643 17153
rect 6012 17116 6040 17144
rect 4908 17088 5120 17116
rect 5644 17088 6040 17116
rect 5092 17048 5120 17088
rect 9858 17076 9864 17128
rect 9916 17076 9922 17128
rect 10980 17116 11008 17170
rect 12161 17153 12173 17187
rect 12207 17153 12219 17187
rect 12161 17147 12219 17153
rect 13906 17144 13912 17196
rect 13964 17184 13970 17196
rect 15028 17193 15056 17292
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 16758 17280 16764 17332
rect 16816 17320 16822 17332
rect 16816 17292 17356 17320
rect 16816 17280 16822 17292
rect 15197 17255 15255 17261
rect 15197 17221 15209 17255
rect 15243 17252 15255 17255
rect 16022 17252 16028 17264
rect 15243 17224 16028 17252
rect 15243 17221 15255 17224
rect 15197 17215 15255 17221
rect 15856 17196 15884 17224
rect 16022 17212 16028 17224
rect 16080 17212 16086 17264
rect 16114 17212 16120 17264
rect 16172 17252 16178 17264
rect 16172 17224 17080 17252
rect 16172 17212 16178 17224
rect 14001 17187 14059 17193
rect 14001 17184 14013 17187
rect 13964 17156 14013 17184
rect 13964 17144 13970 17156
rect 14001 17153 14013 17156
rect 14047 17153 14059 17187
rect 14001 17147 14059 17153
rect 15013 17187 15071 17193
rect 15013 17153 15025 17187
rect 15059 17153 15071 17187
rect 15013 17147 15071 17153
rect 15102 17144 15108 17196
rect 15160 17184 15166 17196
rect 15289 17187 15347 17193
rect 15289 17184 15301 17187
rect 15160 17156 15301 17184
rect 15160 17144 15166 17156
rect 15289 17153 15301 17156
rect 15335 17153 15347 17187
rect 15289 17147 15347 17153
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17153 15439 17187
rect 15381 17147 15439 17153
rect 11054 17116 11060 17128
rect 10980 17088 11060 17116
rect 11054 17076 11060 17088
rect 11112 17076 11118 17128
rect 5166 17048 5172 17060
rect 3344 17020 5028 17048
rect 5092 17020 5172 17048
rect 5000 16992 5028 17020
rect 5166 17008 5172 17020
rect 5224 17008 5230 17060
rect 5258 17008 5264 17060
rect 5316 17048 5322 17060
rect 5316 17020 7788 17048
rect 5316 17008 5322 17020
rect 7760 16992 7788 17020
rect 11238 17008 11244 17060
rect 11296 17048 11302 17060
rect 11333 17051 11391 17057
rect 11333 17048 11345 17051
rect 11296 17020 11345 17048
rect 11296 17008 11302 17020
rect 11333 17017 11345 17020
rect 11379 17017 11391 17051
rect 11333 17011 11391 17017
rect 3326 16940 3332 16992
rect 3384 16980 3390 16992
rect 3881 16983 3939 16989
rect 3881 16980 3893 16983
rect 3384 16952 3893 16980
rect 3384 16940 3390 16952
rect 3881 16949 3893 16952
rect 3927 16949 3939 16983
rect 3881 16943 3939 16949
rect 4982 16940 4988 16992
rect 5040 16940 5046 16992
rect 5810 16940 5816 16992
rect 5868 16940 5874 16992
rect 7742 16940 7748 16992
rect 7800 16940 7806 16992
rect 14090 16940 14096 16992
rect 14148 16980 14154 16992
rect 14645 16983 14703 16989
rect 14645 16980 14657 16983
rect 14148 16952 14657 16980
rect 14148 16940 14154 16952
rect 14645 16949 14657 16952
rect 14691 16949 14703 16983
rect 15396 16980 15424 17147
rect 15838 17144 15844 17196
rect 15896 17144 15902 17196
rect 17052 17193 17080 17224
rect 16945 17187 17003 17193
rect 16945 17184 16957 17187
rect 16592 17156 16957 17184
rect 15470 17076 15476 17128
rect 15528 17076 15534 17128
rect 15488 17048 15516 17076
rect 15565 17051 15623 17057
rect 15565 17048 15577 17051
rect 15488 17020 15577 17048
rect 15565 17017 15577 17020
rect 15611 17017 15623 17051
rect 15856 17048 15884 17144
rect 16592 17128 16620 17156
rect 16945 17153 16957 17156
rect 16991 17153 17003 17187
rect 16945 17147 17003 17153
rect 17037 17187 17095 17193
rect 17037 17153 17049 17187
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 17126 17144 17132 17196
rect 17184 17144 17190 17196
rect 17328 17193 17356 17292
rect 17586 17280 17592 17332
rect 17644 17320 17650 17332
rect 18785 17323 18843 17329
rect 18785 17320 18797 17323
rect 17644 17292 18797 17320
rect 17644 17280 17650 17292
rect 18785 17289 18797 17292
rect 18831 17289 18843 17323
rect 19058 17320 19064 17332
rect 18785 17283 18843 17289
rect 18892 17292 19064 17320
rect 18892 17261 18920 17292
rect 19058 17280 19064 17292
rect 19116 17280 19122 17332
rect 19242 17280 19248 17332
rect 19300 17280 19306 17332
rect 20346 17280 20352 17332
rect 20404 17320 20410 17332
rect 20809 17323 20867 17329
rect 20809 17320 20821 17323
rect 20404 17292 20821 17320
rect 20404 17280 20410 17292
rect 20809 17289 20821 17292
rect 20855 17289 20867 17323
rect 20809 17283 20867 17289
rect 21821 17323 21879 17329
rect 21821 17289 21833 17323
rect 21867 17289 21879 17323
rect 22830 17320 22836 17332
rect 21821 17283 21879 17289
rect 22388 17292 22836 17320
rect 18877 17255 18935 17261
rect 18877 17252 18889 17255
rect 17604 17224 18889 17252
rect 17604 17193 17632 17224
rect 18877 17221 18889 17224
rect 18923 17221 18935 17255
rect 21836 17252 21864 17283
rect 18877 17215 18935 17221
rect 21008 17224 21864 17252
rect 22066 17224 22324 17252
rect 17313 17187 17371 17193
rect 17313 17153 17325 17187
rect 17359 17153 17371 17187
rect 17313 17147 17371 17153
rect 17589 17187 17647 17193
rect 17589 17153 17601 17187
rect 17635 17153 17647 17187
rect 17589 17147 17647 17153
rect 18141 17187 18199 17193
rect 18141 17153 18153 17187
rect 18187 17184 18199 17187
rect 18233 17187 18291 17193
rect 18233 17184 18245 17187
rect 18187 17156 18245 17184
rect 18187 17153 18199 17156
rect 18141 17147 18199 17153
rect 18233 17153 18245 17156
rect 18279 17153 18291 17187
rect 18233 17147 18291 17153
rect 18322 17144 18328 17196
rect 18380 17144 18386 17196
rect 18417 17187 18475 17193
rect 18417 17153 18429 17187
rect 18463 17153 18475 17187
rect 18417 17147 18475 17153
rect 16574 17076 16580 17128
rect 16632 17076 16638 17128
rect 16669 17119 16727 17125
rect 16669 17085 16681 17119
rect 16715 17116 16727 17119
rect 18340 17116 18368 17144
rect 16715 17088 18368 17116
rect 16715 17085 16727 17088
rect 16669 17079 16727 17085
rect 18432 17048 18460 17147
rect 18506 17144 18512 17196
rect 18564 17144 18570 17196
rect 18601 17187 18659 17193
rect 18601 17153 18613 17187
rect 18647 17153 18659 17187
rect 18601 17147 18659 17153
rect 15856 17020 18460 17048
rect 15565 17011 15623 17017
rect 16482 16980 16488 16992
rect 15396 16952 16488 16980
rect 14645 16943 14703 16949
rect 16482 16940 16488 16952
rect 16540 16980 16546 16992
rect 18616 16980 18644 17147
rect 19058 17144 19064 17196
rect 19116 17144 19122 17196
rect 21008 17193 21036 17224
rect 20993 17187 21051 17193
rect 20993 17153 21005 17187
rect 21039 17153 21051 17187
rect 20993 17147 21051 17153
rect 21269 17187 21327 17193
rect 21269 17153 21281 17187
rect 21315 17184 21327 17187
rect 21818 17184 21824 17196
rect 21315 17156 21824 17184
rect 21315 17153 21327 17156
rect 21269 17147 21327 17153
rect 21818 17144 21824 17156
rect 21876 17184 21882 17196
rect 22066 17184 22094 17224
rect 21876 17156 22094 17184
rect 21876 17144 21882 17156
rect 22186 17144 22192 17196
rect 22244 17144 22250 17196
rect 22296 17193 22324 17224
rect 22281 17187 22339 17193
rect 22281 17153 22293 17187
rect 22327 17153 22339 17187
rect 22281 17147 22339 17153
rect 21361 17119 21419 17125
rect 21361 17085 21373 17119
rect 21407 17116 21419 17119
rect 22388 17116 22416 17292
rect 22830 17280 22836 17292
rect 22888 17280 22894 17332
rect 23385 17323 23443 17329
rect 23385 17289 23397 17323
rect 23431 17320 23443 17323
rect 23566 17320 23572 17332
rect 23431 17292 23572 17320
rect 23431 17289 23443 17292
rect 23385 17283 23443 17289
rect 23566 17280 23572 17292
rect 23624 17280 23630 17332
rect 25130 17320 25136 17332
rect 23768 17292 25136 17320
rect 22554 17212 22560 17264
rect 22612 17252 22618 17264
rect 23658 17252 23664 17264
rect 22612 17224 23664 17252
rect 22612 17212 22618 17224
rect 23658 17212 23664 17224
rect 23716 17212 23722 17264
rect 23768 17261 23796 17292
rect 25130 17280 25136 17292
rect 25188 17280 25194 17332
rect 25406 17280 25412 17332
rect 25464 17320 25470 17332
rect 25869 17323 25927 17329
rect 25869 17320 25881 17323
rect 25464 17292 25881 17320
rect 25464 17280 25470 17292
rect 25869 17289 25881 17292
rect 25915 17289 25927 17323
rect 25869 17283 25927 17289
rect 26234 17280 26240 17332
rect 26292 17280 26298 17332
rect 26602 17280 26608 17332
rect 26660 17320 26666 17332
rect 26973 17323 27031 17329
rect 26973 17320 26985 17323
rect 26660 17292 26985 17320
rect 26660 17280 26666 17292
rect 26973 17289 26985 17292
rect 27019 17289 27031 17323
rect 26973 17283 27031 17289
rect 27540 17292 28028 17320
rect 23753 17255 23811 17261
rect 23753 17221 23765 17255
rect 23799 17221 23811 17255
rect 23753 17215 23811 17221
rect 25498 17212 25504 17264
rect 25556 17252 25562 17264
rect 25593 17255 25651 17261
rect 25593 17252 25605 17255
rect 25556 17224 25605 17252
rect 25556 17212 25562 17224
rect 25593 17221 25605 17224
rect 25639 17221 25651 17255
rect 26252 17252 26280 17280
rect 27540 17264 27568 17292
rect 26252 17224 27476 17252
rect 25593 17215 25651 17221
rect 22830 17144 22836 17196
rect 22888 17144 22894 17196
rect 23474 17144 23480 17196
rect 23532 17144 23538 17196
rect 24762 17144 24768 17196
rect 24820 17144 24826 17196
rect 21407 17088 22416 17116
rect 22465 17119 22523 17125
rect 21407 17085 21419 17088
rect 21361 17079 21419 17085
rect 22465 17085 22477 17119
rect 22511 17085 22523 17119
rect 22465 17079 22523 17085
rect 23109 17119 23167 17125
rect 23109 17085 23121 17119
rect 23155 17116 23167 17119
rect 23382 17116 23388 17128
rect 23155 17088 23388 17116
rect 23155 17085 23167 17088
rect 23109 17079 23167 17085
rect 21637 17051 21695 17057
rect 21637 17017 21649 17051
rect 21683 17048 21695 17051
rect 22278 17048 22284 17060
rect 21683 17020 22284 17048
rect 21683 17017 21695 17020
rect 21637 17011 21695 17017
rect 22278 17008 22284 17020
rect 22336 17008 22342 17060
rect 22480 17048 22508 17079
rect 23382 17076 23388 17088
rect 23440 17076 23446 17128
rect 24780 17048 24808 17144
rect 24872 17116 24900 17170
rect 25222 17144 25228 17196
rect 25280 17184 25286 17196
rect 25406 17184 25412 17196
rect 25280 17156 25412 17184
rect 25280 17144 25286 17156
rect 25406 17144 25412 17156
rect 25464 17144 25470 17196
rect 26050 17144 26056 17196
rect 26108 17144 26114 17196
rect 26237 17187 26295 17193
rect 26237 17153 26249 17187
rect 26283 17153 26295 17187
rect 26237 17147 26295 17153
rect 26329 17187 26387 17193
rect 26329 17153 26341 17187
rect 26375 17153 26387 17187
rect 26329 17147 26387 17153
rect 26421 17187 26479 17193
rect 26421 17153 26433 17187
rect 26467 17184 26479 17187
rect 27157 17187 27215 17193
rect 26467 17156 27016 17184
rect 26467 17153 26479 17156
rect 26421 17147 26479 17153
rect 24946 17116 24952 17128
rect 24872 17088 24952 17116
rect 24946 17076 24952 17088
rect 25004 17076 25010 17128
rect 25958 17116 25964 17128
rect 25240 17088 25964 17116
rect 25240 17057 25268 17088
rect 25958 17076 25964 17088
rect 26016 17116 26022 17128
rect 26252 17116 26280 17147
rect 26016 17088 26280 17116
rect 26016 17076 26022 17088
rect 25225 17051 25283 17057
rect 25225 17048 25237 17051
rect 22480 17020 23612 17048
rect 24780 17020 25237 17048
rect 23584 16992 23612 17020
rect 25225 17017 25237 17020
rect 25271 17017 25283 17051
rect 25866 17048 25872 17060
rect 25225 17011 25283 17017
rect 25700 17020 25872 17048
rect 16540 16952 18644 16980
rect 16540 16940 16546 16952
rect 23106 16940 23112 16992
rect 23164 16940 23170 16992
rect 23566 16940 23572 16992
rect 23624 16940 23630 16992
rect 24854 16940 24860 16992
rect 24912 16980 24918 16992
rect 25700 16980 25728 17020
rect 25866 17008 25872 17020
rect 25924 17008 25930 17060
rect 26344 17048 26372 17147
rect 26988 17128 27016 17156
rect 27157 17153 27169 17187
rect 27203 17184 27215 17187
rect 27246 17184 27252 17196
rect 27203 17156 27252 17184
rect 27203 17153 27215 17156
rect 27157 17147 27215 17153
rect 27246 17144 27252 17156
rect 27304 17144 27310 17196
rect 27448 17193 27476 17224
rect 27522 17212 27528 17264
rect 27580 17212 27586 17264
rect 27433 17187 27491 17193
rect 27433 17153 27445 17187
rect 27479 17153 27491 17187
rect 27433 17147 27491 17153
rect 27617 17187 27675 17193
rect 27617 17153 27629 17187
rect 27663 17184 27675 17187
rect 27798 17184 27804 17196
rect 27663 17156 27804 17184
rect 27663 17153 27675 17156
rect 27617 17147 27675 17153
rect 27798 17144 27804 17156
rect 27856 17144 27862 17196
rect 27890 17144 27896 17196
rect 27948 17144 27954 17196
rect 28000 17184 28028 17292
rect 28442 17212 28448 17264
rect 28500 17212 28506 17264
rect 28261 17187 28319 17193
rect 28000 17156 28212 17184
rect 26513 17119 26571 17125
rect 26513 17085 26525 17119
rect 26559 17116 26571 17119
rect 26694 17116 26700 17128
rect 26559 17088 26700 17116
rect 26559 17085 26571 17088
rect 26513 17079 26571 17085
rect 26694 17076 26700 17088
rect 26752 17076 26758 17128
rect 26970 17076 26976 17128
rect 27028 17076 27034 17128
rect 27341 17119 27399 17125
rect 27341 17085 27353 17119
rect 27387 17085 27399 17119
rect 27341 17079 27399 17085
rect 26789 17051 26847 17057
rect 26789 17048 26801 17051
rect 26344 17020 26801 17048
rect 26789 17017 26801 17020
rect 26835 17048 26847 17051
rect 27154 17048 27160 17060
rect 26835 17020 27160 17048
rect 26835 17017 26847 17020
rect 26789 17011 26847 17017
rect 27154 17008 27160 17020
rect 27212 17008 27218 17060
rect 27249 17051 27307 17057
rect 27249 17017 27261 17051
rect 27295 17017 27307 17051
rect 27356 17048 27384 17079
rect 27522 17076 27528 17128
rect 27580 17116 27586 17128
rect 28184 17125 28212 17156
rect 28261 17153 28273 17187
rect 28307 17184 28319 17187
rect 28350 17184 28356 17196
rect 28307 17156 28356 17184
rect 28307 17153 28319 17156
rect 28261 17147 28319 17153
rect 28350 17144 28356 17156
rect 28408 17144 28414 17196
rect 28077 17119 28135 17125
rect 28077 17116 28089 17119
rect 27580 17088 28089 17116
rect 27580 17076 27586 17088
rect 28077 17085 28089 17088
rect 28123 17085 28135 17119
rect 28077 17079 28135 17085
rect 28169 17119 28227 17125
rect 28169 17085 28181 17119
rect 28215 17116 28227 17119
rect 28215 17088 28396 17116
rect 28215 17085 28227 17088
rect 28169 17079 28227 17085
rect 27709 17051 27767 17057
rect 27709 17048 27721 17051
rect 27356 17020 27721 17048
rect 27249 17011 27307 17017
rect 27709 17017 27721 17020
rect 27755 17017 27767 17051
rect 27709 17011 27767 17017
rect 24912 16952 25728 16980
rect 25777 16983 25835 16989
rect 24912 16940 24918 16952
rect 25777 16949 25789 16983
rect 25823 16980 25835 16983
rect 26418 16980 26424 16992
rect 25823 16952 26424 16980
rect 25823 16949 25835 16952
rect 25777 16943 25835 16949
rect 26418 16940 26424 16952
rect 26476 16940 26482 16992
rect 26510 16940 26516 16992
rect 26568 16940 26574 16992
rect 27264 16980 27292 17011
rect 28368 16992 28396 17088
rect 28442 17076 28448 17128
rect 28500 17116 28506 17128
rect 28626 17116 28632 17128
rect 28500 17088 28632 17116
rect 28500 17076 28506 17088
rect 28626 17076 28632 17088
rect 28684 17076 28690 17128
rect 27982 16980 27988 16992
rect 27264 16952 27988 16980
rect 27982 16940 27988 16952
rect 28040 16940 28046 16992
rect 28350 16940 28356 16992
rect 28408 16940 28414 16992
rect 28626 16940 28632 16992
rect 28684 16940 28690 16992
rect 1104 16890 29440 16912
rect 1104 16838 4491 16890
rect 4543 16838 4555 16890
rect 4607 16838 4619 16890
rect 4671 16838 4683 16890
rect 4735 16838 4747 16890
rect 4799 16838 11574 16890
rect 11626 16838 11638 16890
rect 11690 16838 11702 16890
rect 11754 16838 11766 16890
rect 11818 16838 11830 16890
rect 11882 16838 18657 16890
rect 18709 16838 18721 16890
rect 18773 16838 18785 16890
rect 18837 16838 18849 16890
rect 18901 16838 18913 16890
rect 18965 16838 25740 16890
rect 25792 16838 25804 16890
rect 25856 16838 25868 16890
rect 25920 16838 25932 16890
rect 25984 16838 25996 16890
rect 26048 16838 29440 16890
rect 1104 16816 29440 16838
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 6273 16779 6331 16785
rect 6273 16776 6285 16779
rect 5592 16748 6285 16776
rect 5592 16736 5598 16748
rect 6273 16745 6285 16748
rect 6319 16745 6331 16779
rect 6273 16739 6331 16745
rect 14642 16736 14648 16788
rect 14700 16736 14706 16788
rect 15102 16736 15108 16788
rect 15160 16776 15166 16788
rect 20438 16776 20444 16788
rect 15160 16748 20444 16776
rect 15160 16736 15166 16748
rect 20438 16736 20444 16748
rect 20496 16736 20502 16788
rect 22005 16779 22063 16785
rect 22005 16745 22017 16779
rect 22051 16776 22063 16779
rect 22186 16776 22192 16788
rect 22051 16748 22192 16776
rect 22051 16745 22063 16748
rect 22005 16739 22063 16745
rect 22186 16736 22192 16748
rect 22244 16736 22250 16788
rect 22278 16736 22284 16788
rect 22336 16776 22342 16788
rect 22373 16779 22431 16785
rect 22373 16776 22385 16779
rect 22336 16748 22385 16776
rect 22336 16736 22342 16748
rect 22373 16745 22385 16748
rect 22419 16745 22431 16779
rect 22373 16739 22431 16745
rect 22554 16736 22560 16788
rect 22612 16776 22618 16788
rect 22741 16779 22799 16785
rect 22741 16776 22753 16779
rect 22612 16748 22753 16776
rect 22612 16736 22618 16748
rect 22741 16745 22753 16748
rect 22787 16745 22799 16779
rect 22741 16739 22799 16745
rect 22830 16736 22836 16788
rect 22888 16776 22894 16788
rect 23109 16779 23167 16785
rect 23109 16776 23121 16779
rect 22888 16748 23121 16776
rect 22888 16736 22894 16748
rect 23109 16745 23121 16748
rect 23155 16745 23167 16779
rect 23109 16739 23167 16745
rect 23750 16736 23756 16788
rect 23808 16736 23814 16788
rect 24397 16779 24455 16785
rect 24397 16745 24409 16779
rect 24443 16776 24455 16779
rect 25314 16776 25320 16788
rect 24443 16748 25320 16776
rect 24443 16745 24455 16748
rect 24397 16739 24455 16745
rect 25314 16736 25320 16748
rect 25372 16736 25378 16788
rect 26145 16779 26203 16785
rect 26145 16745 26157 16779
rect 26191 16776 26203 16779
rect 26786 16776 26792 16788
rect 26191 16748 26792 16776
rect 26191 16745 26203 16748
rect 26145 16739 26203 16745
rect 26786 16736 26792 16748
rect 26844 16736 26850 16788
rect 26970 16736 26976 16788
rect 27028 16776 27034 16788
rect 27065 16779 27123 16785
rect 27065 16776 27077 16779
rect 27028 16748 27077 16776
rect 27028 16736 27034 16748
rect 27065 16745 27077 16748
rect 27111 16776 27123 16779
rect 27522 16776 27528 16788
rect 27111 16748 27528 16776
rect 27111 16745 27123 16748
rect 27065 16739 27123 16745
rect 27522 16736 27528 16748
rect 27580 16736 27586 16788
rect 27798 16736 27804 16788
rect 27856 16736 27862 16788
rect 27890 16736 27896 16788
rect 27948 16776 27954 16788
rect 28261 16779 28319 16785
rect 28261 16776 28273 16779
rect 27948 16748 28273 16776
rect 27948 16736 27954 16748
rect 28261 16745 28273 16748
rect 28307 16745 28319 16779
rect 28261 16739 28319 16745
rect 5074 16668 5080 16720
rect 5132 16708 5138 16720
rect 6914 16708 6920 16720
rect 5132 16680 6920 16708
rect 5132 16668 5138 16680
rect 6914 16668 6920 16680
rect 6972 16668 6978 16720
rect 14366 16668 14372 16720
rect 14424 16708 14430 16720
rect 14550 16708 14556 16720
rect 14424 16680 14556 16708
rect 14424 16668 14430 16680
rect 14550 16668 14556 16680
rect 14608 16708 14614 16720
rect 15120 16708 15148 16736
rect 14608 16680 15148 16708
rect 14608 16668 14614 16680
rect 23290 16668 23296 16720
rect 23348 16708 23354 16720
rect 23661 16711 23719 16717
rect 23661 16708 23673 16711
rect 23348 16680 23673 16708
rect 23348 16668 23354 16680
rect 23661 16677 23673 16680
rect 23707 16677 23719 16711
rect 23661 16671 23719 16677
rect 24964 16680 26188 16708
rect 3145 16643 3203 16649
rect 3145 16609 3157 16643
rect 3191 16640 3203 16643
rect 3789 16643 3847 16649
rect 3789 16640 3801 16643
rect 3191 16612 3801 16640
rect 3191 16609 3203 16612
rect 3145 16603 3203 16609
rect 3789 16609 3801 16612
rect 3835 16609 3847 16643
rect 3789 16603 3847 16609
rect 4246 16600 4252 16652
rect 4304 16640 4310 16652
rect 4890 16640 4896 16652
rect 4304 16612 4896 16640
rect 4304 16600 4310 16612
rect 4890 16600 4896 16612
rect 4948 16640 4954 16652
rect 10689 16643 10747 16649
rect 4948 16612 6500 16640
rect 4948 16600 4954 16612
rect 1394 16532 1400 16584
rect 1452 16532 1458 16584
rect 4985 16575 5043 16581
rect 4985 16541 4997 16575
rect 5031 16541 5043 16575
rect 4985 16535 5043 16541
rect 1670 16464 1676 16516
rect 1728 16464 1734 16516
rect 3878 16504 3884 16516
rect 2898 16476 3884 16504
rect 3878 16464 3884 16476
rect 3936 16464 3942 16516
rect 4430 16396 4436 16448
rect 4488 16396 4494 16448
rect 5000 16436 5028 16535
rect 5074 16532 5080 16584
rect 5132 16572 5138 16584
rect 5276 16581 5304 16612
rect 6472 16584 6500 16612
rect 9784 16612 9996 16640
rect 5169 16575 5227 16581
rect 5169 16572 5181 16575
rect 5132 16544 5181 16572
rect 5132 16532 5138 16544
rect 5169 16541 5181 16544
rect 5215 16541 5227 16575
rect 5169 16535 5227 16541
rect 5261 16575 5319 16581
rect 5261 16541 5273 16575
rect 5307 16541 5319 16575
rect 5261 16535 5319 16541
rect 5350 16532 5356 16584
rect 5408 16532 5414 16584
rect 5718 16532 5724 16584
rect 5776 16532 5782 16584
rect 6454 16532 6460 16584
rect 6512 16532 6518 16584
rect 9674 16532 9680 16584
rect 9732 16572 9738 16584
rect 9784 16572 9812 16612
rect 9732 16544 9812 16572
rect 9732 16532 9738 16544
rect 9858 16532 9864 16584
rect 9916 16532 9922 16584
rect 9968 16572 9996 16612
rect 10689 16609 10701 16643
rect 10735 16640 10747 16643
rect 10962 16640 10968 16652
rect 10735 16612 10968 16640
rect 10735 16609 10747 16612
rect 10689 16603 10747 16609
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 13998 16640 14004 16652
rect 12268 16612 14004 16640
rect 12268 16584 12296 16612
rect 13998 16600 14004 16612
rect 14056 16640 14062 16652
rect 16574 16640 16580 16652
rect 14056 16612 14504 16640
rect 14056 16600 14062 16612
rect 10229 16575 10287 16581
rect 10229 16572 10241 16575
rect 9968 16544 10241 16572
rect 10229 16541 10241 16544
rect 10275 16541 10287 16575
rect 10229 16535 10287 16541
rect 12250 16532 12256 16584
rect 12308 16532 12314 16584
rect 14090 16532 14096 16584
rect 14148 16532 14154 16584
rect 14476 16581 14504 16612
rect 15120 16612 16580 16640
rect 14461 16575 14519 16581
rect 14461 16541 14473 16575
rect 14507 16541 14519 16575
rect 14461 16535 14519 16541
rect 14642 16532 14648 16584
rect 14700 16572 14706 16584
rect 15010 16572 15016 16584
rect 14700 16544 15016 16572
rect 14700 16532 14706 16544
rect 15010 16532 15016 16544
rect 15068 16572 15074 16584
rect 15120 16581 15148 16612
rect 16574 16600 16580 16612
rect 16632 16640 16638 16652
rect 19058 16640 19064 16652
rect 16632 16612 19064 16640
rect 16632 16600 16638 16612
rect 19058 16600 19064 16612
rect 19116 16600 19122 16652
rect 21818 16600 21824 16652
rect 21876 16640 21882 16652
rect 22833 16643 22891 16649
rect 22833 16640 22845 16643
rect 21876 16612 22845 16640
rect 21876 16600 21882 16612
rect 22833 16609 22845 16612
rect 22879 16640 22891 16643
rect 23845 16643 23903 16649
rect 22879 16612 23520 16640
rect 22879 16609 22891 16612
rect 22833 16603 22891 16609
rect 15105 16575 15163 16581
rect 15105 16572 15117 16575
rect 15068 16544 15117 16572
rect 15068 16532 15074 16544
rect 15105 16541 15117 16544
rect 15151 16541 15163 16575
rect 15105 16535 15163 16541
rect 15197 16575 15255 16581
rect 15197 16541 15209 16575
rect 15243 16541 15255 16575
rect 15197 16535 15255 16541
rect 15289 16575 15347 16581
rect 15289 16541 15301 16575
rect 15335 16541 15347 16575
rect 15289 16535 15347 16541
rect 15473 16575 15531 16581
rect 15473 16541 15485 16575
rect 15519 16572 15531 16575
rect 15654 16572 15660 16584
rect 15519 16544 15660 16572
rect 15519 16541 15531 16544
rect 15473 16535 15531 16541
rect 5368 16504 5396 16532
rect 7466 16504 7472 16516
rect 5368 16476 7472 16504
rect 7466 16464 7472 16476
rect 7524 16464 7530 16516
rect 10042 16464 10048 16516
rect 10100 16464 10106 16516
rect 10137 16507 10195 16513
rect 10137 16473 10149 16507
rect 10183 16504 10195 16507
rect 11241 16507 11299 16513
rect 11241 16504 11253 16507
rect 10183 16476 11253 16504
rect 10183 16473 10195 16476
rect 10137 16467 10195 16473
rect 11241 16473 11253 16476
rect 11287 16473 11299 16507
rect 11241 16467 11299 16473
rect 14277 16507 14335 16513
rect 14277 16473 14289 16507
rect 14323 16473 14335 16507
rect 14277 16467 14335 16473
rect 5442 16436 5448 16448
rect 5000 16408 5448 16436
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 5534 16396 5540 16448
rect 5592 16396 5598 16448
rect 9950 16396 9956 16448
rect 10008 16436 10014 16448
rect 10226 16436 10232 16448
rect 10008 16408 10232 16436
rect 10008 16396 10014 16408
rect 10226 16396 10232 16408
rect 10284 16396 10290 16448
rect 10410 16396 10416 16448
rect 10468 16396 10474 16448
rect 10502 16396 10508 16448
rect 10560 16436 10566 16448
rect 12342 16436 12348 16448
rect 10560 16408 12348 16436
rect 10560 16396 10566 16408
rect 12342 16396 12348 16408
rect 12400 16396 12406 16448
rect 12710 16396 12716 16448
rect 12768 16436 12774 16448
rect 14292 16436 14320 16467
rect 14366 16464 14372 16516
rect 14424 16464 14430 16516
rect 14918 16504 14924 16516
rect 14476 16476 14924 16504
rect 14476 16436 14504 16476
rect 14918 16464 14924 16476
rect 14976 16464 14982 16516
rect 15212 16504 15240 16535
rect 15028 16476 15240 16504
rect 15304 16504 15332 16535
rect 15654 16532 15660 16544
rect 15712 16532 15718 16584
rect 22189 16575 22247 16581
rect 22189 16541 22201 16575
rect 22235 16541 22247 16575
rect 22189 16535 22247 16541
rect 22465 16575 22523 16581
rect 22465 16541 22477 16575
rect 22511 16541 22523 16575
rect 22465 16535 22523 16541
rect 15746 16504 15752 16516
rect 15304 16476 15752 16504
rect 15028 16448 15056 16476
rect 15746 16464 15752 16476
rect 15804 16504 15810 16516
rect 17126 16504 17132 16516
rect 15804 16476 17132 16504
rect 15804 16464 15810 16476
rect 17126 16464 17132 16476
rect 17184 16464 17190 16516
rect 12768 16408 14504 16436
rect 12768 16396 12774 16408
rect 14826 16396 14832 16448
rect 14884 16396 14890 16448
rect 15010 16396 15016 16448
rect 15068 16396 15074 16448
rect 22204 16436 22232 16535
rect 22480 16504 22508 16535
rect 22646 16532 22652 16584
rect 22704 16572 22710 16584
rect 23492 16581 23520 16612
rect 23845 16609 23857 16643
rect 23891 16640 23903 16643
rect 23891 16612 23980 16640
rect 23891 16609 23903 16612
rect 23845 16603 23903 16609
rect 23952 16584 23980 16612
rect 22741 16575 22799 16581
rect 22741 16572 22753 16575
rect 22704 16544 22753 16572
rect 22704 16532 22710 16544
rect 22741 16541 22753 16544
rect 22787 16541 22799 16575
rect 22741 16535 22799 16541
rect 23201 16575 23259 16581
rect 23201 16541 23213 16575
rect 23247 16572 23259 16575
rect 23477 16575 23535 16581
rect 23247 16544 23336 16572
rect 23247 16541 23259 16544
rect 23201 16535 23259 16541
rect 22480 16476 23244 16504
rect 23216 16448 23244 16476
rect 23106 16436 23112 16448
rect 22204 16408 23112 16436
rect 23106 16396 23112 16408
rect 23164 16396 23170 16448
rect 23198 16396 23204 16448
rect 23256 16396 23262 16448
rect 23308 16436 23336 16544
rect 23477 16541 23489 16575
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 23569 16575 23627 16581
rect 23569 16541 23581 16575
rect 23615 16572 23627 16575
rect 23658 16572 23664 16584
rect 23615 16544 23664 16572
rect 23615 16541 23627 16544
rect 23569 16535 23627 16541
rect 23658 16532 23664 16544
rect 23716 16532 23722 16584
rect 23934 16532 23940 16584
rect 23992 16532 23998 16584
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16572 24639 16575
rect 24670 16572 24676 16584
rect 24627 16544 24676 16572
rect 24627 16541 24639 16544
rect 24581 16535 24639 16541
rect 24670 16532 24676 16544
rect 24728 16532 24734 16584
rect 24964 16581 24992 16680
rect 25590 16600 25596 16652
rect 25648 16600 25654 16652
rect 26160 16640 26188 16680
rect 26418 16668 26424 16720
rect 26476 16708 26482 16720
rect 26476 16680 28212 16708
rect 26476 16668 26482 16680
rect 26160 16612 27476 16640
rect 24857 16575 24915 16581
rect 24857 16541 24869 16575
rect 24903 16541 24915 16575
rect 24857 16535 24915 16541
rect 24949 16575 25007 16581
rect 24949 16541 24961 16575
rect 24995 16541 25007 16575
rect 24949 16535 25007 16541
rect 23750 16464 23756 16516
rect 23808 16504 23814 16516
rect 24872 16504 24900 16535
rect 25498 16532 25504 16584
rect 25556 16532 25562 16584
rect 25608 16572 25636 16600
rect 26160 16584 26188 16612
rect 25685 16575 25743 16581
rect 25685 16572 25697 16575
rect 25608 16544 25697 16572
rect 25685 16541 25697 16544
rect 25731 16541 25743 16575
rect 25685 16535 25743 16541
rect 26142 16532 26148 16584
rect 26200 16572 26206 16584
rect 27448 16581 27476 16612
rect 27982 16600 27988 16652
rect 28040 16600 28046 16652
rect 26329 16575 26387 16581
rect 26329 16572 26341 16575
rect 26200 16544 26341 16572
rect 26200 16532 26206 16544
rect 26329 16541 26341 16544
rect 26375 16541 26387 16575
rect 26605 16575 26663 16581
rect 26605 16574 26617 16575
rect 26528 16572 26617 16574
rect 26329 16535 26387 16541
rect 26436 16546 26617 16572
rect 26436 16544 26556 16546
rect 25041 16507 25099 16513
rect 25041 16504 25053 16507
rect 23808 16476 25053 16504
rect 23808 16464 23814 16476
rect 25041 16473 25053 16476
rect 25087 16473 25099 16507
rect 25041 16467 25099 16473
rect 25593 16507 25651 16513
rect 25593 16473 25605 16507
rect 25639 16504 25651 16507
rect 26436 16504 26464 16544
rect 26605 16541 26617 16546
rect 26651 16541 26663 16575
rect 26605 16535 26663 16541
rect 27433 16575 27491 16581
rect 27433 16541 27445 16575
rect 27479 16541 27491 16575
rect 27433 16535 27491 16541
rect 25639 16476 26464 16504
rect 25639 16473 25651 16476
rect 25593 16467 25651 16473
rect 26694 16464 26700 16516
rect 26752 16464 26758 16516
rect 26881 16507 26939 16513
rect 26881 16473 26893 16507
rect 26927 16473 26939 16507
rect 27448 16504 27476 16535
rect 27614 16532 27620 16584
rect 27672 16532 27678 16584
rect 27709 16575 27767 16581
rect 27709 16541 27721 16575
rect 27755 16572 27767 16575
rect 27890 16572 27896 16584
rect 27755 16544 27896 16572
rect 27755 16541 27767 16544
rect 27709 16535 27767 16541
rect 27890 16532 27896 16544
rect 27948 16532 27954 16584
rect 28000 16572 28028 16600
rect 28184 16591 28212 16680
rect 28169 16585 28227 16591
rect 28073 16572 28131 16575
rect 28000 16569 28131 16572
rect 28000 16544 28085 16569
rect 28073 16535 28085 16544
rect 28119 16535 28131 16569
rect 28169 16551 28181 16585
rect 28215 16551 28227 16585
rect 28169 16545 28227 16551
rect 28073 16529 28131 16535
rect 28350 16532 28356 16584
rect 28408 16581 28414 16584
rect 28408 16572 28419 16581
rect 28408 16544 28453 16572
rect 28408 16535 28419 16544
rect 28408 16532 28414 16535
rect 28626 16532 28632 16584
rect 28684 16532 28690 16584
rect 27801 16507 27859 16513
rect 27801 16504 27813 16507
rect 27448 16476 27813 16504
rect 26881 16467 26939 16473
rect 27801 16473 27813 16476
rect 27847 16473 27859 16507
rect 27801 16467 27859 16473
rect 24765 16439 24823 16445
rect 24765 16436 24777 16439
rect 23308 16408 24777 16436
rect 24765 16405 24777 16408
rect 24811 16436 24823 16439
rect 26050 16436 26056 16448
rect 24811 16408 26056 16436
rect 24811 16405 24823 16408
rect 24765 16399 24823 16405
rect 26050 16396 26056 16408
rect 26108 16396 26114 16448
rect 26418 16396 26424 16448
rect 26476 16436 26482 16448
rect 26513 16439 26571 16445
rect 26513 16436 26525 16439
rect 26476 16408 26525 16436
rect 26476 16396 26482 16408
rect 26513 16405 26525 16408
rect 26559 16405 26571 16439
rect 26513 16399 26571 16405
rect 26602 16396 26608 16448
rect 26660 16436 26666 16448
rect 26896 16436 26924 16467
rect 26660 16408 26924 16436
rect 26660 16396 26666 16408
rect 27246 16396 27252 16448
rect 27304 16396 27310 16448
rect 27982 16396 27988 16448
rect 28040 16436 28046 16448
rect 28644 16436 28672 16532
rect 28040 16408 28672 16436
rect 28040 16396 28046 16408
rect 1104 16346 29595 16368
rect 1104 16294 8032 16346
rect 8084 16294 8096 16346
rect 8148 16294 8160 16346
rect 8212 16294 8224 16346
rect 8276 16294 8288 16346
rect 8340 16294 15115 16346
rect 15167 16294 15179 16346
rect 15231 16294 15243 16346
rect 15295 16294 15307 16346
rect 15359 16294 15371 16346
rect 15423 16294 22198 16346
rect 22250 16294 22262 16346
rect 22314 16294 22326 16346
rect 22378 16294 22390 16346
rect 22442 16294 22454 16346
rect 22506 16294 29281 16346
rect 29333 16294 29345 16346
rect 29397 16294 29409 16346
rect 29461 16294 29473 16346
rect 29525 16294 29537 16346
rect 29589 16294 29595 16346
rect 1104 16272 29595 16294
rect 1397 16235 1455 16241
rect 1397 16201 1409 16235
rect 1443 16232 1455 16235
rect 1670 16232 1676 16244
rect 1443 16204 1676 16232
rect 1443 16201 1455 16204
rect 1397 16195 1455 16201
rect 1670 16192 1676 16204
rect 1728 16192 1734 16244
rect 4430 16232 4436 16244
rect 2792 16204 4436 16232
rect 2792 16173 2820 16204
rect 4430 16192 4436 16204
rect 4488 16192 4494 16244
rect 4982 16192 4988 16244
rect 5040 16192 5046 16244
rect 5442 16192 5448 16244
rect 5500 16232 5506 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 5500 16204 6193 16232
rect 5500 16192 5506 16204
rect 6181 16201 6193 16204
rect 6227 16201 6239 16235
rect 6181 16195 6239 16201
rect 6270 16192 6276 16244
rect 6328 16232 6334 16244
rect 6328 16204 6868 16232
rect 6328 16192 6334 16204
rect 2777 16167 2835 16173
rect 2777 16133 2789 16167
rect 2823 16133 2835 16167
rect 2777 16127 2835 16133
rect 5736 16136 6500 16164
rect 5736 16108 5764 16136
rect 934 16056 940 16108
rect 992 16096 998 16108
rect 1581 16099 1639 16105
rect 1581 16096 1593 16099
rect 992 16068 1593 16096
rect 992 16056 998 16068
rect 1581 16065 1593 16068
rect 1627 16065 1639 16099
rect 1581 16059 1639 16065
rect 3878 16056 3884 16108
rect 3936 16096 3942 16108
rect 5442 16096 5448 16108
rect 3936 16068 5448 16096
rect 3936 16056 3942 16068
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 5537 16099 5595 16105
rect 5537 16065 5549 16099
rect 5583 16096 5595 16099
rect 5626 16096 5632 16108
rect 5583 16068 5632 16096
rect 5583 16065 5595 16068
rect 5537 16059 5595 16065
rect 5626 16056 5632 16068
rect 5684 16056 5690 16108
rect 5718 16056 5724 16108
rect 5776 16056 5782 16108
rect 6178 16056 6184 16108
rect 6236 16096 6242 16108
rect 6472 16105 6500 16136
rect 6546 16124 6552 16176
rect 6604 16164 6610 16176
rect 6641 16167 6699 16173
rect 6641 16164 6653 16167
rect 6604 16136 6653 16164
rect 6604 16124 6610 16136
rect 6641 16133 6653 16136
rect 6687 16133 6699 16167
rect 6641 16127 6699 16133
rect 6840 16105 6868 16204
rect 7558 16192 7564 16244
rect 7616 16232 7622 16244
rect 7653 16235 7711 16241
rect 7653 16232 7665 16235
rect 7616 16204 7665 16232
rect 7616 16192 7622 16204
rect 7653 16201 7665 16204
rect 7699 16201 7711 16235
rect 7653 16195 7711 16201
rect 7760 16204 12296 16232
rect 7760 16176 7788 16204
rect 6914 16124 6920 16176
rect 6972 16164 6978 16176
rect 7285 16167 7343 16173
rect 7285 16164 7297 16167
rect 6972 16136 7297 16164
rect 6972 16124 6978 16136
rect 7285 16133 7297 16136
rect 7331 16133 7343 16167
rect 7285 16127 7343 16133
rect 7377 16167 7435 16173
rect 7377 16133 7389 16167
rect 7423 16164 7435 16167
rect 7742 16164 7748 16176
rect 7423 16136 7748 16164
rect 7423 16133 7435 16136
rect 7377 16127 7435 16133
rect 7742 16124 7748 16136
rect 7800 16124 7806 16176
rect 9309 16167 9367 16173
rect 9309 16164 9321 16167
rect 8036 16136 9321 16164
rect 6365 16099 6423 16105
rect 6365 16096 6377 16099
rect 6236 16068 6377 16096
rect 6236 16056 6242 16068
rect 6365 16065 6377 16068
rect 6411 16065 6423 16099
rect 6365 16059 6423 16065
rect 6458 16099 6516 16105
rect 6458 16065 6470 16099
rect 6504 16065 6516 16099
rect 6458 16059 6516 16065
rect 6733 16099 6791 16105
rect 6733 16065 6745 16099
rect 6779 16065 6791 16099
rect 6733 16059 6791 16065
rect 6830 16099 6888 16105
rect 6830 16065 6842 16099
rect 6876 16065 6888 16099
rect 6830 16059 6888 16065
rect 7101 16099 7159 16105
rect 7101 16065 7113 16099
rect 7147 16096 7159 16099
rect 7147 16068 7328 16096
rect 7147 16065 7159 16068
rect 7101 16059 7159 16065
rect 1394 15988 1400 16040
rect 1452 16028 1458 16040
rect 2501 16031 2559 16037
rect 2501 16028 2513 16031
rect 1452 16000 2513 16028
rect 1452 15988 1458 16000
rect 2501 15997 2513 16000
rect 2547 15997 2559 16031
rect 2501 15991 2559 15997
rect 4433 16031 4491 16037
rect 4433 15997 4445 16031
rect 4479 15997 4491 16031
rect 4433 15991 4491 15997
rect 4338 15920 4344 15972
rect 4396 15960 4402 15972
rect 4448 15960 4476 15991
rect 6748 15960 6776 16059
rect 7300 16028 7328 16068
rect 7466 16056 7472 16108
rect 7524 16056 7530 16108
rect 7926 16056 7932 16108
rect 7984 16056 7990 16108
rect 8036 16028 8064 16136
rect 9309 16133 9321 16136
rect 9355 16133 9367 16167
rect 12161 16167 12219 16173
rect 12161 16164 12173 16167
rect 9309 16127 9367 16133
rect 9876 16136 12173 16164
rect 9876 16105 9904 16136
rect 12161 16133 12173 16136
rect 12207 16133 12219 16167
rect 12268 16164 12296 16204
rect 22830 16192 22836 16244
rect 22888 16232 22894 16244
rect 22888 16204 24854 16232
rect 22888 16192 22894 16204
rect 12268 16136 12388 16164
rect 12161 16127 12219 16133
rect 9861 16099 9919 16105
rect 9861 16065 9873 16099
rect 9907 16065 9919 16099
rect 9861 16059 9919 16065
rect 10042 16056 10048 16108
rect 10100 16056 10106 16108
rect 10134 16056 10140 16108
rect 10192 16056 10198 16108
rect 10229 16099 10287 16105
rect 10229 16065 10241 16099
rect 10275 16096 10287 16099
rect 10318 16096 10324 16108
rect 10275 16068 10324 16096
rect 10275 16065 10287 16068
rect 10229 16059 10287 16065
rect 10318 16056 10324 16068
rect 10376 16056 10382 16108
rect 7300 16000 8064 16028
rect 8202 15988 8208 16040
rect 8260 15988 8266 16040
rect 8662 15988 8668 16040
rect 8720 15988 8726 16040
rect 10502 16028 10508 16040
rect 9048 16000 10508 16028
rect 4396 15932 6776 15960
rect 7009 15963 7067 15969
rect 4396 15920 4402 15932
rect 7009 15929 7021 15963
rect 7055 15960 7067 15963
rect 8386 15960 8392 15972
rect 7055 15932 8392 15960
rect 7055 15929 7067 15932
rect 7009 15923 7067 15929
rect 8386 15920 8392 15932
rect 8444 15920 8450 15972
rect 4249 15895 4307 15901
rect 4249 15861 4261 15895
rect 4295 15892 4307 15895
rect 9048 15892 9076 16000
rect 10502 15988 10508 16000
rect 10560 15988 10566 16040
rect 11054 15988 11060 16040
rect 11112 16028 11118 16040
rect 11517 16031 11575 16037
rect 11517 16028 11529 16031
rect 11112 16000 11529 16028
rect 11112 15988 11118 16000
rect 11517 15997 11529 16000
rect 11563 15997 11575 16031
rect 12360 16028 12388 16136
rect 12894 16124 12900 16176
rect 12952 16164 12958 16176
rect 13265 16167 13323 16173
rect 12952 16136 13216 16164
rect 12952 16124 12958 16136
rect 13188 16108 13216 16136
rect 13265 16133 13277 16167
rect 13311 16164 13323 16167
rect 16025 16167 16083 16173
rect 16025 16164 16037 16167
rect 13311 16136 13952 16164
rect 13311 16133 13323 16136
rect 13265 16127 13323 16133
rect 13924 16108 13952 16136
rect 14016 16136 16037 16164
rect 12618 16056 12624 16108
rect 12676 16096 12682 16108
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 12676 16068 13001 16096
rect 12676 16056 12682 16068
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 13170 16056 13176 16108
rect 13228 16056 13234 16108
rect 13354 16056 13360 16108
rect 13412 16056 13418 16108
rect 13906 16056 13912 16108
rect 13964 16056 13970 16108
rect 13630 16028 13636 16040
rect 12360 16000 13636 16028
rect 11517 15991 11575 15997
rect 13630 15988 13636 16000
rect 13688 16028 13694 16040
rect 14016 16028 14044 16136
rect 16025 16133 16037 16136
rect 16071 16133 16083 16167
rect 16025 16127 16083 16133
rect 23198 16124 23204 16176
rect 23256 16164 23262 16176
rect 23293 16167 23351 16173
rect 23293 16164 23305 16167
rect 23256 16136 23305 16164
rect 23256 16124 23262 16136
rect 23293 16133 23305 16136
rect 23339 16133 23351 16167
rect 24826 16164 24854 16204
rect 26694 16192 26700 16244
rect 26752 16192 26758 16244
rect 27338 16192 27344 16244
rect 27396 16232 27402 16244
rect 27798 16232 27804 16244
rect 27396 16204 27804 16232
rect 27396 16192 27402 16204
rect 27798 16192 27804 16204
rect 27856 16192 27862 16244
rect 26712 16164 26740 16192
rect 24826 16136 26740 16164
rect 23293 16127 23351 16133
rect 14826 16056 14832 16108
rect 14884 16096 14890 16108
rect 15470 16096 15476 16108
rect 14884 16068 15476 16096
rect 14884 16056 14890 16068
rect 15470 16056 15476 16068
rect 15528 16056 15534 16108
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16096 15715 16099
rect 15749 16099 15807 16105
rect 15749 16096 15761 16099
rect 15703 16068 15761 16096
rect 15703 16065 15715 16068
rect 15657 16059 15715 16065
rect 15749 16065 15761 16068
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 15838 16056 15844 16108
rect 15896 16096 15902 16108
rect 15933 16099 15991 16105
rect 15933 16096 15945 16099
rect 15896 16068 15945 16096
rect 15896 16056 15902 16068
rect 15933 16065 15945 16068
rect 15979 16065 15991 16099
rect 15933 16059 15991 16065
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 16482 16096 16488 16108
rect 16163 16068 16488 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 16482 16056 16488 16068
rect 16540 16056 16546 16108
rect 23477 16099 23535 16105
rect 23477 16065 23489 16099
rect 23523 16096 23535 16099
rect 23934 16096 23940 16108
rect 23523 16068 23940 16096
rect 23523 16065 23535 16068
rect 23477 16059 23535 16065
rect 23934 16056 23940 16068
rect 23992 16056 23998 16108
rect 25700 16105 25728 16136
rect 25685 16099 25743 16105
rect 25685 16065 25697 16099
rect 25731 16065 25743 16099
rect 25685 16059 25743 16065
rect 25869 16099 25927 16105
rect 25869 16065 25881 16099
rect 25915 16096 25927 16099
rect 26602 16096 26608 16108
rect 25915 16068 26608 16096
rect 25915 16065 25927 16068
rect 25869 16059 25927 16065
rect 13688 16000 14044 16028
rect 13688 15988 13694 16000
rect 15010 15988 15016 16040
rect 15068 16028 15074 16040
rect 15105 16031 15163 16037
rect 15105 16028 15117 16031
rect 15068 16000 15117 16028
rect 15068 15988 15074 16000
rect 15105 15997 15117 16000
rect 15151 16028 15163 16031
rect 15151 16000 16160 16028
rect 15151 15997 15163 16000
rect 15105 15991 15163 15997
rect 9858 15920 9864 15972
rect 9916 15960 9922 15972
rect 10134 15960 10140 15972
rect 9916 15932 10140 15960
rect 9916 15920 9922 15932
rect 10134 15920 10140 15932
rect 10192 15920 10198 15972
rect 11164 15932 12296 15960
rect 4295 15864 9076 15892
rect 4295 15861 4307 15864
rect 4249 15855 4307 15861
rect 9950 15852 9956 15904
rect 10008 15892 10014 15904
rect 11164 15901 11192 15932
rect 10413 15895 10471 15901
rect 10413 15892 10425 15895
rect 10008 15864 10425 15892
rect 10008 15852 10014 15864
rect 10413 15861 10425 15864
rect 10459 15861 10471 15895
rect 10413 15855 10471 15861
rect 11149 15895 11207 15901
rect 11149 15861 11161 15895
rect 11195 15861 11207 15895
rect 12268 15892 12296 15932
rect 12342 15920 12348 15972
rect 12400 15960 12406 15972
rect 13078 15960 13084 15972
rect 12400 15932 13084 15960
rect 12400 15920 12406 15932
rect 13078 15920 13084 15932
rect 13136 15920 13142 15972
rect 13464 15932 15976 15960
rect 13464 15892 13492 15932
rect 15948 15904 15976 15932
rect 16132 15904 16160 16000
rect 25498 15988 25504 16040
rect 25556 16028 25562 16040
rect 25884 16028 25912 16059
rect 26602 16056 26608 16068
rect 26660 16056 26666 16108
rect 25556 16000 25912 16028
rect 25556 15988 25562 16000
rect 23382 15920 23388 15972
rect 23440 15960 23446 15972
rect 23658 15960 23664 15972
rect 23440 15932 23664 15960
rect 23440 15920 23446 15932
rect 23658 15920 23664 15932
rect 23716 15960 23722 15972
rect 27356 15960 27384 16192
rect 23716 15932 27384 15960
rect 23716 15920 23722 15932
rect 12268 15864 13492 15892
rect 13541 15895 13599 15901
rect 11149 15855 11207 15861
rect 13541 15861 13553 15895
rect 13587 15892 13599 15895
rect 13814 15892 13820 15904
rect 13587 15864 13820 15892
rect 13587 15861 13599 15864
rect 13541 15855 13599 15861
rect 13814 15852 13820 15864
rect 13872 15852 13878 15904
rect 15470 15852 15476 15904
rect 15528 15892 15534 15904
rect 15746 15892 15752 15904
rect 15528 15864 15752 15892
rect 15528 15852 15534 15864
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 15930 15852 15936 15904
rect 15988 15852 15994 15904
rect 16114 15852 16120 15904
rect 16172 15852 16178 15904
rect 16298 15852 16304 15904
rect 16356 15852 16362 15904
rect 25777 15895 25835 15901
rect 25777 15861 25789 15895
rect 25823 15892 25835 15895
rect 26142 15892 26148 15904
rect 25823 15864 26148 15892
rect 25823 15861 25835 15864
rect 25777 15855 25835 15861
rect 26142 15852 26148 15864
rect 26200 15852 26206 15904
rect 1104 15802 29440 15824
rect 1104 15750 4491 15802
rect 4543 15750 4555 15802
rect 4607 15750 4619 15802
rect 4671 15750 4683 15802
rect 4735 15750 4747 15802
rect 4799 15750 11574 15802
rect 11626 15750 11638 15802
rect 11690 15750 11702 15802
rect 11754 15750 11766 15802
rect 11818 15750 11830 15802
rect 11882 15750 18657 15802
rect 18709 15750 18721 15802
rect 18773 15750 18785 15802
rect 18837 15750 18849 15802
rect 18901 15750 18913 15802
rect 18965 15750 25740 15802
rect 25792 15750 25804 15802
rect 25856 15750 25868 15802
rect 25920 15750 25932 15802
rect 25984 15750 25996 15802
rect 26048 15750 29440 15802
rect 1104 15728 29440 15750
rect 3605 15691 3663 15697
rect 3605 15657 3617 15691
rect 3651 15688 3663 15691
rect 4338 15688 4344 15700
rect 3651 15660 4344 15688
rect 3651 15657 3663 15660
rect 3605 15651 3663 15657
rect 4338 15648 4344 15660
rect 4396 15648 4402 15700
rect 5718 15648 5724 15700
rect 5776 15688 5782 15700
rect 5997 15691 6055 15697
rect 5997 15688 6009 15691
rect 5776 15660 6009 15688
rect 5776 15648 5782 15660
rect 5997 15657 6009 15660
rect 6043 15657 6055 15691
rect 7926 15688 7932 15700
rect 5997 15651 6055 15657
rect 6104 15660 7932 15688
rect 6104 15620 6132 15660
rect 7926 15648 7932 15660
rect 7984 15688 7990 15700
rect 8389 15691 8447 15697
rect 7984 15660 8340 15688
rect 7984 15648 7990 15660
rect 5552 15592 6132 15620
rect 1394 15512 1400 15564
rect 1452 15552 1458 15564
rect 1857 15555 1915 15561
rect 1857 15552 1869 15555
rect 1452 15524 1869 15552
rect 1452 15512 1458 15524
rect 1857 15521 1869 15524
rect 1903 15521 1915 15555
rect 1857 15515 1915 15521
rect 2133 15555 2191 15561
rect 2133 15521 2145 15555
rect 2179 15552 2191 15555
rect 3326 15552 3332 15564
rect 2179 15524 3332 15552
rect 2179 15521 2191 15524
rect 2133 15515 2191 15521
rect 3326 15512 3332 15524
rect 3384 15512 3390 15564
rect 3234 15444 3240 15496
rect 3292 15484 3298 15496
rect 3878 15484 3884 15496
rect 3292 15456 3884 15484
rect 3292 15444 3298 15456
rect 3878 15444 3884 15456
rect 3936 15444 3942 15496
rect 4062 15444 4068 15496
rect 4120 15484 4126 15496
rect 4249 15487 4307 15493
rect 4249 15484 4261 15487
rect 4120 15456 4261 15484
rect 4120 15444 4126 15456
rect 4249 15453 4261 15456
rect 4295 15453 4307 15487
rect 5552 15484 5580 15592
rect 6917 15555 6975 15561
rect 6917 15521 6929 15555
rect 6963 15552 6975 15555
rect 7558 15552 7564 15564
rect 6963 15524 7564 15552
rect 6963 15521 6975 15524
rect 6917 15515 6975 15521
rect 7558 15512 7564 15524
rect 7616 15512 7622 15564
rect 5552 15456 5658 15484
rect 4249 15447 4307 15453
rect 5810 15444 5816 15496
rect 5868 15444 5874 15496
rect 6638 15444 6644 15496
rect 6696 15444 6702 15496
rect 7926 15444 7932 15496
rect 7984 15484 7990 15496
rect 8202 15484 8208 15496
rect 7984 15456 8208 15484
rect 7984 15444 7990 15456
rect 8202 15444 8208 15456
rect 8260 15444 8266 15496
rect 4525 15419 4583 15425
rect 4525 15385 4537 15419
rect 4571 15385 4583 15419
rect 4525 15379 4583 15385
rect 4540 15348 4568 15379
rect 5828 15348 5856 15444
rect 8312 15416 8340 15660
rect 8389 15657 8401 15691
rect 8435 15688 8447 15691
rect 8662 15688 8668 15700
rect 8435 15660 8668 15688
rect 8435 15657 8447 15660
rect 8389 15651 8447 15657
rect 8662 15648 8668 15660
rect 8720 15648 8726 15700
rect 9480 15691 9538 15697
rect 9480 15657 9492 15691
rect 9526 15688 9538 15691
rect 9950 15688 9956 15700
rect 9526 15660 9956 15688
rect 9526 15657 9538 15660
rect 9480 15651 9538 15657
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 10778 15648 10784 15700
rect 10836 15688 10842 15700
rect 10965 15691 11023 15697
rect 10965 15688 10977 15691
rect 10836 15660 10977 15688
rect 10836 15648 10842 15660
rect 10965 15657 10977 15660
rect 11011 15688 11023 15691
rect 11054 15688 11060 15700
rect 11011 15660 11060 15688
rect 11011 15657 11023 15660
rect 10965 15651 11023 15657
rect 11054 15648 11060 15660
rect 11112 15648 11118 15700
rect 11698 15648 11704 15700
rect 11756 15688 11762 15700
rect 12158 15688 12164 15700
rect 11756 15660 12164 15688
rect 11756 15648 11762 15660
rect 12158 15648 12164 15660
rect 12216 15648 12222 15700
rect 16114 15648 16120 15700
rect 16172 15648 16178 15700
rect 16298 15648 16304 15700
rect 16356 15648 16362 15700
rect 16408 15660 17908 15688
rect 13909 15623 13967 15629
rect 13909 15620 13921 15623
rect 11900 15592 13921 15620
rect 10134 15512 10140 15564
rect 10192 15552 10198 15564
rect 10192 15524 10732 15552
rect 10192 15512 10198 15524
rect 9214 15444 9220 15496
rect 9272 15444 9278 15496
rect 10704 15484 10732 15524
rect 11900 15493 11928 15592
rect 13909 15589 13921 15592
rect 13955 15589 13967 15623
rect 13909 15583 13967 15589
rect 12618 15512 12624 15564
rect 12676 15512 12682 15564
rect 13078 15512 13084 15564
rect 13136 15512 13142 15564
rect 14645 15555 14703 15561
rect 14645 15521 14657 15555
rect 14691 15552 14703 15555
rect 16316 15552 16344 15648
rect 14691 15524 16344 15552
rect 14691 15521 14703 15524
rect 14645 15515 14703 15521
rect 11885 15487 11943 15493
rect 10704 15456 11836 15484
rect 11808 15428 11836 15456
rect 11885 15453 11897 15487
rect 11931 15453 11943 15487
rect 12161 15487 12219 15493
rect 12161 15484 12173 15487
rect 11885 15447 11943 15453
rect 11992 15456 12173 15484
rect 9582 15416 9588 15428
rect 8312 15388 9588 15416
rect 9582 15376 9588 15388
rect 9640 15416 9646 15428
rect 9950 15416 9956 15428
rect 9640 15388 9956 15416
rect 9640 15376 9646 15388
rect 9950 15376 9956 15388
rect 10008 15376 10014 15428
rect 11790 15376 11796 15428
rect 11848 15416 11854 15428
rect 11992 15416 12020 15456
rect 12161 15453 12173 15456
rect 12207 15453 12219 15487
rect 12161 15447 12219 15453
rect 12250 15444 12256 15496
rect 12308 15444 12314 15496
rect 12710 15444 12716 15496
rect 12768 15444 12774 15496
rect 11848 15388 12020 15416
rect 12069 15419 12127 15425
rect 11848 15376 11854 15388
rect 12069 15385 12081 15419
rect 12115 15416 12127 15419
rect 12728 15416 12756 15444
rect 12115 15388 12756 15416
rect 13096 15416 13124 15512
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15484 13415 15487
rect 13906 15484 13912 15496
rect 13403 15456 13912 15484
rect 13403 15453 13415 15456
rect 13357 15447 13415 15453
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 14366 15444 14372 15496
rect 14424 15444 14430 15496
rect 15746 15444 15752 15496
rect 15804 15484 15810 15496
rect 16114 15484 16120 15496
rect 15804 15456 16120 15484
rect 15804 15444 15810 15456
rect 16114 15444 16120 15456
rect 16172 15484 16178 15496
rect 16408 15484 16436 15660
rect 16485 15555 16543 15561
rect 16485 15521 16497 15555
rect 16531 15552 16543 15555
rect 17402 15552 17408 15564
rect 16531 15524 17408 15552
rect 16531 15521 16543 15524
rect 16485 15515 16543 15521
rect 17402 15512 17408 15524
rect 17460 15512 17466 15564
rect 16172 15456 16436 15484
rect 17880 15470 17908 15660
rect 23566 15648 23572 15700
rect 23624 15648 23630 15700
rect 26142 15648 26148 15700
rect 26200 15688 26206 15700
rect 26237 15691 26295 15697
rect 26237 15688 26249 15691
rect 26200 15660 26249 15688
rect 26200 15648 26206 15660
rect 26237 15657 26249 15660
rect 26283 15657 26295 15691
rect 26970 15688 26976 15700
rect 26237 15651 26295 15657
rect 26344 15660 26976 15688
rect 18506 15580 18512 15632
rect 18564 15620 18570 15632
rect 18785 15623 18843 15629
rect 18785 15620 18797 15623
rect 18564 15592 18797 15620
rect 18564 15580 18570 15592
rect 18785 15589 18797 15592
rect 18831 15620 18843 15623
rect 19978 15620 19984 15632
rect 18831 15592 19984 15620
rect 18831 15589 18843 15592
rect 18785 15583 18843 15589
rect 19978 15580 19984 15592
rect 20036 15620 20042 15632
rect 23201 15623 23259 15629
rect 20036 15592 20208 15620
rect 20036 15580 20042 15592
rect 17954 15512 17960 15564
rect 18012 15552 18018 15564
rect 18693 15555 18751 15561
rect 18693 15552 18705 15555
rect 18012 15524 18705 15552
rect 18012 15512 18018 15524
rect 18693 15521 18705 15524
rect 18739 15521 18751 15555
rect 18693 15515 18751 15521
rect 19720 15524 20024 15552
rect 16172 15444 16178 15456
rect 18138 15444 18144 15496
rect 18196 15484 18202 15496
rect 19720 15493 19748 15524
rect 19996 15493 20024 15524
rect 20180 15493 20208 15592
rect 23201 15589 23213 15623
rect 23247 15620 23259 15623
rect 23290 15620 23296 15632
rect 23247 15592 23296 15620
rect 23247 15589 23259 15592
rect 23201 15583 23259 15589
rect 23290 15580 23296 15592
rect 23348 15580 23354 15632
rect 23400 15592 24716 15620
rect 22646 15512 22652 15564
rect 22704 15552 22710 15564
rect 23106 15552 23112 15564
rect 22704 15524 23112 15552
rect 22704 15512 22710 15524
rect 23106 15512 23112 15524
rect 23164 15552 23170 15564
rect 23400 15552 23428 15592
rect 24688 15564 24716 15592
rect 23164 15524 23428 15552
rect 23164 15512 23170 15524
rect 18417 15487 18475 15493
rect 18417 15484 18429 15487
rect 18196 15456 18429 15484
rect 18196 15444 18202 15456
rect 18417 15453 18429 15456
rect 18463 15453 18475 15487
rect 18417 15447 18475 15453
rect 19613 15487 19671 15493
rect 19613 15453 19625 15487
rect 19659 15484 19671 15487
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 19659 15456 19717 15484
rect 19659 15453 19671 15456
rect 19613 15447 19671 15453
rect 19705 15453 19717 15456
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 19889 15487 19947 15493
rect 19889 15453 19901 15487
rect 19935 15453 19947 15487
rect 19889 15447 19947 15453
rect 19981 15487 20039 15493
rect 19981 15453 19993 15487
rect 20027 15453 20039 15487
rect 19981 15447 20039 15453
rect 20165 15487 20223 15493
rect 20165 15453 20177 15487
rect 20211 15453 20223 15487
rect 20165 15447 20223 15453
rect 13096 15388 15056 15416
rect 12115 15385 12127 15388
rect 12069 15379 12127 15385
rect 4540 15320 5856 15348
rect 6914 15308 6920 15360
rect 6972 15348 6978 15360
rect 12084 15348 12112 15379
rect 6972 15320 12112 15348
rect 6972 15308 6978 15320
rect 12434 15308 12440 15360
rect 12492 15308 12498 15360
rect 13170 15308 13176 15360
rect 13228 15308 13234 15360
rect 15028 15348 15056 15388
rect 15930 15376 15936 15428
rect 15988 15416 15994 15428
rect 16761 15419 16819 15425
rect 16761 15416 16773 15419
rect 15988 15388 16773 15416
rect 15988 15376 15994 15388
rect 16761 15385 16773 15388
rect 16807 15385 16819 15419
rect 19058 15416 19064 15428
rect 16761 15379 16819 15385
rect 18064 15388 19064 15416
rect 18064 15348 18092 15388
rect 19058 15376 19064 15388
rect 19116 15416 19122 15428
rect 19245 15419 19303 15425
rect 19245 15416 19257 15419
rect 19116 15388 19257 15416
rect 19116 15376 19122 15388
rect 19245 15385 19257 15388
rect 19291 15385 19303 15419
rect 19245 15379 19303 15385
rect 19426 15376 19432 15428
rect 19484 15376 19490 15428
rect 19904 15416 19932 15447
rect 23198 15444 23204 15496
rect 23256 15444 23262 15496
rect 23400 15493 23428 15524
rect 23750 15512 23756 15564
rect 23808 15512 23814 15564
rect 24026 15512 24032 15564
rect 24084 15512 24090 15564
rect 24670 15512 24676 15564
rect 24728 15552 24734 15564
rect 26234 15552 26240 15564
rect 24728 15524 26240 15552
rect 24728 15512 24734 15524
rect 23385 15487 23443 15493
rect 23385 15453 23397 15487
rect 23431 15453 23443 15487
rect 23385 15447 23443 15453
rect 23845 15487 23903 15493
rect 23845 15453 23857 15487
rect 23891 15453 23903 15487
rect 23845 15447 23903 15453
rect 23860 15416 23888 15447
rect 23934 15444 23940 15496
rect 23992 15484 23998 15496
rect 23992 15456 24532 15484
rect 23992 15444 23998 15456
rect 24118 15416 24124 15428
rect 19904 15388 24124 15416
rect 24118 15376 24124 15388
rect 24176 15376 24182 15428
rect 15028 15320 18092 15348
rect 18138 15308 18144 15360
rect 18196 15348 18202 15360
rect 18233 15351 18291 15357
rect 18233 15348 18245 15351
rect 18196 15320 18245 15348
rect 18196 15308 18202 15320
rect 18233 15317 18245 15320
rect 18279 15317 18291 15351
rect 18233 15311 18291 15317
rect 19518 15308 19524 15360
rect 19576 15348 19582 15360
rect 19797 15351 19855 15357
rect 19797 15348 19809 15351
rect 19576 15320 19809 15348
rect 19576 15308 19582 15320
rect 19797 15317 19809 15320
rect 19843 15317 19855 15351
rect 19797 15311 19855 15317
rect 20070 15308 20076 15360
rect 20128 15308 20134 15360
rect 24504 15348 24532 15456
rect 26068 15425 26096 15524
rect 26234 15512 26240 15524
rect 26292 15512 26298 15564
rect 26053 15419 26111 15425
rect 26053 15385 26065 15419
rect 26099 15385 26111 15419
rect 26053 15379 26111 15385
rect 26142 15348 26148 15360
rect 24504 15320 26148 15348
rect 26142 15308 26148 15320
rect 26200 15308 26206 15360
rect 26253 15351 26311 15357
rect 26253 15317 26265 15351
rect 26299 15348 26311 15351
rect 26344 15348 26372 15660
rect 26970 15648 26976 15660
rect 27028 15688 27034 15700
rect 27338 15688 27344 15700
rect 27028 15660 27344 15688
rect 27028 15648 27034 15660
rect 27338 15648 27344 15660
rect 27396 15648 27402 15700
rect 26421 15623 26479 15629
rect 26421 15589 26433 15623
rect 26467 15589 26479 15623
rect 26421 15583 26479 15589
rect 26436 15552 26464 15583
rect 26510 15580 26516 15632
rect 26568 15580 26574 15632
rect 26786 15580 26792 15632
rect 26844 15580 26850 15632
rect 28166 15620 28172 15632
rect 26896 15592 28172 15620
rect 26436 15524 26556 15552
rect 26528 15493 26556 15524
rect 26804 15493 26832 15580
rect 26896 15493 26924 15592
rect 28166 15580 28172 15592
rect 28224 15620 28230 15632
rect 28350 15620 28356 15632
rect 28224 15592 28356 15620
rect 28224 15580 28230 15592
rect 28350 15580 28356 15592
rect 28408 15580 28414 15632
rect 27157 15555 27215 15561
rect 27157 15521 27169 15555
rect 27203 15552 27215 15555
rect 27706 15552 27712 15564
rect 27203 15524 27712 15552
rect 27203 15521 27215 15524
rect 27157 15515 27215 15521
rect 27706 15512 27712 15524
rect 27764 15512 27770 15564
rect 26513 15487 26571 15493
rect 26513 15453 26525 15487
rect 26559 15453 26571 15487
rect 26513 15447 26571 15453
rect 26789 15487 26847 15493
rect 26789 15453 26801 15487
rect 26835 15453 26847 15487
rect 26789 15447 26847 15453
rect 26881 15487 26939 15493
rect 26881 15453 26893 15487
rect 26927 15453 26939 15487
rect 26881 15447 26939 15453
rect 27246 15444 27252 15496
rect 27304 15444 27310 15496
rect 27433 15487 27491 15493
rect 27433 15453 27445 15487
rect 27479 15453 27491 15487
rect 27433 15447 27491 15453
rect 27448 15416 27476 15447
rect 26712 15388 27476 15416
rect 26299 15320 26372 15348
rect 26299 15317 26311 15320
rect 26253 15311 26311 15317
rect 26510 15308 26516 15360
rect 26568 15348 26574 15360
rect 26712 15357 26740 15388
rect 26697 15351 26755 15357
rect 26697 15348 26709 15351
rect 26568 15320 26709 15348
rect 26568 15308 26574 15320
rect 26697 15317 26709 15320
rect 26743 15317 26755 15351
rect 26697 15311 26755 15317
rect 27154 15308 27160 15360
rect 27212 15308 27218 15360
rect 27246 15308 27252 15360
rect 27304 15348 27310 15360
rect 27341 15351 27399 15357
rect 27341 15348 27353 15351
rect 27304 15320 27353 15348
rect 27304 15308 27310 15320
rect 27341 15317 27353 15320
rect 27387 15317 27399 15351
rect 27341 15311 27399 15317
rect 1104 15258 29595 15280
rect 1104 15206 8032 15258
rect 8084 15206 8096 15258
rect 8148 15206 8160 15258
rect 8212 15206 8224 15258
rect 8276 15206 8288 15258
rect 8340 15206 15115 15258
rect 15167 15206 15179 15258
rect 15231 15206 15243 15258
rect 15295 15206 15307 15258
rect 15359 15206 15371 15258
rect 15423 15206 22198 15258
rect 22250 15206 22262 15258
rect 22314 15206 22326 15258
rect 22378 15206 22390 15258
rect 22442 15206 22454 15258
rect 22506 15206 29281 15258
rect 29333 15206 29345 15258
rect 29397 15206 29409 15258
rect 29461 15206 29473 15258
rect 29525 15206 29537 15258
rect 29589 15206 29595 15258
rect 1104 15184 29595 15206
rect 5718 15104 5724 15156
rect 5776 15144 5782 15156
rect 5813 15147 5871 15153
rect 5813 15144 5825 15147
rect 5776 15116 5825 15144
rect 5776 15104 5782 15116
rect 5813 15113 5825 15116
rect 5859 15113 5871 15147
rect 5813 15107 5871 15113
rect 6638 15104 6644 15156
rect 6696 15104 6702 15156
rect 7466 15104 7472 15156
rect 7524 15144 7530 15156
rect 7524 15116 8340 15144
rect 7524 15104 7530 15116
rect 6656 15076 6684 15104
rect 6564 15048 6684 15076
rect 8312 15076 8340 15116
rect 8662 15104 8668 15156
rect 8720 15104 8726 15156
rect 9398 15104 9404 15156
rect 9456 15104 9462 15156
rect 10410 15144 10416 15156
rect 9508 15116 10416 15144
rect 8680 15076 8708 15104
rect 8757 15079 8815 15085
rect 8757 15076 8769 15079
rect 8312 15048 8616 15076
rect 8680 15048 8769 15076
rect 5442 14968 5448 15020
rect 5500 15008 5506 15020
rect 6564 15017 6592 15048
rect 8588 15020 8616 15048
rect 8757 15045 8769 15048
rect 8803 15045 8815 15079
rect 9416 15076 9444 15104
rect 9508 15085 9536 15116
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 10962 15104 10968 15156
rect 11020 15104 11026 15156
rect 13170 15144 13176 15156
rect 11624 15116 13176 15144
rect 8757 15039 8815 15045
rect 9232 15048 9444 15076
rect 9493 15079 9551 15085
rect 6549 15011 6607 15017
rect 5500 14980 5672 15008
rect 5500 14968 5506 14980
rect 1394 14900 1400 14952
rect 1452 14940 1458 14952
rect 4062 14940 4068 14952
rect 1452 14912 4068 14940
rect 1452 14900 1458 14912
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 4341 14943 4399 14949
rect 4341 14909 4353 14943
rect 4387 14940 4399 14943
rect 5534 14940 5540 14952
rect 4387 14912 5540 14940
rect 4387 14909 4399 14912
rect 4341 14903 4399 14909
rect 5534 14900 5540 14912
rect 5592 14900 5598 14952
rect 5644 14804 5672 14980
rect 6549 14977 6561 15011
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 7926 14968 7932 15020
rect 7984 14968 7990 15020
rect 8386 14968 8392 15020
rect 8444 14968 8450 15020
rect 8482 15011 8540 15017
rect 8482 14977 8494 15011
rect 8528 14977 8540 15011
rect 8482 14971 8540 14977
rect 6822 14900 6828 14952
rect 6880 14900 6886 14952
rect 7944 14804 7972 14968
rect 8496 14940 8524 14971
rect 8570 14968 8576 15020
rect 8628 15008 8634 15020
rect 8665 15011 8723 15017
rect 8665 15008 8677 15011
rect 8628 14980 8677 15008
rect 8628 14968 8634 14980
rect 8665 14977 8677 14980
rect 8711 14977 8723 15011
rect 8665 14971 8723 14977
rect 8895 15011 8953 15017
rect 8895 14977 8907 15011
rect 8941 15008 8953 15011
rect 9232 15008 9260 15048
rect 9493 15045 9505 15079
rect 9539 15045 9551 15079
rect 9493 15039 9551 15045
rect 9950 15036 9956 15088
rect 10008 15036 10014 15088
rect 11422 15008 11428 15020
rect 8941 14980 9260 15008
rect 10704 14980 11428 15008
rect 8941 14977 8953 14980
rect 8895 14971 8953 14977
rect 8312 14912 8524 14940
rect 5644 14776 7972 14804
rect 8110 14764 8116 14816
rect 8168 14804 8174 14816
rect 8312 14813 8340 14912
rect 9214 14900 9220 14952
rect 9272 14900 9278 14952
rect 10502 14900 10508 14952
rect 10560 14940 10566 14952
rect 10704 14940 10732 14980
rect 11422 14968 11428 14980
rect 11480 14968 11486 15020
rect 11517 15011 11575 15017
rect 11517 14977 11529 15011
rect 11563 15008 11575 15011
rect 11624 15008 11652 15116
rect 13170 15104 13176 15116
rect 13228 15104 13234 15156
rect 13906 15104 13912 15156
rect 13964 15104 13970 15156
rect 15654 15144 15660 15156
rect 14016 15116 15660 15144
rect 11698 15036 11704 15088
rect 11756 15036 11762 15088
rect 11790 15036 11796 15088
rect 11848 15036 11854 15088
rect 12342 15076 12348 15088
rect 11924 15048 12348 15076
rect 11924 15017 11952 15048
rect 12342 15036 12348 15048
rect 12400 15036 12406 15088
rect 12434 15036 12440 15088
rect 12492 15036 12498 15088
rect 11563 14980 11652 15008
rect 11909 15011 11967 15017
rect 11563 14977 11575 14980
rect 11517 14971 11575 14977
rect 11909 14977 11921 15011
rect 11955 14977 11967 15011
rect 11909 14971 11967 14977
rect 13446 14968 13452 15020
rect 13504 15008 13510 15020
rect 13504 14980 13570 15008
rect 13504 14968 13510 14980
rect 10560 14912 10732 14940
rect 10560 14900 10566 14912
rect 11330 14900 11336 14952
rect 11388 14940 11394 14952
rect 12161 14943 12219 14949
rect 12161 14940 12173 14943
rect 11388 14912 12173 14940
rect 11388 14900 11394 14912
rect 12161 14909 12173 14912
rect 12207 14909 12219 14943
rect 14016 14940 14044 15116
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 16206 15104 16212 15156
rect 16264 15104 16270 15156
rect 20806 15144 20812 15156
rect 18248 15116 20812 15144
rect 15746 15036 15752 15088
rect 15804 15036 15810 15088
rect 16224 15008 16252 15104
rect 16390 15036 16396 15088
rect 16448 15076 16454 15088
rect 18248 15085 18276 15116
rect 20806 15104 20812 15116
rect 20864 15104 20870 15156
rect 24762 15104 24768 15156
rect 24820 15144 24826 15156
rect 24854 15144 24860 15156
rect 24820 15116 24860 15144
rect 24820 15104 24826 15116
rect 24854 15104 24860 15116
rect 24912 15144 24918 15156
rect 24912 15116 26556 15144
rect 24912 15104 24918 15116
rect 16669 15079 16727 15085
rect 16669 15076 16681 15079
rect 16448 15048 16681 15076
rect 16448 15036 16454 15048
rect 16669 15045 16681 15048
rect 16715 15076 16727 15079
rect 18233 15079 18291 15085
rect 18233 15076 18245 15079
rect 16715 15048 18245 15076
rect 16715 15045 16727 15048
rect 16669 15039 16727 15045
rect 18233 15045 18245 15048
rect 18279 15045 18291 15079
rect 18233 15039 18291 15045
rect 19061 15079 19119 15085
rect 19061 15045 19073 15079
rect 19107 15076 19119 15079
rect 19334 15076 19340 15088
rect 19107 15048 19340 15076
rect 19107 15045 19119 15048
rect 19061 15039 19119 15045
rect 19334 15036 19340 15048
rect 19392 15076 19398 15088
rect 19392 15048 19932 15076
rect 19392 15036 19398 15048
rect 16301 15011 16359 15017
rect 16301 15008 16313 15011
rect 16224 14980 16313 15008
rect 16301 14977 16313 14980
rect 16347 14977 16359 15011
rect 16301 14971 16359 14977
rect 17681 15011 17739 15017
rect 17681 14977 17693 15011
rect 17727 15008 17739 15011
rect 18138 15008 18144 15020
rect 17727 14980 18144 15008
rect 17727 14977 17739 14980
rect 17681 14971 17739 14977
rect 18138 14968 18144 14980
rect 18196 14968 18202 15020
rect 19429 15011 19487 15017
rect 19429 14977 19441 15011
rect 19475 15008 19487 15011
rect 19518 15008 19524 15020
rect 19475 14980 19524 15008
rect 19475 14977 19487 14980
rect 19429 14971 19487 14977
rect 19518 14968 19524 14980
rect 19576 14968 19582 15020
rect 19613 15011 19671 15017
rect 19613 14977 19625 15011
rect 19659 14977 19671 15011
rect 19613 14971 19671 14977
rect 12161 14903 12219 14909
rect 12268 14912 14044 14940
rect 9033 14875 9091 14881
rect 9033 14841 9045 14875
rect 9079 14841 9091 14875
rect 9033 14835 9091 14841
rect 8297 14807 8355 14813
rect 8297 14804 8309 14807
rect 8168 14776 8309 14804
rect 8168 14764 8174 14776
rect 8297 14773 8309 14776
rect 8343 14773 8355 14807
rect 9048 14804 9076 14835
rect 11422 14832 11428 14884
rect 11480 14872 11486 14884
rect 12069 14875 12127 14881
rect 12069 14872 12081 14875
rect 11480 14844 12081 14872
rect 11480 14832 11486 14844
rect 12069 14841 12081 14844
rect 12115 14841 12127 14875
rect 12069 14835 12127 14841
rect 12268 14804 12296 14912
rect 14366 14900 14372 14952
rect 14424 14940 14430 14952
rect 14461 14943 14519 14949
rect 14461 14940 14473 14943
rect 14424 14912 14473 14940
rect 14424 14900 14430 14912
rect 14461 14909 14473 14912
rect 14507 14909 14519 14943
rect 14461 14903 14519 14909
rect 14737 14943 14795 14949
rect 14737 14909 14749 14943
rect 14783 14940 14795 14943
rect 15470 14940 15476 14952
rect 14783 14912 15476 14940
rect 14783 14909 14795 14912
rect 14737 14903 14795 14909
rect 9048 14776 12296 14804
rect 14476 14804 14504 14903
rect 15470 14900 15476 14912
rect 15528 14900 15534 14952
rect 17402 14900 17408 14952
rect 17460 14900 17466 14952
rect 19628 14940 19656 14971
rect 19702 14968 19708 15020
rect 19760 14968 19766 15020
rect 19904 15017 19932 15048
rect 24026 15036 24032 15088
rect 24084 15076 24090 15088
rect 26528 15085 26556 15116
rect 27154 15104 27160 15156
rect 27212 15104 27218 15156
rect 27338 15104 27344 15156
rect 27396 15104 27402 15156
rect 27586 15116 28028 15144
rect 24995 15079 25053 15085
rect 24995 15076 25007 15079
rect 24084 15048 25007 15076
rect 24084 15036 24090 15048
rect 24995 15045 25007 15048
rect 25041 15076 25053 15079
rect 26513 15079 26571 15085
rect 25041 15048 26464 15076
rect 25041 15045 25053 15048
rect 24995 15039 25053 15045
rect 19889 15011 19947 15017
rect 19889 14977 19901 15011
rect 19935 14977 19947 15011
rect 21450 15008 21456 15020
rect 21298 14980 21456 15008
rect 19889 14971 19947 14977
rect 21450 14968 21456 14980
rect 21508 14968 21514 15020
rect 22097 15011 22155 15017
rect 22097 14977 22109 15011
rect 22143 14977 22155 15011
rect 22097 14971 22155 14977
rect 19794 14940 19800 14952
rect 19352 14912 19800 14940
rect 19352 14884 19380 14912
rect 19794 14900 19800 14912
rect 19852 14900 19858 14952
rect 20162 14900 20168 14952
rect 20220 14900 20226 14952
rect 21637 14943 21695 14949
rect 21637 14909 21649 14943
rect 21683 14940 21695 14943
rect 22112 14940 22140 14971
rect 22922 14968 22928 15020
rect 22980 14968 22986 15020
rect 23290 14968 23296 15020
rect 23348 14968 23354 15020
rect 23382 14968 23388 15020
rect 23440 15008 23446 15020
rect 23753 15011 23811 15017
rect 23753 15008 23765 15011
rect 23440 14980 23765 15008
rect 23440 14968 23446 14980
rect 23753 14977 23765 14980
rect 23799 14977 23811 15011
rect 23753 14971 23811 14977
rect 24670 14968 24676 15020
rect 24728 14968 24734 15020
rect 24762 14968 24768 15020
rect 24820 14968 24826 15020
rect 26436 15017 26464 15048
rect 26513 15045 26525 15079
rect 26559 15076 26571 15079
rect 27172 15076 27200 15104
rect 27249 15079 27307 15085
rect 27249 15076 27261 15079
rect 26559 15048 26648 15076
rect 27172 15048 27261 15076
rect 26559 15045 26571 15048
rect 26513 15039 26571 15045
rect 24857 15011 24915 15017
rect 24857 14977 24869 15011
rect 24903 14977 24915 15011
rect 24857 14971 24915 14977
rect 25133 15011 25191 15017
rect 25133 14977 25145 15011
rect 25179 15008 25191 15011
rect 26053 15011 26111 15017
rect 26053 15008 26065 15011
rect 25179 14980 26065 15008
rect 25179 14977 25191 14980
rect 25133 14971 25191 14977
rect 26053 14977 26065 14980
rect 26099 14977 26111 15011
rect 26053 14971 26111 14977
rect 26145 15011 26203 15017
rect 26145 14977 26157 15011
rect 26191 14977 26203 15011
rect 26145 14971 26203 14977
rect 26421 15011 26479 15017
rect 26421 14977 26433 15011
rect 26467 15008 26479 15011
rect 26467 14980 26556 15008
rect 26467 14977 26479 14980
rect 26421 14971 26479 14977
rect 21683 14912 22140 14940
rect 22281 14943 22339 14949
rect 21683 14909 21695 14912
rect 21637 14903 21695 14909
rect 22281 14909 22293 14943
rect 22327 14909 22339 14943
rect 22281 14903 22339 14909
rect 23308 14940 23336 14968
rect 24872 14940 24900 14971
rect 23308 14912 24900 14940
rect 17954 14832 17960 14884
rect 18012 14832 18018 14884
rect 19334 14832 19340 14884
rect 19392 14832 19398 14884
rect 14734 14804 14740 14816
rect 14476 14776 14740 14804
rect 8297 14767 8355 14773
rect 14734 14764 14740 14776
rect 14792 14764 14798 14816
rect 15102 14764 15108 14816
rect 15160 14804 15166 14816
rect 16209 14807 16267 14813
rect 16209 14804 16221 14807
rect 15160 14776 16221 14804
rect 15160 14764 15166 14776
rect 16209 14773 16221 14776
rect 16255 14773 16267 14807
rect 16209 14767 16267 14773
rect 16393 14807 16451 14813
rect 16393 14773 16405 14807
rect 16439 14804 16451 14807
rect 16574 14804 16580 14816
rect 16439 14776 16580 14804
rect 16439 14773 16451 14776
rect 16393 14767 16451 14773
rect 16574 14764 16580 14776
rect 16632 14764 16638 14816
rect 18138 14764 18144 14816
rect 18196 14764 18202 14816
rect 19245 14807 19303 14813
rect 19245 14773 19257 14807
rect 19291 14804 19303 14807
rect 19610 14804 19616 14816
rect 19291 14776 19616 14804
rect 19291 14773 19303 14776
rect 19245 14767 19303 14773
rect 19610 14764 19616 14776
rect 19668 14764 19674 14816
rect 19812 14804 19840 14900
rect 21542 14804 21548 14816
rect 19812 14776 21548 14804
rect 21542 14764 21548 14776
rect 21600 14804 21606 14816
rect 22296 14804 22324 14903
rect 23308 14872 23336 14912
rect 25498 14900 25504 14952
rect 25556 14900 25562 14952
rect 23032 14844 23336 14872
rect 23032 14816 23060 14844
rect 23934 14832 23940 14884
rect 23992 14872 23998 14884
rect 26160 14872 26188 14971
rect 23992 14844 26188 14872
rect 26528 14872 26556 14980
rect 26620 14940 26648 15048
rect 27249 15045 27261 15048
rect 27295 15045 27307 15079
rect 27356 15076 27384 15104
rect 27586 15076 27614 15116
rect 27356 15048 27614 15076
rect 27709 15079 27767 15085
rect 27249 15039 27307 15045
rect 27709 15045 27721 15079
rect 27755 15076 27767 15079
rect 27798 15076 27804 15088
rect 27755 15048 27804 15076
rect 27755 15045 27767 15048
rect 27709 15039 27767 15045
rect 27798 15036 27804 15048
rect 27856 15036 27862 15088
rect 27154 14968 27160 15020
rect 27212 14968 27218 15020
rect 28000 15017 28028 15116
rect 27341 15011 27399 15017
rect 27341 14977 27353 15011
rect 27387 14977 27399 15011
rect 27459 15011 27517 15017
rect 27459 15008 27471 15011
rect 27341 14971 27399 14977
rect 27448 14977 27471 15008
rect 27505 14977 27517 15011
rect 27448 14971 27517 14977
rect 27893 15011 27951 15017
rect 27893 14977 27905 15011
rect 27939 14977 27951 15011
rect 27893 14971 27951 14977
rect 27985 15011 28043 15017
rect 27985 14977 27997 15011
rect 28031 14977 28043 15011
rect 27985 14971 28043 14977
rect 27356 14940 27384 14971
rect 26620 14912 27384 14940
rect 27448 14872 27476 14971
rect 27617 14943 27675 14949
rect 27617 14909 27629 14943
rect 27663 14940 27675 14943
rect 27908 14940 27936 14971
rect 28166 14968 28172 15020
rect 28224 14968 28230 15020
rect 28184 14940 28212 14968
rect 27663 14912 28212 14940
rect 27663 14909 27675 14912
rect 27617 14903 27675 14909
rect 26528 14844 27476 14872
rect 23992 14832 23998 14844
rect 27706 14832 27712 14884
rect 27764 14832 27770 14884
rect 21600 14776 22324 14804
rect 21600 14764 21606 14776
rect 23014 14764 23020 14816
rect 23072 14764 23078 14816
rect 24486 14764 24492 14816
rect 24544 14764 24550 14816
rect 26973 14807 27031 14813
rect 26973 14773 26985 14807
rect 27019 14804 27031 14807
rect 27062 14804 27068 14816
rect 27019 14776 27068 14804
rect 27019 14773 27031 14776
rect 26973 14767 27031 14773
rect 27062 14764 27068 14776
rect 27120 14764 27126 14816
rect 1104 14714 29440 14736
rect 1104 14662 4491 14714
rect 4543 14662 4555 14714
rect 4607 14662 4619 14714
rect 4671 14662 4683 14714
rect 4735 14662 4747 14714
rect 4799 14662 11574 14714
rect 11626 14662 11638 14714
rect 11690 14662 11702 14714
rect 11754 14662 11766 14714
rect 11818 14662 11830 14714
rect 11882 14662 18657 14714
rect 18709 14662 18721 14714
rect 18773 14662 18785 14714
rect 18837 14662 18849 14714
rect 18901 14662 18913 14714
rect 18965 14662 25740 14714
rect 25792 14662 25804 14714
rect 25856 14662 25868 14714
rect 25920 14662 25932 14714
rect 25984 14662 25996 14714
rect 26048 14662 29440 14714
rect 1104 14640 29440 14662
rect 6822 14560 6828 14612
rect 6880 14600 6886 14612
rect 7653 14603 7711 14609
rect 7653 14600 7665 14603
rect 6880 14572 7665 14600
rect 6880 14560 6886 14572
rect 7653 14569 7665 14572
rect 7699 14569 7711 14603
rect 7653 14563 7711 14569
rect 11422 14560 11428 14612
rect 11480 14600 11486 14612
rect 11480 14572 11744 14600
rect 11480 14560 11486 14572
rect 10134 14532 10140 14544
rect 7392 14504 10140 14532
rect 7392 14476 7420 14504
rect 10134 14492 10140 14504
rect 10192 14492 10198 14544
rect 7006 14424 7012 14476
rect 7064 14464 7070 14476
rect 7374 14464 7380 14476
rect 7064 14436 7380 14464
rect 7064 14424 7070 14436
rect 7374 14424 7380 14436
rect 7432 14424 7438 14476
rect 8110 14424 8116 14476
rect 8168 14424 8174 14476
rect 11330 14464 11336 14476
rect 9232 14436 11336 14464
rect 7101 14399 7159 14405
rect 7101 14365 7113 14399
rect 7147 14365 7159 14399
rect 7392 14396 7420 14424
rect 9232 14408 9260 14436
rect 11330 14424 11336 14436
rect 11388 14464 11394 14476
rect 11609 14467 11667 14473
rect 11609 14464 11621 14467
rect 11388 14436 11621 14464
rect 11388 14424 11394 14436
rect 11609 14433 11621 14436
rect 11655 14433 11667 14467
rect 11716 14464 11744 14572
rect 12618 14560 12624 14612
rect 12676 14600 12682 14612
rect 13357 14603 13415 14609
rect 13357 14600 13369 14603
rect 12676 14572 13369 14600
rect 12676 14560 12682 14572
rect 13357 14569 13369 14572
rect 13403 14569 13415 14603
rect 13357 14563 13415 14569
rect 15102 14560 15108 14612
rect 15160 14560 15166 14612
rect 15378 14560 15384 14612
rect 15436 14600 15442 14612
rect 15654 14600 15660 14612
rect 15436 14572 15660 14600
rect 15436 14560 15442 14572
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 16025 14603 16083 14609
rect 16025 14569 16037 14603
rect 16071 14569 16083 14603
rect 16025 14563 16083 14569
rect 11885 14467 11943 14473
rect 11885 14464 11897 14467
rect 11716 14436 11897 14464
rect 11609 14427 11667 14433
rect 11885 14433 11897 14436
rect 11931 14433 11943 14467
rect 13446 14464 13452 14476
rect 11885 14427 11943 14433
rect 13004 14436 13452 14464
rect 13004 14408 13032 14436
rect 13446 14424 13452 14436
rect 13504 14464 13510 14476
rect 15120 14473 15148 14560
rect 16040 14532 16068 14563
rect 16206 14560 16212 14612
rect 16264 14560 16270 14612
rect 18138 14560 18144 14612
rect 18196 14600 18202 14612
rect 18785 14603 18843 14609
rect 18785 14600 18797 14603
rect 18196 14572 18797 14600
rect 18196 14560 18202 14572
rect 18785 14569 18797 14572
rect 18831 14569 18843 14603
rect 18785 14563 18843 14569
rect 19518 14560 19524 14612
rect 19576 14560 19582 14612
rect 19610 14560 19616 14612
rect 19668 14600 19674 14612
rect 20073 14603 20131 14609
rect 20073 14600 20085 14603
rect 19668 14572 20085 14600
rect 19668 14560 19674 14572
rect 20073 14569 20085 14572
rect 20119 14569 20131 14603
rect 20073 14563 20131 14569
rect 20162 14560 20168 14612
rect 20220 14600 20226 14612
rect 20717 14603 20775 14609
rect 20717 14600 20729 14603
rect 20220 14572 20729 14600
rect 20220 14560 20226 14572
rect 20717 14569 20729 14572
rect 20763 14569 20775 14603
rect 20717 14563 20775 14569
rect 23109 14603 23167 14609
rect 23109 14569 23121 14603
rect 23155 14600 23167 14603
rect 23382 14600 23388 14612
rect 23155 14572 23388 14600
rect 23155 14569 23167 14572
rect 23109 14563 23167 14569
rect 23382 14560 23388 14572
rect 23440 14560 23446 14612
rect 23566 14560 23572 14612
rect 23624 14560 23630 14612
rect 24486 14560 24492 14612
rect 24544 14600 24550 14612
rect 24746 14603 24804 14609
rect 24746 14600 24758 14603
rect 24544 14572 24758 14600
rect 24544 14560 24550 14572
rect 24746 14569 24758 14572
rect 24792 14569 24804 14603
rect 24746 14563 24804 14569
rect 26878 14560 26884 14612
rect 26936 14560 26942 14612
rect 19334 14532 19340 14544
rect 16040 14504 19340 14532
rect 19334 14492 19340 14504
rect 19392 14492 19398 14544
rect 19536 14532 19564 14560
rect 19536 14504 19656 14532
rect 14461 14467 14519 14473
rect 14461 14464 14473 14467
rect 13504 14436 14473 14464
rect 13504 14424 13510 14436
rect 14461 14433 14473 14436
rect 14507 14433 14519 14467
rect 14461 14427 14519 14433
rect 15105 14467 15163 14473
rect 15105 14433 15117 14467
rect 15151 14433 15163 14467
rect 15105 14427 15163 14433
rect 15672 14436 16252 14464
rect 7101 14359 7159 14365
rect 7300 14368 7420 14396
rect 7469 14399 7527 14405
rect 7116 14260 7144 14359
rect 7300 14337 7328 14368
rect 7469 14365 7481 14399
rect 7515 14396 7527 14399
rect 7834 14396 7840 14408
rect 7515 14368 7840 14396
rect 7515 14365 7527 14368
rect 7469 14359 7527 14365
rect 7834 14356 7840 14368
rect 7892 14356 7898 14408
rect 9214 14356 9220 14408
rect 9272 14356 9278 14408
rect 10410 14356 10416 14408
rect 10468 14356 10474 14408
rect 10561 14399 10619 14405
rect 10561 14365 10573 14399
rect 10607 14396 10619 14399
rect 10607 14365 10640 14396
rect 10561 14359 10640 14365
rect 7285 14331 7343 14337
rect 7285 14297 7297 14331
rect 7331 14297 7343 14331
rect 7285 14291 7343 14297
rect 7377 14331 7435 14337
rect 7377 14297 7389 14331
rect 7423 14328 7435 14331
rect 7742 14328 7748 14340
rect 7423 14300 7748 14328
rect 7423 14297 7435 14300
rect 7377 14291 7435 14297
rect 7742 14288 7748 14300
rect 7800 14288 7806 14340
rect 8665 14263 8723 14269
rect 8665 14260 8677 14263
rect 7116 14232 8677 14260
rect 8665 14229 8677 14232
rect 8711 14229 8723 14263
rect 10612 14260 10640 14359
rect 10778 14356 10784 14408
rect 10836 14356 10842 14408
rect 10878 14399 10936 14405
rect 10878 14365 10890 14399
rect 10924 14396 10936 14399
rect 11238 14396 11244 14408
rect 10924 14368 11244 14396
rect 10924 14365 10936 14368
rect 10878 14359 10936 14365
rect 11238 14356 11244 14368
rect 11296 14356 11302 14408
rect 12986 14356 12992 14408
rect 13044 14356 13050 14408
rect 14185 14399 14243 14405
rect 14185 14365 14197 14399
rect 14231 14396 14243 14399
rect 14274 14396 14280 14408
rect 14231 14368 14280 14396
rect 14231 14365 14243 14368
rect 14185 14359 14243 14365
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 14642 14356 14648 14408
rect 14700 14396 14706 14408
rect 15672 14396 15700 14436
rect 14700 14368 15700 14396
rect 14700 14356 14706 14368
rect 15746 14356 15752 14408
rect 15804 14356 15810 14408
rect 10686 14288 10692 14340
rect 10744 14328 10750 14340
rect 11146 14328 11152 14340
rect 10744 14300 11152 14328
rect 10744 14288 10750 14300
rect 11146 14288 11152 14300
rect 11204 14288 11210 14340
rect 16224 14328 16252 14436
rect 16298 14424 16304 14476
rect 16356 14464 16362 14476
rect 16393 14467 16451 14473
rect 16393 14464 16405 14467
rect 16356 14436 16405 14464
rect 16356 14424 16362 14436
rect 16393 14433 16405 14436
rect 16439 14433 16451 14467
rect 16393 14427 16451 14433
rect 16574 14356 16580 14408
rect 16632 14396 16638 14408
rect 18509 14399 18567 14405
rect 18509 14396 18521 14399
rect 16632 14368 18521 14396
rect 16632 14356 16638 14368
rect 18509 14365 18521 14368
rect 18555 14365 18567 14399
rect 18509 14359 18567 14365
rect 18598 14356 18604 14408
rect 18656 14356 18662 14408
rect 18877 14399 18935 14405
rect 18877 14365 18889 14399
rect 18923 14396 18935 14399
rect 19058 14396 19064 14408
rect 18923 14368 19064 14396
rect 18923 14365 18935 14368
rect 18877 14359 18935 14365
rect 19058 14356 19064 14368
rect 19116 14356 19122 14408
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14365 19487 14399
rect 19628 14396 19656 14504
rect 19702 14492 19708 14544
rect 19760 14532 19766 14544
rect 19978 14532 19984 14544
rect 19760 14504 19984 14532
rect 19760 14492 19766 14504
rect 19978 14492 19984 14504
rect 20036 14492 20042 14544
rect 20625 14535 20683 14541
rect 20625 14501 20637 14535
rect 20671 14501 20683 14535
rect 22281 14535 22339 14541
rect 22281 14532 22293 14535
rect 20625 14495 20683 14501
rect 22066 14504 22293 14532
rect 19889 14467 19947 14473
rect 19889 14433 19901 14467
rect 19935 14464 19947 14467
rect 19996 14464 20024 14492
rect 19935 14436 20024 14464
rect 19935 14433 19947 14436
rect 19889 14427 19947 14433
rect 19731 14399 19789 14405
rect 19731 14396 19743 14399
rect 19628 14368 19743 14396
rect 19429 14359 19487 14365
rect 19731 14365 19743 14368
rect 19777 14365 19789 14399
rect 19996 14396 20024 14436
rect 20349 14399 20407 14405
rect 19996 14368 20300 14396
rect 19731 14359 19789 14365
rect 17034 14328 17040 14340
rect 16224 14300 17040 14328
rect 17034 14288 17040 14300
rect 17092 14288 17098 14340
rect 10962 14260 10968 14272
rect 10612 14232 10968 14260
rect 8665 14223 8723 14229
rect 10962 14220 10968 14232
rect 11020 14220 11026 14272
rect 11054 14220 11060 14272
rect 11112 14220 11118 14272
rect 14826 14220 14832 14272
rect 14884 14260 14890 14272
rect 15657 14263 15715 14269
rect 15657 14260 15669 14263
rect 14884 14232 15669 14260
rect 14884 14220 14890 14232
rect 15657 14229 15669 14232
rect 15703 14229 15715 14263
rect 15657 14223 15715 14229
rect 16758 14220 16764 14272
rect 16816 14220 16822 14272
rect 18322 14220 18328 14272
rect 18380 14220 18386 14272
rect 19242 14220 19248 14272
rect 19300 14220 19306 14272
rect 19444 14260 19472 14359
rect 19518 14288 19524 14340
rect 19576 14288 19582 14340
rect 19613 14331 19671 14337
rect 19613 14297 19625 14331
rect 19659 14328 19671 14331
rect 19886 14328 19892 14340
rect 19659 14300 19892 14328
rect 19659 14297 19671 14300
rect 19613 14291 19671 14297
rect 19886 14288 19892 14300
rect 19944 14288 19950 14340
rect 19978 14288 19984 14340
rect 20036 14288 20042 14340
rect 20070 14260 20076 14272
rect 19444 14232 20076 14260
rect 20070 14220 20076 14232
rect 20128 14220 20134 14272
rect 20272 14260 20300 14368
rect 20349 14365 20361 14399
rect 20395 14365 20407 14399
rect 20349 14359 20407 14365
rect 20441 14399 20499 14405
rect 20441 14365 20453 14399
rect 20487 14396 20499 14399
rect 20530 14396 20536 14408
rect 20487 14368 20536 14396
rect 20487 14365 20499 14368
rect 20441 14359 20499 14365
rect 20364 14328 20392 14359
rect 20530 14356 20536 14368
rect 20588 14356 20594 14408
rect 20640 14396 20668 14495
rect 22066 14464 22094 14504
rect 22281 14501 22293 14504
rect 22327 14501 22339 14535
rect 22281 14495 22339 14501
rect 22646 14492 22652 14544
rect 22704 14492 22710 14544
rect 22664 14464 22692 14492
rect 21192 14436 22094 14464
rect 22296 14436 22692 14464
rect 22741 14467 22799 14473
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 20640 14368 20913 14396
rect 20901 14365 20913 14368
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 21192 14328 21220 14436
rect 21361 14399 21419 14405
rect 21361 14365 21373 14399
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 20364 14300 21220 14328
rect 21376 14260 21404 14359
rect 21542 14356 21548 14408
rect 21600 14356 21606 14408
rect 21634 14356 21640 14408
rect 21692 14356 21698 14408
rect 21730 14399 21788 14405
rect 21730 14365 21742 14399
rect 21776 14365 21788 14399
rect 21730 14359 21788 14365
rect 22143 14399 22201 14405
rect 22143 14365 22155 14399
rect 22189 14396 22201 14399
rect 22296 14396 22324 14436
rect 22741 14433 22753 14467
rect 22787 14464 22799 14467
rect 22830 14464 22836 14476
rect 22787 14436 22836 14464
rect 22787 14433 22799 14436
rect 22741 14427 22799 14433
rect 22830 14424 22836 14436
rect 22888 14464 22894 14476
rect 23934 14464 23940 14476
rect 22888 14436 23940 14464
rect 22888 14424 22894 14436
rect 23934 14424 23940 14436
rect 23992 14424 23998 14476
rect 24486 14424 24492 14476
rect 24544 14464 24550 14476
rect 26789 14467 26847 14473
rect 26789 14464 26801 14467
rect 24544 14436 26801 14464
rect 24544 14424 24550 14436
rect 26789 14433 26801 14436
rect 26835 14464 26847 14467
rect 26896 14464 26924 14560
rect 28166 14492 28172 14544
rect 28224 14532 28230 14544
rect 28224 14504 28856 14532
rect 28224 14492 28230 14504
rect 26835 14436 26924 14464
rect 26835 14433 26847 14436
rect 26789 14427 26847 14433
rect 27062 14424 27068 14476
rect 27120 14424 27126 14476
rect 28828 14473 28856 14504
rect 28813 14467 28871 14473
rect 28813 14433 28825 14467
rect 28859 14433 28871 14467
rect 28813 14427 28871 14433
rect 22189 14368 22324 14396
rect 22373 14399 22431 14405
rect 22189 14365 22201 14368
rect 22143 14359 22201 14365
rect 22373 14365 22385 14399
rect 22419 14365 22431 14399
rect 22373 14359 22431 14365
rect 21453 14331 21511 14337
rect 21453 14297 21465 14331
rect 21499 14328 21511 14331
rect 21744 14328 21772 14359
rect 21499 14300 21772 14328
rect 21499 14297 21511 14300
rect 21453 14291 21511 14297
rect 21910 14288 21916 14340
rect 21968 14288 21974 14340
rect 22005 14331 22063 14337
rect 22005 14297 22017 14331
rect 22051 14328 22063 14331
rect 22388 14328 22416 14359
rect 22554 14356 22560 14408
rect 22612 14356 22618 14408
rect 22646 14356 22652 14408
rect 22704 14356 22710 14408
rect 22922 14356 22928 14408
rect 22980 14356 22986 14408
rect 23477 14399 23535 14405
rect 23477 14365 23489 14399
rect 23523 14396 23535 14399
rect 23658 14396 23664 14408
rect 23523 14368 23664 14396
rect 23523 14365 23535 14368
rect 23477 14359 23535 14365
rect 23658 14356 23664 14368
rect 23716 14356 23722 14408
rect 25866 14356 25872 14408
rect 25924 14356 25930 14408
rect 23106 14328 23112 14340
rect 22051 14300 22324 14328
rect 22388 14300 23112 14328
rect 22051 14297 22063 14300
rect 22005 14291 22063 14297
rect 20272 14232 21404 14260
rect 22296 14260 22324 14300
rect 23106 14288 23112 14300
rect 23164 14288 23170 14340
rect 26513 14331 26571 14337
rect 26513 14297 26525 14331
rect 26559 14297 26571 14331
rect 26513 14291 26571 14297
rect 23842 14260 23848 14272
rect 22296 14232 23848 14260
rect 23842 14220 23848 14232
rect 23900 14220 23906 14272
rect 23934 14220 23940 14272
rect 23992 14220 23998 14272
rect 25498 14220 25504 14272
rect 25556 14260 25562 14272
rect 26528 14260 26556 14291
rect 28074 14288 28080 14340
rect 28132 14288 28138 14340
rect 25556 14232 26556 14260
rect 25556 14220 25562 14232
rect 1104 14170 29595 14192
rect 1104 14118 8032 14170
rect 8084 14118 8096 14170
rect 8148 14118 8160 14170
rect 8212 14118 8224 14170
rect 8276 14118 8288 14170
rect 8340 14118 15115 14170
rect 15167 14118 15179 14170
rect 15231 14118 15243 14170
rect 15295 14118 15307 14170
rect 15359 14118 15371 14170
rect 15423 14118 22198 14170
rect 22250 14118 22262 14170
rect 22314 14118 22326 14170
rect 22378 14118 22390 14170
rect 22442 14118 22454 14170
rect 22506 14118 29281 14170
rect 29333 14118 29345 14170
rect 29397 14118 29409 14170
rect 29461 14118 29473 14170
rect 29525 14118 29537 14170
rect 29589 14118 29595 14170
rect 1104 14096 29595 14118
rect 6362 14016 6368 14068
rect 6420 14016 6426 14068
rect 7834 14016 7840 14068
rect 7892 14056 7898 14068
rect 7892 14028 11928 14056
rect 7892 14016 7898 14028
rect 3234 13988 3240 14000
rect 3082 13960 3240 13988
rect 3234 13948 3240 13960
rect 3292 13948 3298 14000
rect 3510 13948 3516 14000
rect 3568 13948 3574 14000
rect 11900 13988 11928 14028
rect 11974 14016 11980 14068
rect 12032 14056 12038 14068
rect 12032 14028 15240 14056
rect 12032 14016 12038 14028
rect 12618 13988 12624 14000
rect 9876 13960 10916 13988
rect 11900 13960 12624 13988
rect 1394 13880 1400 13932
rect 1452 13920 1458 13932
rect 1581 13923 1639 13929
rect 1581 13920 1593 13923
rect 1452 13892 1593 13920
rect 1452 13880 1458 13892
rect 1581 13889 1593 13892
rect 1627 13889 1639 13923
rect 3528 13920 3556 13948
rect 3605 13923 3663 13929
rect 3605 13920 3617 13923
rect 3528 13892 3617 13920
rect 1581 13883 1639 13889
rect 3605 13889 3617 13892
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 5718 13880 5724 13932
rect 5776 13920 5782 13932
rect 9876 13929 9904 13960
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 5776 13892 6561 13920
rect 5776 13880 5782 13892
rect 6549 13889 6561 13892
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 6733 13923 6791 13929
rect 6733 13889 6745 13923
rect 6779 13920 6791 13923
rect 9861 13923 9919 13929
rect 6779 13892 7512 13920
rect 6779 13889 6791 13892
rect 6733 13883 6791 13889
rect 7484 13864 7512 13892
rect 9861 13889 9873 13923
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 10042 13880 10048 13932
rect 10100 13880 10106 13932
rect 10137 13923 10195 13929
rect 10137 13889 10149 13923
rect 10183 13889 10195 13923
rect 10137 13883 10195 13889
rect 10229 13923 10287 13929
rect 10229 13889 10241 13923
rect 10275 13920 10287 13923
rect 10318 13920 10324 13932
rect 10275 13892 10324 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 1854 13812 1860 13864
rect 1912 13812 1918 13864
rect 6178 13812 6184 13864
rect 6236 13812 6242 13864
rect 6638 13812 6644 13864
rect 6696 13812 6702 13864
rect 6825 13855 6883 13861
rect 6825 13821 6837 13855
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 6196 13784 6224 13812
rect 6362 13784 6368 13796
rect 6196 13756 6368 13784
rect 6362 13744 6368 13756
rect 6420 13784 6426 13796
rect 6840 13784 6868 13815
rect 7466 13812 7472 13864
rect 7524 13812 7530 13864
rect 9950 13812 9956 13864
rect 10008 13812 10014 13864
rect 10152 13852 10180 13883
rect 10318 13880 10324 13892
rect 10376 13920 10382 13932
rect 10594 13920 10600 13932
rect 10376 13892 10600 13920
rect 10376 13880 10382 13892
rect 10594 13880 10600 13892
rect 10652 13880 10658 13932
rect 10152 13824 10732 13852
rect 7558 13784 7564 13796
rect 6420 13756 7564 13784
rect 6420 13744 6426 13756
rect 7558 13744 7564 13756
rect 7616 13744 7622 13796
rect 9968 13784 9996 13812
rect 10704 13784 10732 13824
rect 10778 13812 10784 13864
rect 10836 13812 10842 13864
rect 10888 13852 10916 13960
rect 12618 13948 12624 13960
rect 12676 13948 12682 14000
rect 13814 13948 13820 14000
rect 13872 13988 13878 14000
rect 15212 13997 15240 14028
rect 18322 14016 18328 14068
rect 18380 14016 18386 14068
rect 19426 14016 19432 14068
rect 19484 14016 19490 14068
rect 19518 14016 19524 14068
rect 19576 14016 19582 14068
rect 19978 14016 19984 14068
rect 20036 14056 20042 14068
rect 20533 14059 20591 14065
rect 20533 14056 20545 14059
rect 20036 14028 20545 14056
rect 20036 14016 20042 14028
rect 20533 14025 20545 14028
rect 20579 14025 20591 14059
rect 20533 14019 20591 14025
rect 20622 14016 20628 14068
rect 20680 14056 20686 14068
rect 21545 14059 21603 14065
rect 21545 14056 21557 14059
rect 20680 14028 21557 14056
rect 20680 14016 20686 14028
rect 21545 14025 21557 14028
rect 21591 14025 21603 14059
rect 22554 14056 22560 14068
rect 21545 14019 21603 14025
rect 22066 14028 22560 14056
rect 15197 13991 15255 13997
rect 13872 13960 14228 13988
rect 13872 13948 13878 13960
rect 11054 13880 11060 13932
rect 11112 13920 11118 13932
rect 14200 13929 14228 13960
rect 15197 13957 15209 13991
rect 15243 13988 15255 13991
rect 15378 13988 15384 14000
rect 15243 13960 15384 13988
rect 15243 13957 15255 13960
rect 15197 13951 15255 13957
rect 15378 13948 15384 13960
rect 15436 13948 15442 14000
rect 18340 13988 18368 14016
rect 15580 13960 16160 13988
rect 18340 13960 18920 13988
rect 14093 13923 14151 13929
rect 14093 13920 14105 13923
rect 11112 13892 14105 13920
rect 11112 13880 11118 13892
rect 14093 13889 14105 13892
rect 14139 13889 14151 13923
rect 14093 13883 14151 13889
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13920 14519 13923
rect 14642 13920 14648 13932
rect 14507 13892 14648 13920
rect 14507 13889 14519 13892
rect 14461 13883 14519 13889
rect 14642 13880 14648 13892
rect 14700 13880 14706 13932
rect 14826 13880 14832 13932
rect 14884 13920 14890 13932
rect 14921 13923 14979 13929
rect 14921 13920 14933 13923
rect 14884 13892 14933 13920
rect 14884 13880 14890 13892
rect 14921 13889 14933 13892
rect 14967 13889 14979 13923
rect 14921 13883 14979 13889
rect 15010 13880 15016 13932
rect 15068 13880 15074 13932
rect 15105 13923 15163 13929
rect 15105 13889 15117 13923
rect 15151 13889 15163 13923
rect 15105 13883 15163 13889
rect 15289 13923 15347 13929
rect 15289 13889 15301 13923
rect 15335 13920 15347 13923
rect 15580 13920 15608 13960
rect 15335 13892 15608 13920
rect 16132 13920 16160 13960
rect 16482 13920 16488 13932
rect 16132 13892 16488 13920
rect 15335 13889 15347 13892
rect 15289 13883 15347 13889
rect 11333 13855 11391 13861
rect 11333 13852 11345 13855
rect 10888 13824 11345 13852
rect 11333 13821 11345 13824
rect 11379 13821 11391 13855
rect 12986 13852 12992 13864
rect 11333 13815 11391 13821
rect 11532 13824 12992 13852
rect 11422 13784 11428 13796
rect 9968 13756 10640 13784
rect 10704 13756 11428 13784
rect 5902 13676 5908 13728
rect 5960 13716 5966 13728
rect 6546 13716 6552 13728
rect 5960 13688 6552 13716
rect 5960 13676 5966 13688
rect 6546 13676 6552 13688
rect 6604 13716 6610 13728
rect 10226 13716 10232 13728
rect 6604 13688 10232 13716
rect 6604 13676 6610 13688
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 10410 13676 10416 13728
rect 10468 13676 10474 13728
rect 10612 13716 10640 13756
rect 11422 13744 11428 13756
rect 11480 13744 11486 13796
rect 11532 13716 11560 13824
rect 12986 13812 12992 13824
rect 13044 13812 13050 13864
rect 13909 13855 13967 13861
rect 13909 13821 13921 13855
rect 13955 13852 13967 13855
rect 14369 13855 14427 13861
rect 13955 13824 14320 13852
rect 13955 13821 13967 13824
rect 13909 13815 13967 13821
rect 12066 13744 12072 13796
rect 12124 13784 12130 13796
rect 14090 13784 14096 13796
rect 12124 13756 14096 13784
rect 12124 13744 12130 13756
rect 14090 13744 14096 13756
rect 14148 13744 14154 13796
rect 10612 13688 11560 13716
rect 14292 13716 14320 13824
rect 14369 13821 14381 13855
rect 14415 13852 14427 13855
rect 15028 13852 15056 13880
rect 14415 13824 15056 13852
rect 15120 13852 15148 13883
rect 16482 13880 16488 13892
rect 16540 13920 16546 13932
rect 18601 13923 18659 13929
rect 16540 13892 17080 13920
rect 16540 13880 16546 13892
rect 15930 13852 15936 13864
rect 15120 13824 15936 13852
rect 14415 13821 14427 13824
rect 14369 13815 14427 13821
rect 15930 13812 15936 13824
rect 15988 13852 15994 13864
rect 16850 13852 16856 13864
rect 15988 13824 16856 13852
rect 15988 13812 15994 13824
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 15470 13744 15476 13796
rect 15528 13744 15534 13796
rect 17052 13784 17080 13892
rect 18601 13889 18613 13923
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 18616 13852 18644 13883
rect 18690 13880 18696 13932
rect 18748 13880 18754 13932
rect 18892 13929 18920 13960
rect 18877 13923 18935 13929
rect 18877 13889 18889 13923
rect 18923 13889 18935 13923
rect 18877 13883 18935 13889
rect 18969 13923 19027 13929
rect 18969 13889 18981 13923
rect 19015 13920 19027 13923
rect 19061 13923 19119 13929
rect 19061 13920 19073 13923
rect 19015 13892 19073 13920
rect 19015 13889 19027 13892
rect 18969 13883 19027 13889
rect 19061 13889 19073 13892
rect 19107 13889 19119 13923
rect 19061 13883 19119 13889
rect 19150 13880 19156 13932
rect 19208 13920 19214 13932
rect 19245 13923 19303 13929
rect 19245 13920 19257 13923
rect 19208 13892 19257 13920
rect 19208 13880 19214 13892
rect 19245 13889 19257 13892
rect 19291 13889 19303 13923
rect 19245 13883 19303 13889
rect 19334 13880 19340 13932
rect 19392 13880 19398 13932
rect 19444 13852 19472 14016
rect 19536 13988 19564 14016
rect 20073 13991 20131 13997
rect 20073 13988 20085 13991
rect 19536 13960 20085 13988
rect 20073 13957 20085 13960
rect 20119 13957 20131 13991
rect 22066 13988 22094 14028
rect 22554 14016 22560 14028
rect 22612 14016 22618 14068
rect 23106 14016 23112 14068
rect 23164 14056 23170 14068
rect 23661 14059 23719 14065
rect 23661 14056 23673 14059
rect 23164 14028 23673 14056
rect 23164 14016 23170 14028
rect 23661 14025 23673 14028
rect 23707 14025 23719 14059
rect 23661 14019 23719 14025
rect 23842 14016 23848 14068
rect 23900 14056 23906 14068
rect 25130 14056 25136 14068
rect 23900 14028 25136 14056
rect 23900 14016 23906 14028
rect 25130 14016 25136 14028
rect 25188 14016 25194 14068
rect 20073 13951 20131 13957
rect 20732 13960 22094 13988
rect 20732 13932 20760 13960
rect 23566 13948 23572 14000
rect 23624 13988 23630 14000
rect 24118 13988 24124 14000
rect 23624 13960 24124 13988
rect 23624 13948 23630 13960
rect 24118 13948 24124 13960
rect 24176 13948 24182 14000
rect 19518 13880 19524 13932
rect 19576 13880 19582 13932
rect 19610 13880 19616 13932
rect 19668 13880 19674 13932
rect 19702 13880 19708 13932
rect 19760 13880 19766 13932
rect 19794 13880 19800 13932
rect 19852 13920 19858 13932
rect 19889 13923 19947 13929
rect 19889 13920 19901 13923
rect 19852 13892 19901 13920
rect 19852 13880 19858 13892
rect 19889 13889 19901 13892
rect 19935 13889 19947 13923
rect 19889 13883 19947 13889
rect 20165 13923 20223 13929
rect 20165 13889 20177 13923
rect 20211 13920 20223 13923
rect 20714 13920 20720 13932
rect 20211 13892 20720 13920
rect 20211 13889 20223 13892
rect 20165 13883 20223 13889
rect 20180 13852 20208 13883
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 20806 13880 20812 13932
rect 20864 13920 20870 13932
rect 22649 13923 22707 13929
rect 22649 13920 22661 13923
rect 20864 13892 22661 13920
rect 20864 13880 20870 13892
rect 22649 13889 22661 13892
rect 22695 13889 22707 13923
rect 22649 13883 22707 13889
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 24486 13920 24492 13932
rect 23532 13892 24492 13920
rect 23532 13880 23538 13892
rect 24486 13880 24492 13892
rect 24544 13880 24550 13932
rect 25866 13880 25872 13932
rect 25924 13880 25930 13932
rect 28169 13923 28227 13929
rect 28169 13889 28181 13923
rect 28215 13920 28227 13923
rect 28442 13920 28448 13932
rect 28215 13892 28448 13920
rect 28215 13889 28227 13892
rect 28169 13883 28227 13889
rect 28442 13880 28448 13892
rect 28500 13880 28506 13932
rect 18616 13824 19472 13852
rect 19536 13824 20208 13852
rect 20257 13855 20315 13861
rect 17126 13784 17132 13796
rect 17052 13756 17132 13784
rect 17126 13744 17132 13756
rect 17184 13744 17190 13796
rect 18138 13744 18144 13796
rect 18196 13784 18202 13796
rect 19536 13784 19564 13824
rect 20257 13821 20269 13855
rect 20303 13821 20315 13855
rect 20257 13815 20315 13821
rect 21085 13855 21143 13861
rect 21085 13821 21097 13855
rect 21131 13852 21143 13855
rect 22186 13852 22192 13864
rect 21131 13824 22192 13852
rect 21131 13821 21143 13824
rect 21085 13815 21143 13821
rect 20272 13784 20300 13815
rect 22186 13812 22192 13824
rect 22244 13812 22250 13864
rect 24029 13855 24087 13861
rect 24029 13821 24041 13855
rect 24075 13821 24087 13855
rect 24029 13815 24087 13821
rect 18196 13756 19564 13784
rect 19628 13756 20300 13784
rect 21453 13787 21511 13793
rect 18196 13744 18202 13756
rect 16758 13716 16764 13728
rect 14292 13688 16764 13716
rect 16758 13676 16764 13688
rect 16816 13676 16822 13728
rect 18414 13676 18420 13728
rect 18472 13676 18478 13728
rect 19334 13676 19340 13728
rect 19392 13716 19398 13728
rect 19628 13716 19656 13756
rect 21453 13753 21465 13787
rect 21499 13753 21511 13787
rect 21453 13747 21511 13753
rect 19392 13688 19656 13716
rect 19392 13676 19398 13688
rect 20162 13676 20168 13728
rect 20220 13716 20226 13728
rect 21468 13716 21496 13747
rect 21726 13716 21732 13728
rect 20220 13688 21732 13716
rect 20220 13676 20226 13688
rect 21726 13676 21732 13688
rect 21784 13676 21790 13728
rect 24044 13716 24072 13815
rect 24118 13812 24124 13864
rect 24176 13812 24182 13864
rect 24305 13855 24363 13861
rect 24305 13821 24317 13855
rect 24351 13852 24363 13855
rect 24765 13855 24823 13861
rect 24765 13852 24777 13855
rect 24351 13824 24777 13852
rect 24351 13821 24363 13824
rect 24305 13815 24363 13821
rect 24765 13821 24777 13824
rect 24811 13821 24823 13855
rect 25884 13852 25912 13880
rect 26326 13852 26332 13864
rect 25884 13824 26332 13852
rect 24765 13815 24823 13821
rect 26326 13812 26332 13824
rect 26384 13852 26390 13864
rect 28074 13852 28080 13864
rect 26384 13824 28080 13852
rect 26384 13812 26390 13824
rect 28074 13812 28080 13824
rect 28132 13852 28138 13864
rect 28353 13855 28411 13861
rect 28353 13852 28365 13855
rect 28132 13824 28365 13852
rect 28132 13812 28138 13824
rect 28353 13821 28365 13824
rect 28399 13821 28411 13855
rect 28353 13815 28411 13821
rect 25314 13716 25320 13728
rect 24044 13688 25320 13716
rect 25314 13676 25320 13688
rect 25372 13676 25378 13728
rect 26234 13676 26240 13728
rect 26292 13676 26298 13728
rect 1104 13626 29440 13648
rect 1104 13574 4491 13626
rect 4543 13574 4555 13626
rect 4607 13574 4619 13626
rect 4671 13574 4683 13626
rect 4735 13574 4747 13626
rect 4799 13574 11574 13626
rect 11626 13574 11638 13626
rect 11690 13574 11702 13626
rect 11754 13574 11766 13626
rect 11818 13574 11830 13626
rect 11882 13574 18657 13626
rect 18709 13574 18721 13626
rect 18773 13574 18785 13626
rect 18837 13574 18849 13626
rect 18901 13574 18913 13626
rect 18965 13574 25740 13626
rect 25792 13574 25804 13626
rect 25856 13574 25868 13626
rect 25920 13574 25932 13626
rect 25984 13574 25996 13626
rect 26048 13574 29440 13626
rect 1104 13552 29440 13574
rect 1854 13472 1860 13524
rect 1912 13512 1918 13524
rect 2225 13515 2283 13521
rect 2225 13512 2237 13515
rect 1912 13484 2237 13512
rect 1912 13472 1918 13484
rect 2225 13481 2237 13484
rect 2271 13481 2283 13515
rect 2225 13475 2283 13481
rect 6273 13515 6331 13521
rect 6273 13481 6285 13515
rect 6319 13512 6331 13515
rect 6638 13512 6644 13524
rect 6319 13484 6644 13512
rect 6319 13481 6331 13484
rect 6273 13475 6331 13481
rect 6638 13472 6644 13484
rect 6696 13472 6702 13524
rect 8481 13515 8539 13521
rect 8481 13481 8493 13515
rect 8527 13512 8539 13515
rect 13262 13512 13268 13524
rect 8527 13484 13268 13512
rect 8527 13481 8539 13484
rect 8481 13475 8539 13481
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 16390 13512 16396 13524
rect 15212 13484 16396 13512
rect 2593 13447 2651 13453
rect 2593 13413 2605 13447
rect 2639 13413 2651 13447
rect 2593 13407 2651 13413
rect 2409 13311 2467 13317
rect 2409 13277 2421 13311
rect 2455 13308 2467 13311
rect 2608 13308 2636 13407
rect 5994 13404 6000 13456
rect 6052 13444 6058 13456
rect 6454 13444 6460 13456
rect 6052 13416 6460 13444
rect 6052 13404 6058 13416
rect 6454 13404 6460 13416
rect 6512 13444 6518 13456
rect 9674 13444 9680 13456
rect 6512 13416 9680 13444
rect 6512 13404 6518 13416
rect 9674 13404 9680 13416
rect 9732 13404 9738 13456
rect 9766 13404 9772 13456
rect 9824 13444 9830 13456
rect 12069 13447 12127 13453
rect 12069 13444 12081 13447
rect 9824 13416 12081 13444
rect 9824 13404 9830 13416
rect 12069 13413 12081 13416
rect 12115 13413 12127 13447
rect 12069 13407 12127 13413
rect 12526 13404 12532 13456
rect 12584 13444 12590 13456
rect 15212 13444 15240 13484
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 18506 13472 18512 13524
rect 18564 13512 18570 13524
rect 18785 13515 18843 13521
rect 18785 13512 18797 13515
rect 18564 13484 18797 13512
rect 18564 13472 18570 13484
rect 18785 13481 18797 13484
rect 18831 13481 18843 13515
rect 18785 13475 18843 13481
rect 12584 13416 15240 13444
rect 15289 13447 15347 13453
rect 12584 13404 12590 13416
rect 15289 13413 15301 13447
rect 15335 13444 15347 13447
rect 15746 13444 15752 13456
rect 15335 13416 15752 13444
rect 15335 13413 15347 13416
rect 15289 13407 15347 13413
rect 15746 13404 15752 13416
rect 15804 13404 15810 13456
rect 15841 13447 15899 13453
rect 15841 13413 15853 13447
rect 15887 13444 15899 13447
rect 17862 13444 17868 13456
rect 15887 13416 17868 13444
rect 15887 13413 15899 13416
rect 15841 13407 15899 13413
rect 17862 13404 17868 13416
rect 17920 13404 17926 13456
rect 18800 13444 18828 13475
rect 19518 13472 19524 13524
rect 19576 13512 19582 13524
rect 20438 13512 20444 13524
rect 19576 13484 20444 13512
rect 19576 13472 19582 13484
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 22922 13472 22928 13524
rect 22980 13512 22986 13524
rect 23293 13515 23351 13521
rect 23293 13512 23305 13515
rect 22980 13484 23305 13512
rect 22980 13472 22986 13484
rect 23293 13481 23305 13484
rect 23339 13481 23351 13515
rect 23293 13475 23351 13481
rect 25314 13472 25320 13524
rect 25372 13512 25378 13524
rect 25777 13515 25835 13521
rect 25777 13512 25789 13515
rect 25372 13484 25789 13512
rect 25372 13472 25378 13484
rect 25777 13481 25789 13484
rect 25823 13481 25835 13515
rect 25777 13475 25835 13481
rect 28994 13472 29000 13524
rect 29052 13472 29058 13524
rect 20254 13444 20260 13456
rect 18800 13416 19380 13444
rect 3237 13379 3295 13385
rect 3237 13345 3249 13379
rect 3283 13376 3295 13379
rect 3510 13376 3516 13388
rect 3283 13348 3516 13376
rect 3283 13345 3295 13348
rect 3237 13339 3295 13345
rect 3510 13336 3516 13348
rect 3568 13336 3574 13388
rect 7282 13376 7288 13388
rect 6196 13348 7288 13376
rect 2455 13280 2636 13308
rect 2961 13311 3019 13317
rect 2455 13277 2467 13280
rect 2409 13271 2467 13277
rect 2961 13277 2973 13311
rect 3007 13308 3019 13311
rect 3050 13308 3056 13320
rect 3007 13280 3056 13308
rect 3007 13277 3019 13280
rect 2961 13271 3019 13277
rect 3050 13268 3056 13280
rect 3108 13308 3114 13320
rect 6196 13317 6224 13348
rect 7282 13336 7288 13348
rect 7340 13376 7346 13388
rect 13354 13376 13360 13388
rect 7340 13348 9168 13376
rect 7340 13336 7346 13348
rect 3421 13311 3479 13317
rect 3421 13308 3433 13311
rect 3108 13280 3433 13308
rect 3108 13268 3114 13280
rect 3421 13277 3433 13280
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 3605 13311 3663 13317
rect 3605 13277 3617 13311
rect 3651 13277 3663 13311
rect 3605 13271 3663 13277
rect 6181 13311 6239 13317
rect 6181 13277 6193 13311
rect 6227 13277 6239 13311
rect 6181 13271 6239 13277
rect 6549 13311 6607 13317
rect 6549 13277 6561 13311
rect 6595 13308 6607 13311
rect 6914 13308 6920 13320
rect 6595 13280 6920 13308
rect 6595 13277 6607 13280
rect 6549 13271 6607 13277
rect 3620 13240 3648 13271
rect 6914 13268 6920 13280
rect 6972 13268 6978 13320
rect 7190 13268 7196 13320
rect 7248 13268 7254 13320
rect 7377 13311 7435 13317
rect 7377 13277 7389 13311
rect 7423 13277 7435 13311
rect 7377 13271 7435 13277
rect 7208 13240 7236 13268
rect 3620 13212 7236 13240
rect 3053 13175 3111 13181
rect 3053 13141 3065 13175
rect 3099 13172 3111 13175
rect 3234 13172 3240 13184
rect 3099 13144 3240 13172
rect 3099 13141 3111 13144
rect 3053 13135 3111 13141
rect 3234 13132 3240 13144
rect 3292 13172 3298 13184
rect 3513 13175 3571 13181
rect 3513 13172 3525 13175
rect 3292 13144 3525 13172
rect 3292 13132 3298 13144
rect 3513 13141 3525 13144
rect 3559 13141 3571 13175
rect 3513 13135 3571 13141
rect 7098 13132 7104 13184
rect 7156 13132 7162 13184
rect 7190 13132 7196 13184
rect 7248 13172 7254 13184
rect 7392 13172 7420 13271
rect 7558 13268 7564 13320
rect 7616 13268 7622 13320
rect 8128 13317 8156 13348
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13308 8447 13311
rect 8570 13308 8576 13320
rect 8435 13280 8576 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 7837 13243 7895 13249
rect 7837 13209 7849 13243
rect 7883 13240 7895 13243
rect 8404 13240 8432 13271
rect 8570 13268 8576 13280
rect 8628 13268 8634 13320
rect 9140 13317 9168 13348
rect 9416 13348 13360 13376
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 7883 13212 8432 13240
rect 7883 13209 7895 13212
rect 7837 13203 7895 13209
rect 7466 13172 7472 13184
rect 7248 13144 7472 13172
rect 7248 13132 7254 13144
rect 7466 13132 7472 13144
rect 7524 13172 7530 13184
rect 8956 13172 8984 13271
rect 9416 13184 9444 13348
rect 13354 13336 13360 13348
rect 13412 13376 13418 13388
rect 13412 13348 14504 13376
rect 13412 13336 13418 13348
rect 9674 13268 9680 13320
rect 9732 13308 9738 13320
rect 10318 13308 10324 13320
rect 9732 13280 10324 13308
rect 9732 13268 9738 13280
rect 10318 13268 10324 13280
rect 10376 13308 10382 13320
rect 10413 13311 10471 13317
rect 10413 13308 10425 13311
rect 10376 13280 10425 13308
rect 10376 13268 10382 13280
rect 10413 13277 10425 13280
rect 10459 13277 10471 13311
rect 10413 13271 10471 13277
rect 10502 13268 10508 13320
rect 10560 13308 10566 13320
rect 10560 13280 10605 13308
rect 10560 13268 10566 13280
rect 10778 13268 10784 13320
rect 10836 13268 10842 13320
rect 10878 13311 10936 13317
rect 10878 13277 10890 13311
rect 10924 13308 10936 13311
rect 11238 13308 11244 13320
rect 10924 13280 11244 13308
rect 10924 13277 10936 13280
rect 10878 13271 10936 13277
rect 11238 13268 11244 13280
rect 11296 13268 11302 13320
rect 11422 13268 11428 13320
rect 11480 13308 11486 13320
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 11480 13280 11529 13308
rect 11480 13268 11486 13280
rect 11517 13277 11529 13280
rect 11563 13277 11575 13311
rect 11517 13271 11575 13277
rect 11606 13268 11612 13320
rect 11664 13308 11670 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11664 13280 11897 13308
rect 11664 13268 11670 13280
rect 11885 13277 11897 13280
rect 11931 13277 11943 13311
rect 11885 13271 11943 13277
rect 14476 13252 14504 13348
rect 14642 13336 14648 13388
rect 14700 13376 14706 13388
rect 19352 13385 19380 13416
rect 19444 13416 20260 13444
rect 17313 13379 17371 13385
rect 17313 13376 17325 13379
rect 14700 13348 15792 13376
rect 14700 13336 14706 13348
rect 15764 13317 15792 13348
rect 15856 13348 17325 13376
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 15749 13311 15807 13317
rect 15749 13277 15761 13311
rect 15795 13277 15807 13311
rect 15749 13271 15807 13277
rect 10042 13200 10048 13252
rect 10100 13240 10106 13252
rect 10686 13240 10692 13252
rect 10100 13212 10692 13240
rect 10100 13200 10106 13212
rect 10686 13200 10692 13212
rect 10744 13200 10750 13252
rect 11701 13243 11759 13249
rect 11701 13240 11713 13243
rect 10796 13212 11713 13240
rect 7524 13144 8984 13172
rect 9125 13175 9183 13181
rect 7524 13132 7530 13144
rect 9125 13141 9137 13175
rect 9171 13172 9183 13175
rect 9398 13172 9404 13184
rect 9171 13144 9404 13172
rect 9171 13141 9183 13144
rect 9125 13135 9183 13141
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 10226 13132 10232 13184
rect 10284 13172 10290 13184
rect 10796 13172 10824 13212
rect 11701 13209 11713 13212
rect 11747 13209 11759 13243
rect 11701 13203 11759 13209
rect 11790 13200 11796 13252
rect 11848 13200 11854 13252
rect 11992 13212 12434 13240
rect 10284 13144 10824 13172
rect 11057 13175 11115 13181
rect 10284 13132 10290 13144
rect 11057 13141 11069 13175
rect 11103 13172 11115 13175
rect 11992 13172 12020 13212
rect 11103 13144 12020 13172
rect 12406 13172 12434 13212
rect 14458 13200 14464 13252
rect 14516 13200 14522 13252
rect 15580 13240 15608 13271
rect 15856 13240 15884 13348
rect 17313 13345 17325 13348
rect 17359 13345 17371 13379
rect 17313 13339 17371 13345
rect 19337 13379 19395 13385
rect 19337 13345 19349 13379
rect 19383 13345 19395 13379
rect 19337 13339 19395 13345
rect 16301 13311 16359 13317
rect 16301 13277 16313 13311
rect 16347 13308 16359 13311
rect 16482 13308 16488 13320
rect 16347 13280 16488 13308
rect 16347 13277 16359 13280
rect 16301 13271 16359 13277
rect 16482 13268 16488 13280
rect 16540 13308 16546 13320
rect 16945 13311 17003 13317
rect 16945 13308 16957 13311
rect 16540 13280 16957 13308
rect 16540 13268 16546 13280
rect 16945 13277 16957 13280
rect 16991 13277 17003 13311
rect 16945 13271 17003 13277
rect 17034 13268 17040 13320
rect 17092 13308 17098 13320
rect 17129 13311 17187 13317
rect 17129 13308 17141 13311
rect 17092 13280 17141 13308
rect 17092 13268 17098 13280
rect 17129 13277 17141 13280
rect 17175 13277 17187 13311
rect 17129 13271 17187 13277
rect 15580 13212 15884 13240
rect 16117 13243 16175 13249
rect 16117 13209 16129 13243
rect 16163 13209 16175 13243
rect 17144 13240 17172 13271
rect 18138 13268 18144 13320
rect 18196 13308 18202 13320
rect 18785 13311 18843 13317
rect 18785 13308 18797 13311
rect 18196 13280 18797 13308
rect 18196 13268 18202 13280
rect 18785 13277 18797 13280
rect 18831 13277 18843 13311
rect 18785 13271 18843 13277
rect 18969 13311 19027 13317
rect 18969 13277 18981 13311
rect 19015 13277 19027 13311
rect 18969 13271 19027 13277
rect 18322 13240 18328 13252
rect 16117 13203 16175 13209
rect 16316 13212 16988 13240
rect 17144 13212 18328 13240
rect 16132 13172 16160 13203
rect 16316 13184 16344 13212
rect 12406 13144 16160 13172
rect 11103 13141 11115 13144
rect 11057 13135 11115 13141
rect 16298 13132 16304 13184
rect 16356 13132 16362 13184
rect 16574 13132 16580 13184
rect 16632 13172 16638 13184
rect 16853 13175 16911 13181
rect 16853 13172 16865 13175
rect 16632 13144 16865 13172
rect 16632 13132 16638 13144
rect 16853 13141 16865 13144
rect 16899 13141 16911 13175
rect 16960 13172 16988 13212
rect 18322 13200 18328 13212
rect 18380 13200 18386 13252
rect 18984 13240 19012 13271
rect 19242 13268 19248 13320
rect 19300 13268 19306 13320
rect 19334 13240 19340 13252
rect 18984 13212 19340 13240
rect 19334 13200 19340 13212
rect 19392 13200 19398 13252
rect 17310 13172 17316 13184
rect 16960 13144 17316 13172
rect 16853 13135 16911 13141
rect 17310 13132 17316 13144
rect 17368 13172 17374 13184
rect 19444 13172 19472 13416
rect 20254 13404 20260 13416
rect 20312 13444 20318 13456
rect 22940 13444 22968 13472
rect 20312 13416 22968 13444
rect 20312 13404 20318 13416
rect 22186 13376 22192 13388
rect 22066 13348 22192 13376
rect 19518 13268 19524 13320
rect 19576 13268 19582 13320
rect 21726 13268 21732 13320
rect 21784 13268 21790 13320
rect 21913 13311 21971 13317
rect 21913 13277 21925 13311
rect 21959 13308 21971 13311
rect 22066 13308 22094 13348
rect 22186 13336 22192 13348
rect 22244 13376 22250 13388
rect 22646 13376 22652 13388
rect 22244 13348 22652 13376
rect 22244 13336 22250 13348
rect 22646 13336 22652 13348
rect 22704 13376 22710 13388
rect 22704 13348 23336 13376
rect 22704 13336 22710 13348
rect 23308 13320 23336 13348
rect 25130 13336 25136 13388
rect 25188 13376 25194 13388
rect 25225 13379 25283 13385
rect 25225 13376 25237 13379
rect 25188 13348 25237 13376
rect 25188 13336 25194 13348
rect 25225 13345 25237 13348
rect 25271 13376 25283 13379
rect 26234 13376 26240 13388
rect 25271 13348 26240 13376
rect 25271 13345 25283 13348
rect 25225 13339 25283 13345
rect 26206 13336 26240 13348
rect 26292 13336 26298 13388
rect 21959 13280 22094 13308
rect 22925 13311 22983 13317
rect 21959 13277 21971 13280
rect 21913 13271 21971 13277
rect 22925 13277 22937 13311
rect 22971 13277 22983 13311
rect 22925 13271 22983 13277
rect 22940 13240 22968 13271
rect 23290 13268 23296 13320
rect 23348 13268 23354 13320
rect 23750 13268 23756 13320
rect 23808 13268 23814 13320
rect 26206 13308 26234 13336
rect 28813 13311 28871 13317
rect 28813 13308 28825 13311
rect 26206 13280 28825 13308
rect 28813 13277 28825 13280
rect 28859 13277 28871 13311
rect 28813 13271 28871 13277
rect 23768 13240 23796 13268
rect 22940 13212 23796 13240
rect 17368 13144 19472 13172
rect 17368 13132 17374 13144
rect 19702 13132 19708 13184
rect 19760 13132 19766 13184
rect 21818 13132 21824 13184
rect 21876 13132 21882 13184
rect 1104 13082 29595 13104
rect 1104 13030 8032 13082
rect 8084 13030 8096 13082
rect 8148 13030 8160 13082
rect 8212 13030 8224 13082
rect 8276 13030 8288 13082
rect 8340 13030 15115 13082
rect 15167 13030 15179 13082
rect 15231 13030 15243 13082
rect 15295 13030 15307 13082
rect 15359 13030 15371 13082
rect 15423 13030 22198 13082
rect 22250 13030 22262 13082
rect 22314 13030 22326 13082
rect 22378 13030 22390 13082
rect 22442 13030 22454 13082
rect 22506 13030 29281 13082
rect 29333 13030 29345 13082
rect 29397 13030 29409 13082
rect 29461 13030 29473 13082
rect 29525 13030 29537 13082
rect 29589 13030 29595 13082
rect 1104 13008 29595 13030
rect 5166 12968 5172 12980
rect 1780 12940 5172 12968
rect 1394 12792 1400 12844
rect 1452 12832 1458 12844
rect 1780 12841 1808 12940
rect 5166 12928 5172 12940
rect 5224 12968 5230 12980
rect 7098 12968 7104 12980
rect 5224 12940 5396 12968
rect 5224 12928 5230 12940
rect 3510 12860 3516 12912
rect 3568 12860 3574 12912
rect 5368 12909 5396 12940
rect 5920 12940 7104 12968
rect 5920 12909 5948 12940
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 7190 12928 7196 12980
rect 7248 12928 7254 12980
rect 10410 12968 10416 12980
rect 9508 12940 10416 12968
rect 5353 12903 5411 12909
rect 5353 12869 5365 12903
rect 5399 12869 5411 12903
rect 5353 12863 5411 12869
rect 5905 12903 5963 12909
rect 5905 12869 5917 12903
rect 5951 12869 5963 12903
rect 5905 12863 5963 12869
rect 6730 12860 6736 12912
rect 6788 12860 6794 12912
rect 1765 12835 1823 12841
rect 1765 12832 1777 12835
rect 1452 12804 1777 12832
rect 1452 12792 1458 12804
rect 1765 12801 1777 12804
rect 1811 12801 1823 12835
rect 1765 12795 1823 12801
rect 3142 12792 3148 12844
rect 3200 12792 3206 12844
rect 3528 12832 3556 12860
rect 3881 12835 3939 12841
rect 3881 12832 3893 12835
rect 3528 12804 3893 12832
rect 3881 12801 3893 12804
rect 3927 12801 3939 12835
rect 3881 12795 3939 12801
rect 4065 12835 4123 12841
rect 4065 12801 4077 12835
rect 4111 12801 4123 12835
rect 4065 12795 4123 12801
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 4890 12832 4896 12844
rect 4663 12804 4896 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 2038 12724 2044 12776
rect 2096 12724 2102 12776
rect 3789 12767 3847 12773
rect 3789 12733 3801 12767
rect 3835 12764 3847 12767
rect 4080 12764 4108 12795
rect 4890 12792 4896 12804
rect 4948 12792 4954 12844
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12801 5871 12835
rect 5813 12795 5871 12801
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12832 6055 12835
rect 6454 12832 6460 12844
rect 6043 12804 6460 12832
rect 6043 12801 6055 12804
rect 5997 12795 6055 12801
rect 5644 12764 5672 12795
rect 3835 12736 5672 12764
rect 5828 12764 5856 12795
rect 6454 12792 6460 12804
rect 6512 12792 6518 12844
rect 6546 12764 6552 12776
rect 5828 12736 6552 12764
rect 3835 12733 3847 12736
rect 3789 12727 3847 12733
rect 3896 12640 3924 12736
rect 6012 12708 6040 12736
rect 6546 12724 6552 12736
rect 6604 12724 6610 12776
rect 6748 12764 6776 12860
rect 7009 12835 7067 12841
rect 7009 12801 7021 12835
rect 7055 12832 7067 12835
rect 7208 12832 7236 12928
rect 9508 12909 9536 12940
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 10778 12928 10784 12980
rect 10836 12968 10842 12980
rect 10965 12971 11023 12977
rect 10965 12968 10977 12971
rect 10836 12940 10977 12968
rect 10836 12928 10842 12940
rect 10965 12937 10977 12940
rect 11011 12937 11023 12971
rect 10965 12931 11023 12937
rect 11790 12928 11796 12980
rect 11848 12968 11854 12980
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 11848 12940 12173 12968
rect 11848 12928 11854 12940
rect 12161 12937 12173 12940
rect 12207 12937 12219 12971
rect 12161 12931 12219 12937
rect 13262 12928 13268 12980
rect 13320 12968 13326 12980
rect 13320 12940 14320 12968
rect 13320 12928 13326 12940
rect 9493 12903 9551 12909
rect 9493 12869 9505 12903
rect 9539 12869 9551 12903
rect 9493 12863 9551 12869
rect 9950 12860 9956 12912
rect 10008 12860 10014 12912
rect 11422 12860 11428 12912
rect 11480 12860 11486 12912
rect 14292 12909 14320 12940
rect 14642 12928 14648 12980
rect 14700 12928 14706 12980
rect 17221 12971 17279 12977
rect 17221 12968 17233 12971
rect 15028 12940 17233 12968
rect 15028 12909 15056 12940
rect 17221 12937 17233 12940
rect 17267 12937 17279 12971
rect 18414 12968 18420 12980
rect 17221 12931 17279 12937
rect 18340 12940 18420 12968
rect 14001 12903 14059 12909
rect 14001 12900 14013 12903
rect 12268 12872 14013 12900
rect 7055 12804 7236 12832
rect 7055 12801 7067 12804
rect 7009 12795 7067 12801
rect 7282 12792 7288 12844
rect 7340 12792 7346 12844
rect 7558 12792 7564 12844
rect 7616 12792 7622 12844
rect 11440 12832 11468 12860
rect 12268 12841 12296 12872
rect 14001 12869 14013 12872
rect 14047 12869 14059 12903
rect 14001 12863 14059 12869
rect 14277 12903 14335 12909
rect 14277 12869 14289 12903
rect 14323 12869 14335 12903
rect 14277 12863 14335 12869
rect 15013 12903 15071 12909
rect 15013 12869 15025 12903
rect 15059 12869 15071 12903
rect 15013 12863 15071 12869
rect 16482 12860 16488 12912
rect 16540 12860 16546 12912
rect 16574 12860 16580 12912
rect 16632 12860 16638 12912
rect 17402 12900 17408 12912
rect 16776 12872 17408 12900
rect 12253 12835 12311 12841
rect 7760 12804 9168 12832
rect 11440 12804 12204 12832
rect 7193 12767 7251 12773
rect 7193 12764 7205 12767
rect 6748 12736 7205 12764
rect 7193 12733 7205 12736
rect 7239 12764 7251 12767
rect 7760 12764 7788 12804
rect 7239 12736 7788 12764
rect 7837 12767 7895 12773
rect 7239 12733 7251 12736
rect 7193 12727 7251 12733
rect 7837 12733 7849 12767
rect 7883 12764 7895 12767
rect 7883 12736 9076 12764
rect 7883 12733 7895 12736
rect 7837 12727 7895 12733
rect 5994 12656 6000 12708
rect 6052 12656 6058 12708
rect 6270 12656 6276 12708
rect 6328 12696 6334 12708
rect 7852 12696 7880 12727
rect 6328 12668 7880 12696
rect 6328 12656 6334 12668
rect 3878 12588 3884 12640
rect 3936 12588 3942 12640
rect 4246 12588 4252 12640
rect 4304 12588 4310 12640
rect 6178 12588 6184 12640
rect 6236 12588 6242 12640
rect 9048 12628 9076 12736
rect 9140 12696 9168 12804
rect 9214 12724 9220 12776
rect 9272 12724 9278 12776
rect 10042 12764 10048 12776
rect 9324 12736 10048 12764
rect 9324 12696 9352 12736
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 10226 12724 10232 12776
rect 10284 12764 10290 12776
rect 10502 12764 10508 12776
rect 10284 12736 10508 12764
rect 10284 12724 10290 12736
rect 10502 12724 10508 12736
rect 10560 12764 10566 12776
rect 11517 12767 11575 12773
rect 11517 12764 11529 12767
rect 10560 12736 11529 12764
rect 10560 12724 10566 12736
rect 11517 12733 11529 12736
rect 11563 12733 11575 12767
rect 12176 12764 12204 12804
rect 12253 12801 12265 12835
rect 12299 12801 12311 12835
rect 12253 12795 12311 12801
rect 12342 12792 12348 12844
rect 12400 12832 12406 12844
rect 12437 12835 12495 12841
rect 12437 12832 12449 12835
rect 12400 12804 12449 12832
rect 12400 12792 12406 12804
rect 12437 12801 12449 12804
rect 12483 12801 12495 12835
rect 12437 12795 12495 12801
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12801 12587 12835
rect 12529 12795 12587 12801
rect 12544 12764 12572 12795
rect 12618 12792 12624 12844
rect 12676 12792 12682 12844
rect 13449 12835 13507 12841
rect 13449 12801 13461 12835
rect 13495 12832 13507 12835
rect 13814 12832 13820 12844
rect 13495 12804 13820 12832
rect 13495 12801 13507 12804
rect 13449 12795 13507 12801
rect 13814 12792 13820 12804
rect 13872 12832 13878 12844
rect 14093 12835 14151 12841
rect 14093 12832 14105 12835
rect 13872 12804 14105 12832
rect 13872 12792 13878 12804
rect 14093 12801 14105 12804
rect 14139 12801 14151 12835
rect 14093 12795 14151 12801
rect 14366 12792 14372 12844
rect 14424 12792 14430 12844
rect 14458 12792 14464 12844
rect 14516 12792 14522 12844
rect 16114 12792 16120 12844
rect 16172 12792 16178 12844
rect 13998 12764 14004 12776
rect 12176 12736 14004 12764
rect 11517 12727 11575 12733
rect 13998 12724 14004 12736
rect 14056 12764 14062 12776
rect 14642 12764 14648 12776
rect 14056 12736 14648 12764
rect 14056 12724 14062 12736
rect 14642 12724 14648 12736
rect 14700 12724 14706 12776
rect 14734 12724 14740 12776
rect 14792 12764 14798 12776
rect 16500 12773 16528 12860
rect 16592 12832 16620 12860
rect 16669 12835 16727 12841
rect 16669 12832 16681 12835
rect 16592 12804 16681 12832
rect 16669 12801 16681 12804
rect 16715 12801 16727 12835
rect 16669 12795 16727 12801
rect 16485 12767 16543 12773
rect 14792 12736 16436 12764
rect 14792 12724 14798 12736
rect 9140 12668 9352 12696
rect 16408 12696 16436 12736
rect 16485 12733 16497 12767
rect 16531 12733 16543 12767
rect 16485 12727 16543 12733
rect 16574 12724 16580 12776
rect 16632 12764 16638 12776
rect 16776 12764 16804 12872
rect 17402 12860 17408 12872
rect 17460 12900 17466 12912
rect 18340 12909 18368 12940
rect 18414 12928 18420 12940
rect 18472 12928 18478 12980
rect 19610 12928 19616 12980
rect 19668 12968 19674 12980
rect 19978 12968 19984 12980
rect 19668 12940 19984 12968
rect 19668 12928 19674 12940
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 21177 12971 21235 12977
rect 21177 12937 21189 12971
rect 21223 12968 21235 12971
rect 21634 12968 21640 12980
rect 21223 12940 21640 12968
rect 21223 12937 21235 12940
rect 21177 12931 21235 12937
rect 21634 12928 21640 12940
rect 21692 12928 21698 12980
rect 18325 12903 18383 12909
rect 17460 12872 18092 12900
rect 17460 12860 17466 12872
rect 16850 12792 16856 12844
rect 16908 12792 16914 12844
rect 16942 12792 16948 12844
rect 17000 12792 17006 12844
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12832 17095 12835
rect 17126 12832 17132 12844
rect 17083 12804 17132 12832
rect 17083 12801 17095 12804
rect 17037 12795 17095 12801
rect 17126 12792 17132 12804
rect 17184 12792 17190 12844
rect 18064 12773 18092 12872
rect 18325 12869 18337 12903
rect 18371 12869 18383 12903
rect 18325 12863 18383 12869
rect 20806 12860 20812 12912
rect 20864 12900 20870 12912
rect 22005 12903 22063 12909
rect 22005 12900 22017 12903
rect 20864 12872 22017 12900
rect 20864 12860 20870 12872
rect 22005 12869 22017 12872
rect 22051 12869 22063 12903
rect 22005 12863 22063 12869
rect 16632 12736 16804 12764
rect 18049 12767 18107 12773
rect 16632 12724 16638 12736
rect 18049 12733 18061 12767
rect 18095 12733 18107 12767
rect 18049 12727 18107 12733
rect 16592 12696 16620 12724
rect 16408 12668 16620 12696
rect 10502 12628 10508 12640
rect 9048 12600 10508 12628
rect 10502 12588 10508 12600
rect 10560 12628 10566 12640
rect 11238 12628 11244 12640
rect 10560 12600 11244 12628
rect 10560 12588 10566 12600
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 12802 12588 12808 12640
rect 12860 12588 12866 12640
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 14366 12628 14372 12640
rect 13964 12600 14372 12628
rect 13964 12588 13970 12600
rect 14366 12588 14372 12600
rect 14424 12588 14430 12640
rect 16114 12588 16120 12640
rect 16172 12628 16178 12640
rect 17954 12628 17960 12640
rect 16172 12600 17960 12628
rect 16172 12588 16178 12600
rect 17954 12588 17960 12600
rect 18012 12628 18018 12640
rect 19444 12628 19472 12818
rect 20714 12792 20720 12844
rect 20772 12832 20778 12844
rect 21453 12835 21511 12841
rect 21453 12832 21465 12835
rect 20772 12804 21465 12832
rect 20772 12792 20778 12804
rect 21453 12801 21465 12804
rect 21499 12801 21511 12835
rect 21453 12795 21511 12801
rect 21542 12792 21548 12844
rect 21600 12792 21606 12844
rect 21818 12792 21824 12844
rect 21876 12832 21882 12844
rect 23017 12835 23075 12841
rect 23017 12832 23029 12835
rect 21876 12804 23029 12832
rect 21876 12792 21882 12804
rect 23017 12801 23029 12804
rect 23063 12801 23075 12835
rect 23017 12795 23075 12801
rect 23201 12835 23259 12841
rect 23201 12801 23213 12835
rect 23247 12832 23259 12835
rect 23382 12832 23388 12844
rect 23247 12804 23388 12832
rect 23247 12801 23259 12804
rect 23201 12795 23259 12801
rect 20073 12767 20131 12773
rect 20073 12733 20085 12767
rect 20119 12764 20131 12767
rect 20254 12764 20260 12776
rect 20119 12736 20260 12764
rect 20119 12733 20131 12736
rect 20073 12727 20131 12733
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12733 21419 12767
rect 21560 12764 21588 12792
rect 22186 12764 22192 12776
rect 21560 12736 22192 12764
rect 21361 12727 21419 12733
rect 21376 12696 21404 12727
rect 22186 12724 22192 12736
rect 22244 12724 22250 12776
rect 22738 12724 22744 12776
rect 22796 12724 22802 12776
rect 22922 12724 22928 12776
rect 22980 12764 22986 12776
rect 23216 12764 23244 12795
rect 23382 12792 23388 12804
rect 23440 12792 23446 12844
rect 22980 12736 23244 12764
rect 22980 12724 22986 12736
rect 22646 12696 22652 12708
rect 21376 12668 22652 12696
rect 22646 12656 22652 12668
rect 22704 12656 22710 12708
rect 21542 12628 21548 12640
rect 18012 12600 21548 12628
rect 18012 12588 18018 12600
rect 21542 12588 21548 12600
rect 21600 12588 21606 12640
rect 21634 12588 21640 12640
rect 21692 12628 21698 12640
rect 23017 12631 23075 12637
rect 23017 12628 23029 12631
rect 21692 12600 23029 12628
rect 21692 12588 21698 12600
rect 23017 12597 23029 12600
rect 23063 12597 23075 12631
rect 23017 12591 23075 12597
rect 23382 12588 23388 12640
rect 23440 12588 23446 12640
rect 1104 12538 29440 12560
rect 1104 12486 4491 12538
rect 4543 12486 4555 12538
rect 4607 12486 4619 12538
rect 4671 12486 4683 12538
rect 4735 12486 4747 12538
rect 4799 12486 11574 12538
rect 11626 12486 11638 12538
rect 11690 12486 11702 12538
rect 11754 12486 11766 12538
rect 11818 12486 11830 12538
rect 11882 12486 18657 12538
rect 18709 12486 18721 12538
rect 18773 12486 18785 12538
rect 18837 12486 18849 12538
rect 18901 12486 18913 12538
rect 18965 12486 25740 12538
rect 25792 12486 25804 12538
rect 25856 12486 25868 12538
rect 25920 12486 25932 12538
rect 25984 12486 25996 12538
rect 26048 12486 29440 12538
rect 1104 12464 29440 12486
rect 2038 12384 2044 12436
rect 2096 12424 2102 12436
rect 2685 12427 2743 12433
rect 2685 12424 2697 12427
rect 2096 12396 2697 12424
rect 2096 12384 2102 12396
rect 2685 12393 2697 12396
rect 2731 12393 2743 12427
rect 2685 12387 2743 12393
rect 6914 12384 6920 12436
rect 6972 12384 6978 12436
rect 7558 12384 7564 12436
rect 7616 12424 7622 12436
rect 7929 12427 7987 12433
rect 7929 12424 7941 12427
rect 7616 12396 7941 12424
rect 7616 12384 7622 12396
rect 7929 12393 7941 12396
rect 7975 12393 7987 12427
rect 7929 12387 7987 12393
rect 10226 12384 10232 12436
rect 10284 12424 10290 12436
rect 10965 12427 11023 12433
rect 10965 12424 10977 12427
rect 10284 12396 10977 12424
rect 10284 12384 10290 12396
rect 10965 12393 10977 12396
rect 11011 12393 11023 12427
rect 10965 12387 11023 12393
rect 12250 12384 12256 12436
rect 12308 12424 12314 12436
rect 12308 12396 15240 12424
rect 12308 12384 12314 12396
rect 4246 12356 4252 12368
rect 2976 12328 4252 12356
rect 2976 12229 3004 12328
rect 4246 12316 4252 12328
rect 4304 12316 4310 12368
rect 3510 12248 3516 12300
rect 3568 12248 3574 12300
rect 4525 12291 4583 12297
rect 4525 12257 4537 12291
rect 4571 12288 4583 12291
rect 4982 12288 4988 12300
rect 4571 12260 4988 12288
rect 4571 12257 4583 12260
rect 4525 12251 4583 12257
rect 4982 12248 4988 12260
rect 5040 12248 5046 12300
rect 5166 12248 5172 12300
rect 5224 12248 5230 12300
rect 5445 12291 5503 12297
rect 5445 12257 5457 12291
rect 5491 12288 5503 12291
rect 6178 12288 6184 12300
rect 5491 12260 6184 12288
rect 5491 12257 5503 12260
rect 5445 12251 5503 12257
rect 6178 12248 6184 12260
rect 6236 12248 6242 12300
rect 6932 12288 6960 12384
rect 7190 12316 7196 12368
rect 7248 12356 7254 12368
rect 15102 12356 15108 12368
rect 7248 12328 7788 12356
rect 7248 12316 7254 12328
rect 7377 12291 7435 12297
rect 7377 12288 7389 12291
rect 6932 12260 7389 12288
rect 7377 12257 7389 12260
rect 7423 12257 7435 12291
rect 7377 12251 7435 12257
rect 7466 12248 7472 12300
rect 7524 12288 7530 12300
rect 7561 12291 7619 12297
rect 7561 12288 7573 12291
rect 7524 12260 7573 12288
rect 7524 12248 7530 12260
rect 7561 12257 7573 12260
rect 7607 12257 7619 12291
rect 7561 12251 7619 12257
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12189 2927 12223
rect 2869 12183 2927 12189
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12189 3019 12223
rect 2961 12183 3019 12189
rect 2884 12084 2912 12183
rect 3050 12180 3056 12232
rect 3108 12180 3114 12232
rect 3234 12229 3240 12232
rect 3191 12223 3240 12229
rect 3191 12189 3203 12223
rect 3237 12189 3240 12223
rect 3191 12183 3240 12189
rect 3234 12180 3240 12183
rect 3292 12180 3298 12232
rect 3329 12223 3387 12229
rect 3329 12189 3341 12223
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 3421 12223 3479 12229
rect 3421 12189 3433 12223
rect 3467 12220 3479 12223
rect 3528 12220 3556 12248
rect 3467 12192 3556 12220
rect 3605 12223 3663 12229
rect 3467 12189 3479 12192
rect 3421 12183 3479 12189
rect 3605 12189 3617 12223
rect 3651 12220 3663 12223
rect 3651 12192 3924 12220
rect 3651 12189 3663 12192
rect 3605 12183 3663 12189
rect 3344 12152 3372 12183
rect 3620 12152 3648 12183
rect 3344 12124 3648 12152
rect 3896 12096 3924 12192
rect 4430 12180 4436 12232
rect 4488 12180 4494 12232
rect 4614 12180 4620 12232
rect 4672 12180 4678 12232
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 4724 12152 4752 12183
rect 7190 12180 7196 12232
rect 7248 12180 7254 12232
rect 7285 12223 7343 12229
rect 7285 12189 7297 12223
rect 7331 12220 7343 12223
rect 7484 12220 7512 12248
rect 7760 12229 7788 12328
rect 13740 12328 15108 12356
rect 9214 12248 9220 12300
rect 9272 12288 9278 12300
rect 11793 12291 11851 12297
rect 11793 12288 11805 12291
rect 9272 12260 11805 12288
rect 9272 12248 9278 12260
rect 11793 12257 11805 12260
rect 11839 12288 11851 12291
rect 12066 12288 12072 12300
rect 11839 12260 12072 12288
rect 11839 12257 11851 12260
rect 11793 12251 11851 12257
rect 12066 12248 12072 12260
rect 12124 12288 12130 12300
rect 12161 12291 12219 12297
rect 12161 12288 12173 12291
rect 12124 12260 12173 12288
rect 12124 12248 12130 12260
rect 12161 12257 12173 12260
rect 12207 12257 12219 12291
rect 12161 12251 12219 12257
rect 12437 12291 12495 12297
rect 12437 12257 12449 12291
rect 12483 12288 12495 12291
rect 13740 12288 13768 12328
rect 15102 12316 15108 12328
rect 15160 12316 15166 12368
rect 12483 12260 13768 12288
rect 12483 12257 12495 12260
rect 12437 12251 12495 12257
rect 7331 12192 7512 12220
rect 7745 12223 7803 12229
rect 7331 12189 7343 12192
rect 7285 12183 7343 12189
rect 7745 12189 7757 12223
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 13906 12180 13912 12232
rect 13964 12220 13970 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13964 12192 14105 12220
rect 13964 12180 13970 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 14642 12180 14648 12232
rect 14700 12180 14706 12232
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12220 14795 12223
rect 14829 12223 14887 12229
rect 14829 12220 14841 12223
rect 14783 12192 14841 12220
rect 14783 12189 14795 12192
rect 14737 12183 14795 12189
rect 14829 12189 14841 12192
rect 14875 12189 14887 12223
rect 14829 12183 14887 12189
rect 14918 12180 14924 12232
rect 14976 12220 14982 12232
rect 15212 12229 15240 12396
rect 15286 12316 15292 12368
rect 15344 12356 15350 12368
rect 15381 12359 15439 12365
rect 15381 12356 15393 12359
rect 15344 12328 15393 12356
rect 15344 12316 15350 12328
rect 15381 12325 15393 12328
rect 15427 12325 15439 12359
rect 15381 12319 15439 12325
rect 15746 12316 15752 12368
rect 15804 12356 15810 12368
rect 15804 12328 16712 12356
rect 15804 12316 15810 12328
rect 16684 12232 16712 12328
rect 22922 12316 22928 12368
rect 22980 12356 22986 12368
rect 23290 12356 23296 12368
rect 22980 12328 23296 12356
rect 22980 12316 22986 12328
rect 23290 12316 23296 12328
rect 23348 12316 23354 12368
rect 16758 12248 16764 12300
rect 16816 12248 16822 12300
rect 23014 12248 23020 12300
rect 23072 12248 23078 12300
rect 23382 12248 23388 12300
rect 23440 12288 23446 12300
rect 23440 12260 24072 12288
rect 23440 12248 23446 12260
rect 15013 12223 15071 12229
rect 15013 12220 15025 12223
rect 14976 12192 15025 12220
rect 14976 12180 14982 12192
rect 15013 12189 15025 12192
rect 15059 12189 15071 12223
rect 15013 12183 15071 12189
rect 15197 12223 15255 12229
rect 15197 12189 15209 12223
rect 15243 12189 15255 12223
rect 15197 12183 15255 12189
rect 16114 12180 16120 12232
rect 16172 12180 16178 12232
rect 16666 12180 16672 12232
rect 16724 12180 16730 12232
rect 19702 12180 19708 12232
rect 19760 12220 19766 12232
rect 19981 12223 20039 12229
rect 19981 12220 19993 12223
rect 19760 12192 19993 12220
rect 19760 12180 19766 12192
rect 19981 12189 19993 12192
rect 20027 12189 20039 12223
rect 19981 12183 20039 12189
rect 22186 12180 22192 12232
rect 22244 12220 22250 12232
rect 22557 12223 22615 12229
rect 22557 12220 22569 12223
rect 22244 12192 22569 12220
rect 22244 12180 22250 12192
rect 22557 12189 22569 12192
rect 22603 12189 22615 12223
rect 22557 12183 22615 12189
rect 5350 12152 5356 12164
rect 4724 12124 5356 12152
rect 5350 12112 5356 12124
rect 5408 12152 5414 12164
rect 9493 12155 9551 12161
rect 5408 12124 5672 12152
rect 6670 12124 7696 12152
rect 5408 12112 5414 12124
rect 3513 12087 3571 12093
rect 3513 12084 3525 12087
rect 2884 12056 3525 12084
rect 3513 12053 3525 12056
rect 3559 12053 3571 12087
rect 3513 12047 3571 12053
rect 3878 12044 3884 12096
rect 3936 12044 3942 12096
rect 4249 12087 4307 12093
rect 4249 12053 4261 12087
rect 4295 12084 4307 12087
rect 5534 12084 5540 12096
rect 4295 12056 5540 12084
rect 4295 12053 4307 12056
rect 4249 12047 4307 12053
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 5644 12084 5672 12124
rect 6362 12084 6368 12096
rect 5644 12056 6368 12084
rect 6362 12044 6368 12056
rect 6420 12044 6426 12096
rect 7006 12044 7012 12096
rect 7064 12044 7070 12096
rect 7668 12084 7696 12124
rect 9493 12121 9505 12155
rect 9539 12152 9551 12155
rect 9766 12152 9772 12164
rect 9539 12124 9772 12152
rect 9539 12121 9551 12124
rect 9493 12115 9551 12121
rect 9766 12112 9772 12124
rect 9824 12112 9830 12164
rect 10042 12112 10048 12164
rect 10100 12112 10106 12164
rect 10962 12112 10968 12164
rect 11020 12152 11026 12164
rect 11057 12155 11115 12161
rect 11057 12152 11069 12155
rect 11020 12124 11069 12152
rect 11020 12112 11026 12124
rect 11057 12121 11069 12124
rect 11103 12152 11115 12155
rect 12526 12152 12532 12164
rect 11103 12124 12532 12152
rect 11103 12121 11115 12124
rect 11057 12115 11115 12121
rect 12526 12112 12532 12124
rect 12584 12112 12590 12164
rect 13722 12152 13728 12164
rect 13662 12124 13728 12152
rect 13722 12112 13728 12124
rect 13780 12112 13786 12164
rect 9582 12084 9588 12096
rect 7668 12056 9588 12084
rect 9582 12044 9588 12056
rect 9640 12084 9646 12096
rect 9858 12084 9864 12096
rect 9640 12056 9864 12084
rect 9640 12044 9646 12056
rect 9858 12044 9864 12056
rect 9916 12044 9922 12096
rect 13924 12093 13952 12180
rect 14660 12152 14688 12180
rect 15105 12155 15163 12161
rect 15105 12152 15117 12155
rect 14660 12124 15117 12152
rect 15105 12121 15117 12124
rect 15151 12152 15163 12155
rect 16942 12152 16948 12164
rect 15151 12124 16948 12152
rect 15151 12121 15163 12124
rect 15105 12115 15163 12121
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 22572 12152 22600 12183
rect 22646 12180 22652 12232
rect 22704 12220 22710 12232
rect 22925 12223 22983 12229
rect 22925 12220 22937 12223
rect 22704 12192 22937 12220
rect 22704 12180 22710 12192
rect 22925 12189 22937 12192
rect 22971 12220 22983 12223
rect 23290 12220 23296 12232
rect 22971 12192 23296 12220
rect 22971 12189 22983 12192
rect 22925 12183 22983 12189
rect 23290 12180 23296 12192
rect 23348 12180 23354 12232
rect 24044 12229 24072 12260
rect 24029 12223 24087 12229
rect 24029 12189 24041 12223
rect 24075 12189 24087 12223
rect 24029 12183 24087 12189
rect 22572 12124 22692 12152
rect 22664 12096 22692 12124
rect 23014 12112 23020 12164
rect 23072 12152 23078 12164
rect 23385 12155 23443 12161
rect 23385 12152 23397 12155
rect 23072 12124 23397 12152
rect 23072 12112 23078 12124
rect 23385 12121 23397 12124
rect 23431 12121 23443 12155
rect 23385 12115 23443 12121
rect 23750 12112 23756 12164
rect 23808 12152 23814 12164
rect 23808 12124 24348 12152
rect 23808 12112 23814 12124
rect 24320 12096 24348 12124
rect 13909 12087 13967 12093
rect 13909 12053 13921 12087
rect 13955 12053 13967 12087
rect 13909 12047 13967 12053
rect 16025 12087 16083 12093
rect 16025 12053 16037 12087
rect 16071 12084 16083 12087
rect 16758 12084 16764 12096
rect 16071 12056 16764 12084
rect 16071 12053 16083 12056
rect 16025 12047 16083 12053
rect 16758 12044 16764 12056
rect 16816 12044 16822 12096
rect 19794 12044 19800 12096
rect 19852 12044 19858 12096
rect 22646 12044 22652 12096
rect 22704 12044 22710 12096
rect 22830 12044 22836 12096
rect 22888 12084 22894 12096
rect 23474 12084 23480 12096
rect 22888 12056 23480 12084
rect 22888 12044 22894 12056
rect 23474 12044 23480 12056
rect 23532 12044 23538 12096
rect 23842 12044 23848 12096
rect 23900 12044 23906 12096
rect 24302 12044 24308 12096
rect 24360 12044 24366 12096
rect 1104 11994 29595 12016
rect 1104 11942 8032 11994
rect 8084 11942 8096 11994
rect 8148 11942 8160 11994
rect 8212 11942 8224 11994
rect 8276 11942 8288 11994
rect 8340 11942 15115 11994
rect 15167 11942 15179 11994
rect 15231 11942 15243 11994
rect 15295 11942 15307 11994
rect 15359 11942 15371 11994
rect 15423 11942 22198 11994
rect 22250 11942 22262 11994
rect 22314 11942 22326 11994
rect 22378 11942 22390 11994
rect 22442 11942 22454 11994
rect 22506 11942 29281 11994
rect 29333 11942 29345 11994
rect 29397 11942 29409 11994
rect 29461 11942 29473 11994
rect 29525 11942 29537 11994
rect 29589 11942 29595 11994
rect 1104 11920 29595 11942
rect 4065 11883 4123 11889
rect 4065 11849 4077 11883
rect 4111 11880 4123 11883
rect 4430 11880 4436 11892
rect 4111 11852 4436 11880
rect 4111 11849 4123 11852
rect 4065 11843 4123 11849
rect 4430 11840 4436 11852
rect 4488 11840 4494 11892
rect 4982 11840 4988 11892
rect 5040 11880 5046 11892
rect 7009 11883 7067 11889
rect 7009 11880 7021 11883
rect 5040 11852 7021 11880
rect 5040 11840 5046 11852
rect 7009 11849 7021 11852
rect 7055 11880 7067 11883
rect 7190 11880 7196 11892
rect 7055 11852 7196 11880
rect 7055 11849 7067 11852
rect 7009 11843 7067 11849
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 7466 11840 7472 11892
rect 7524 11880 7530 11892
rect 10226 11880 10232 11892
rect 7524 11852 10232 11880
rect 7524 11840 7530 11852
rect 10226 11840 10232 11852
rect 10284 11880 10290 11892
rect 12710 11880 12716 11892
rect 10284 11852 10916 11880
rect 10284 11840 10290 11852
rect 3142 11772 3148 11824
rect 3200 11772 3206 11824
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 992 11716 1409 11744
rect 992 11704 998 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11744 1823 11747
rect 2222 11744 2228 11756
rect 1811 11716 2228 11744
rect 1811 11713 1823 11716
rect 1765 11707 1823 11713
rect 2222 11704 2228 11716
rect 2280 11704 2286 11756
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11744 4307 11747
rect 4448 11744 4476 11840
rect 4890 11772 4896 11824
rect 4948 11772 4954 11824
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 6457 11815 6515 11821
rect 6457 11812 6469 11815
rect 6420 11784 6469 11812
rect 6420 11772 6426 11784
rect 6457 11781 6469 11784
rect 6503 11781 6515 11815
rect 7484 11812 7512 11840
rect 6457 11775 6515 11781
rect 6845 11784 7512 11812
rect 4295 11716 4476 11744
rect 4295 11713 4307 11716
rect 4249 11707 4307 11713
rect 2317 11679 2375 11685
rect 2317 11645 2329 11679
rect 2363 11645 2375 11679
rect 2317 11639 2375 11645
rect 2593 11679 2651 11685
rect 2593 11645 2605 11679
rect 2639 11676 2651 11679
rect 4338 11676 4344 11688
rect 2639 11648 4344 11676
rect 2639 11645 2651 11648
rect 2593 11639 2651 11645
rect 2222 11500 2228 11552
rect 2280 11540 2286 11552
rect 2332 11540 2360 11639
rect 4338 11636 4344 11648
rect 4396 11636 4402 11688
rect 5442 11676 5448 11688
rect 4632 11648 5448 11676
rect 4632 11608 4660 11648
rect 5442 11636 5448 11648
rect 5500 11676 5506 11688
rect 5629 11679 5687 11685
rect 5629 11676 5641 11679
rect 5500 11648 5641 11676
rect 5500 11636 5506 11648
rect 5629 11645 5641 11648
rect 5675 11645 5687 11679
rect 5629 11639 5687 11645
rect 4172 11580 4660 11608
rect 4172 11540 4200 11580
rect 4706 11568 4712 11620
rect 4764 11608 4770 11620
rect 6454 11608 6460 11620
rect 4764 11580 6460 11608
rect 4764 11568 4770 11580
rect 6454 11568 6460 11580
rect 6512 11608 6518 11620
rect 6845 11608 6873 11784
rect 9858 11772 9864 11824
rect 9916 11772 9922 11824
rect 10888 11821 10916 11852
rect 12360 11852 12716 11880
rect 12360 11821 12388 11852
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 13814 11840 13820 11892
rect 13872 11840 13878 11892
rect 16224 11852 16620 11880
rect 10873 11815 10931 11821
rect 10873 11781 10885 11815
rect 10919 11781 10931 11815
rect 10873 11775 10931 11781
rect 12345 11815 12403 11821
rect 12345 11781 12357 11815
rect 12391 11781 12403 11815
rect 12345 11775 12403 11781
rect 13909 11815 13967 11821
rect 13909 11781 13921 11815
rect 13955 11812 13967 11815
rect 14274 11812 14280 11824
rect 13955 11784 14280 11812
rect 13955 11781 13967 11784
rect 13909 11775 13967 11781
rect 14274 11772 14280 11784
rect 14332 11772 14338 11824
rect 16224 11821 16252 11852
rect 16209 11815 16267 11821
rect 16209 11781 16221 11815
rect 16255 11781 16267 11815
rect 16592 11812 16620 11852
rect 19978 11840 19984 11892
rect 20036 11840 20042 11892
rect 23290 11840 23296 11892
rect 23348 11880 23354 11892
rect 23753 11883 23811 11889
rect 23753 11880 23765 11883
rect 23348 11852 23765 11880
rect 23348 11840 23354 11852
rect 23753 11849 23765 11852
rect 23799 11849 23811 11883
rect 23753 11843 23811 11849
rect 21726 11812 21732 11824
rect 16592 11784 21732 11812
rect 16209 11775 16267 11781
rect 21726 11772 21732 11784
rect 21784 11772 21790 11824
rect 24118 11812 24124 11824
rect 22572 11784 24124 11812
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11744 6975 11747
rect 7282 11744 7288 11756
rect 6963 11716 7288 11744
rect 6963 11713 6975 11716
rect 6917 11707 6975 11713
rect 7282 11704 7288 11716
rect 7340 11744 7346 11756
rect 7561 11747 7619 11753
rect 7561 11744 7573 11747
rect 7340 11716 7573 11744
rect 7340 11704 7346 11716
rect 7561 11713 7573 11716
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 10459 11747 10517 11753
rect 10459 11713 10471 11747
rect 10505 11744 10517 11747
rect 10597 11747 10655 11753
rect 10597 11744 10609 11747
rect 10505 11716 10609 11744
rect 10505 11713 10517 11716
rect 10459 11707 10517 11713
rect 10597 11713 10609 11716
rect 10643 11713 10655 11747
rect 10597 11707 10655 11713
rect 12066 11704 12072 11756
rect 12124 11704 12130 11756
rect 13722 11744 13728 11756
rect 13478 11730 13728 11744
rect 13464 11716 13728 11730
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11676 8723 11679
rect 8938 11676 8944 11688
rect 8711 11648 8944 11676
rect 8711 11645 8723 11648
rect 8665 11639 8723 11645
rect 8938 11636 8944 11648
rect 8996 11636 9002 11688
rect 9033 11679 9091 11685
rect 9033 11645 9045 11679
rect 9079 11676 9091 11679
rect 9766 11676 9772 11688
rect 9079 11648 9772 11676
rect 9079 11645 9091 11648
rect 9033 11639 9091 11645
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 12986 11636 12992 11688
rect 13044 11676 13050 11688
rect 13464 11676 13492 11716
rect 13722 11704 13728 11716
rect 13780 11704 13786 11756
rect 14090 11704 14096 11756
rect 14148 11744 14154 11756
rect 14642 11744 14648 11756
rect 14148 11716 14648 11744
rect 14148 11704 14154 11716
rect 14642 11704 14648 11716
rect 14700 11704 14706 11756
rect 15470 11704 15476 11756
rect 15528 11744 15534 11756
rect 15746 11744 15752 11756
rect 15528 11716 15752 11744
rect 15528 11704 15534 11716
rect 15746 11704 15752 11716
rect 15804 11744 15810 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15804 11716 15945 11744
rect 15804 11704 15810 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 16117 11747 16175 11753
rect 16117 11713 16129 11747
rect 16163 11713 16175 11747
rect 16117 11707 16175 11713
rect 13044 11648 13492 11676
rect 13044 11636 13050 11648
rect 15838 11636 15844 11688
rect 15896 11676 15902 11688
rect 16132 11676 16160 11707
rect 16298 11704 16304 11756
rect 16356 11704 16362 11756
rect 16684 11716 18184 11744
rect 16390 11676 16396 11688
rect 15896 11648 16396 11676
rect 15896 11636 15902 11648
rect 16390 11636 16396 11648
rect 16448 11676 16454 11688
rect 16684 11676 16712 11716
rect 16448 11648 16712 11676
rect 17037 11679 17095 11685
rect 16448 11636 16454 11648
rect 17037 11645 17049 11679
rect 17083 11676 17095 11679
rect 18046 11676 18052 11688
rect 17083 11648 18052 11676
rect 17083 11645 17095 11648
rect 17037 11639 17095 11645
rect 18046 11636 18052 11648
rect 18104 11636 18110 11688
rect 18156 11676 18184 11716
rect 18506 11704 18512 11756
rect 18564 11704 18570 11756
rect 19334 11704 19340 11756
rect 19392 11704 19398 11756
rect 19797 11747 19855 11753
rect 19797 11713 19809 11747
rect 19843 11744 19855 11747
rect 20257 11747 20315 11753
rect 19843 11716 20116 11744
rect 19843 11713 19855 11716
rect 19797 11707 19855 11713
rect 18156 11648 19472 11676
rect 6512 11580 6873 11608
rect 14200 11580 16620 11608
rect 6512 11568 6518 11580
rect 2280 11512 4200 11540
rect 2280 11500 2286 11512
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 4801 11543 4859 11549
rect 4801 11540 4813 11543
rect 4304 11512 4813 11540
rect 4304 11500 4310 11512
rect 4801 11509 4813 11512
rect 4847 11509 4859 11543
rect 4801 11503 4859 11509
rect 7190 11500 7196 11552
rect 7248 11500 7254 11552
rect 7374 11500 7380 11552
rect 7432 11540 7438 11552
rect 8205 11543 8263 11549
rect 8205 11540 8217 11543
rect 7432 11512 8217 11540
rect 7432 11500 7438 11512
rect 8205 11509 8217 11512
rect 8251 11509 8263 11543
rect 8205 11503 8263 11509
rect 11146 11500 11152 11552
rect 11204 11540 11210 11552
rect 14200 11540 14228 11580
rect 11204 11512 14228 11540
rect 11204 11500 11210 11512
rect 14274 11500 14280 11552
rect 14332 11540 14338 11552
rect 14734 11540 14740 11552
rect 14332 11512 14740 11540
rect 14332 11500 14338 11512
rect 14734 11500 14740 11512
rect 14792 11500 14798 11552
rect 16114 11500 16120 11552
rect 16172 11540 16178 11552
rect 16485 11543 16543 11549
rect 16485 11540 16497 11543
rect 16172 11512 16497 11540
rect 16172 11500 16178 11512
rect 16485 11509 16497 11512
rect 16531 11509 16543 11543
rect 16592 11540 16620 11580
rect 16666 11568 16672 11620
rect 16724 11608 16730 11620
rect 18417 11611 18475 11617
rect 18417 11608 18429 11611
rect 16724 11580 18429 11608
rect 16724 11568 16730 11580
rect 18417 11577 18429 11580
rect 18463 11577 18475 11611
rect 18417 11571 18475 11577
rect 19444 11552 19472 11648
rect 20088 11620 20116 11716
rect 20257 11713 20269 11747
rect 20303 11744 20315 11747
rect 20346 11744 20352 11756
rect 20303 11716 20352 11744
rect 20303 11713 20315 11716
rect 20257 11707 20315 11713
rect 20346 11704 20352 11716
rect 20404 11704 20410 11756
rect 20533 11747 20591 11753
rect 20533 11713 20545 11747
rect 20579 11713 20591 11747
rect 20533 11707 20591 11713
rect 20070 11568 20076 11620
rect 20128 11568 20134 11620
rect 20254 11568 20260 11620
rect 20312 11608 20318 11620
rect 20548 11608 20576 11707
rect 21744 11676 21772 11772
rect 22572 11756 22600 11784
rect 24118 11772 24124 11784
rect 24176 11772 24182 11824
rect 21821 11747 21879 11753
rect 21821 11713 21833 11747
rect 21867 11744 21879 11747
rect 22094 11744 22100 11756
rect 21867 11716 22100 11744
rect 21867 11713 21879 11716
rect 21821 11707 21879 11713
rect 22094 11704 22100 11716
rect 22152 11704 22158 11756
rect 22554 11704 22560 11756
rect 22612 11704 22618 11756
rect 22646 11704 22652 11756
rect 22704 11744 22710 11756
rect 22833 11747 22891 11753
rect 22833 11744 22845 11747
rect 22704 11716 22845 11744
rect 22704 11704 22710 11716
rect 22833 11713 22845 11716
rect 22879 11713 22891 11747
rect 22833 11707 22891 11713
rect 23290 11704 23296 11756
rect 23348 11744 23354 11756
rect 23477 11747 23535 11753
rect 23477 11744 23489 11747
rect 23348 11716 23489 11744
rect 23348 11704 23354 11716
rect 23477 11713 23489 11716
rect 23523 11744 23535 11747
rect 23937 11747 23995 11753
rect 23937 11744 23949 11747
rect 23523 11716 23949 11744
rect 23523 11713 23535 11716
rect 23477 11707 23535 11713
rect 23937 11713 23949 11716
rect 23983 11713 23995 11747
rect 23937 11707 23995 11713
rect 24026 11704 24032 11756
rect 24084 11744 24090 11756
rect 24213 11747 24271 11753
rect 24213 11744 24225 11747
rect 24084 11716 24225 11744
rect 24084 11704 24090 11716
rect 24213 11713 24225 11716
rect 24259 11713 24271 11747
rect 24213 11707 24271 11713
rect 25685 11747 25743 11753
rect 25685 11713 25697 11747
rect 25731 11713 25743 11747
rect 25685 11707 25743 11713
rect 21744 11648 22876 11676
rect 22554 11608 22560 11620
rect 20312 11580 22560 11608
rect 20312 11568 20318 11580
rect 22554 11568 22560 11580
rect 22612 11568 22618 11620
rect 22848 11608 22876 11648
rect 22922 11636 22928 11688
rect 22980 11676 22986 11688
rect 23017 11679 23075 11685
rect 23017 11676 23029 11679
rect 22980 11648 23029 11676
rect 22980 11636 22986 11648
rect 23017 11645 23029 11648
rect 23063 11645 23075 11679
rect 23017 11639 23075 11645
rect 23569 11679 23627 11685
rect 23569 11645 23581 11679
rect 23615 11676 23627 11679
rect 23658 11676 23664 11688
rect 23615 11648 23664 11676
rect 23615 11645 23627 11648
rect 23569 11639 23627 11645
rect 23658 11636 23664 11648
rect 23716 11636 23722 11688
rect 24302 11636 24308 11688
rect 24360 11676 24366 11688
rect 25593 11679 25651 11685
rect 25593 11676 25605 11679
rect 24360 11648 25605 11676
rect 24360 11636 24366 11648
rect 25593 11645 25605 11648
rect 25639 11645 25651 11679
rect 25593 11639 25651 11645
rect 25700 11608 25728 11707
rect 26694 11608 26700 11620
rect 22848 11580 26700 11608
rect 26694 11568 26700 11580
rect 26752 11568 26758 11620
rect 16942 11540 16948 11552
rect 16592 11512 16948 11540
rect 16485 11503 16543 11509
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 17586 11500 17592 11552
rect 17644 11500 17650 11552
rect 19426 11500 19432 11552
rect 19484 11540 19490 11552
rect 21450 11540 21456 11552
rect 19484 11512 21456 11540
rect 19484 11500 19490 11512
rect 21450 11500 21456 11512
rect 21508 11500 21514 11552
rect 24118 11500 24124 11552
rect 24176 11500 24182 11552
rect 24397 11543 24455 11549
rect 24397 11509 24409 11543
rect 24443 11540 24455 11543
rect 25590 11540 25596 11552
rect 24443 11512 25596 11540
rect 24443 11509 24455 11512
rect 24397 11503 24455 11509
rect 25590 11500 25596 11512
rect 25648 11500 25654 11552
rect 26053 11543 26111 11549
rect 26053 11509 26065 11543
rect 26099 11540 26111 11543
rect 26234 11540 26240 11552
rect 26099 11512 26240 11540
rect 26099 11509 26111 11512
rect 26053 11503 26111 11509
rect 26234 11500 26240 11512
rect 26292 11500 26298 11552
rect 1104 11450 29440 11472
rect 1104 11398 4491 11450
rect 4543 11398 4555 11450
rect 4607 11398 4619 11450
rect 4671 11398 4683 11450
rect 4735 11398 4747 11450
rect 4799 11398 11574 11450
rect 11626 11398 11638 11450
rect 11690 11398 11702 11450
rect 11754 11398 11766 11450
rect 11818 11398 11830 11450
rect 11882 11398 18657 11450
rect 18709 11398 18721 11450
rect 18773 11398 18785 11450
rect 18837 11398 18849 11450
rect 18901 11398 18913 11450
rect 18965 11398 25740 11450
rect 25792 11398 25804 11450
rect 25856 11398 25868 11450
rect 25920 11398 25932 11450
rect 25984 11398 25996 11450
rect 26048 11398 29440 11450
rect 1104 11376 29440 11398
rect 2120 11339 2178 11345
rect 2120 11305 2132 11339
rect 2166 11336 2178 11339
rect 4154 11336 4160 11348
rect 2166 11308 4160 11336
rect 2166 11305 2178 11308
rect 2120 11299 2178 11305
rect 4154 11296 4160 11308
rect 4212 11296 4218 11348
rect 4338 11296 4344 11348
rect 4396 11296 4402 11348
rect 4890 11296 4896 11348
rect 4948 11336 4954 11348
rect 5708 11339 5766 11345
rect 4948 11308 5580 11336
rect 4948 11296 4954 11308
rect 3605 11271 3663 11277
rect 3605 11237 3617 11271
rect 3651 11268 3663 11271
rect 4246 11268 4252 11280
rect 3651 11240 4252 11268
rect 3651 11237 3663 11240
rect 3605 11231 3663 11237
rect 4246 11228 4252 11240
rect 4304 11228 4310 11280
rect 4798 11268 4804 11280
rect 4448 11240 4804 11268
rect 1857 11203 1915 11209
rect 1857 11169 1869 11203
rect 1903 11200 1915 11203
rect 2222 11200 2228 11212
rect 1903 11172 2228 11200
rect 1903 11169 1915 11172
rect 1857 11163 1915 11169
rect 2222 11160 2228 11172
rect 2280 11160 2286 11212
rect 4062 11200 4068 11212
rect 3804 11172 4068 11200
rect 3142 11092 3148 11144
rect 3200 11132 3206 11144
rect 3804 11141 3832 11172
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 3789 11135 3847 11141
rect 3200 11104 3266 11132
rect 3200 11092 3206 11104
rect 3789 11101 3801 11135
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 3970 11092 3976 11144
rect 4028 11092 4034 11144
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4448 11132 4476 11240
rect 4798 11228 4804 11240
rect 4856 11268 4862 11280
rect 5166 11268 5172 11280
rect 4856 11240 5172 11268
rect 4856 11228 4862 11240
rect 5166 11228 5172 11240
rect 5224 11228 5230 11280
rect 5074 11160 5080 11212
rect 5132 11160 5138 11212
rect 5442 11160 5448 11212
rect 5500 11160 5506 11212
rect 5552 11200 5580 11308
rect 5708 11305 5720 11339
rect 5754 11336 5766 11339
rect 7837 11339 7895 11345
rect 7837 11336 7849 11339
rect 5754 11308 7849 11336
rect 5754 11305 5766 11308
rect 5708 11299 5766 11305
rect 7837 11305 7849 11308
rect 7883 11305 7895 11339
rect 17586 11336 17592 11348
rect 7837 11299 7895 11305
rect 15948 11308 17592 11336
rect 7193 11271 7251 11277
rect 7193 11237 7205 11271
rect 7239 11268 7251 11271
rect 7282 11268 7288 11280
rect 7239 11240 7288 11268
rect 7239 11237 7251 11240
rect 7193 11231 7251 11237
rect 7282 11228 7288 11240
rect 7340 11228 7346 11280
rect 9674 11228 9680 11280
rect 9732 11268 9738 11280
rect 10502 11268 10508 11280
rect 9732 11240 10508 11268
rect 9732 11228 9738 11240
rect 10502 11228 10508 11240
rect 10560 11228 10566 11280
rect 5552 11172 9674 11200
rect 4203 11104 4476 11132
rect 4525 11135 4583 11141
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4525 11101 4537 11135
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 3878 11024 3884 11076
rect 3936 11064 3942 11076
rect 4065 11067 4123 11073
rect 4065 11064 4077 11067
rect 3936 11036 4077 11064
rect 3936 11024 3942 11036
rect 4065 11033 4077 11036
rect 4111 11033 4123 11067
rect 4065 11027 4123 11033
rect 4080 10996 4108 11027
rect 4246 11024 4252 11076
rect 4304 11064 4310 11076
rect 4540 11064 4568 11095
rect 4798 11092 4804 11144
rect 4856 11132 4862 11144
rect 5092 11132 5120 11160
rect 4856 11104 5120 11132
rect 7285 11135 7343 11141
rect 4856 11092 4862 11104
rect 7285 11101 7297 11135
rect 7331 11132 7343 11135
rect 7374 11132 7380 11144
rect 7331 11104 7380 11132
rect 7331 11101 7343 11104
rect 7285 11095 7343 11101
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 7466 11092 7472 11144
rect 7524 11092 7530 11144
rect 7653 11135 7711 11141
rect 7653 11101 7665 11135
rect 7699 11132 7711 11135
rect 7834 11132 7840 11144
rect 7699 11104 7840 11132
rect 7699 11101 7711 11104
rect 7653 11095 7711 11101
rect 7834 11092 7840 11104
rect 7892 11092 7898 11144
rect 9646 11132 9674 11172
rect 9953 11135 10011 11141
rect 9953 11132 9965 11135
rect 9646 11104 9965 11132
rect 9953 11101 9965 11104
rect 9999 11132 10011 11135
rect 10962 11132 10968 11144
rect 9999 11104 10968 11132
rect 9999 11101 10011 11104
rect 9953 11095 10011 11101
rect 10962 11092 10968 11104
rect 11020 11092 11026 11144
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11132 15715 11135
rect 15948 11132 15976 11308
rect 17586 11296 17592 11308
rect 17644 11296 17650 11348
rect 18046 11296 18052 11348
rect 18104 11296 18110 11348
rect 19794 11296 19800 11348
rect 19852 11336 19858 11348
rect 20238 11339 20296 11345
rect 20238 11336 20250 11339
rect 19852 11308 20250 11336
rect 19852 11296 19858 11308
rect 20238 11305 20250 11308
rect 20284 11305 20296 11339
rect 20238 11299 20296 11305
rect 21634 11296 21640 11348
rect 21692 11336 21698 11348
rect 21910 11336 21916 11348
rect 21692 11308 21916 11336
rect 21692 11296 21698 11308
rect 21910 11296 21916 11308
rect 21968 11336 21974 11348
rect 22097 11339 22155 11345
rect 22097 11336 22109 11339
rect 21968 11308 22109 11336
rect 21968 11296 21974 11308
rect 22097 11305 22109 11308
rect 22143 11336 22155 11339
rect 22143 11308 24716 11336
rect 22143 11305 22155 11308
rect 22097 11299 22155 11305
rect 16209 11271 16267 11277
rect 16209 11237 16221 11271
rect 16255 11237 16267 11271
rect 19518 11268 19524 11280
rect 16209 11231 16267 11237
rect 18892 11240 19524 11268
rect 15703 11104 15976 11132
rect 15703 11101 15715 11104
rect 15657 11095 15715 11101
rect 16022 11092 16028 11144
rect 16080 11092 16086 11144
rect 7098 11064 7104 11076
rect 4304 11036 5948 11064
rect 6946 11036 7104 11064
rect 4304 11024 4310 11036
rect 5920 11008 5948 11036
rect 7098 11024 7104 11036
rect 7156 11024 7162 11076
rect 7561 11067 7619 11073
rect 7561 11033 7573 11067
rect 7607 11064 7619 11067
rect 7607 11036 7696 11064
rect 7607 11033 7619 11036
rect 7561 11027 7619 11033
rect 7668 11008 7696 11036
rect 8938 11024 8944 11076
rect 8996 11064 9002 11076
rect 10689 11067 10747 11073
rect 10689 11064 10701 11067
rect 8996 11036 10701 11064
rect 8996 11024 9002 11036
rect 10689 11033 10701 11036
rect 10735 11033 10747 11067
rect 10689 11027 10747 11033
rect 13630 11024 13636 11076
rect 13688 11064 13694 11076
rect 14366 11064 14372 11076
rect 13688 11036 14372 11064
rect 13688 11024 13694 11036
rect 14366 11024 14372 11036
rect 14424 11024 14430 11076
rect 15841 11067 15899 11073
rect 15841 11033 15853 11067
rect 15887 11033 15899 11067
rect 15841 11027 15899 11033
rect 4614 10996 4620 11008
rect 4080 10968 4620 10996
rect 4614 10956 4620 10968
rect 4672 10956 4678 11008
rect 4706 10956 4712 11008
rect 4764 10996 4770 11008
rect 5077 10999 5135 11005
rect 5077 10996 5089 10999
rect 4764 10968 5089 10996
rect 4764 10956 4770 10968
rect 5077 10965 5089 10968
rect 5123 10965 5135 10999
rect 5077 10959 5135 10965
rect 5902 10956 5908 11008
rect 5960 10956 5966 11008
rect 7650 10956 7656 11008
rect 7708 10996 7714 11008
rect 12434 10996 12440 11008
rect 7708 10968 12440 10996
rect 7708 10956 7714 10968
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 15856 10996 15884 11027
rect 15930 11024 15936 11076
rect 15988 11024 15994 11076
rect 16224 11064 16252 11231
rect 16301 11203 16359 11209
rect 16301 11169 16313 11203
rect 16347 11200 16359 11203
rect 16574 11200 16580 11212
rect 16347 11172 16580 11200
rect 16347 11169 16359 11172
rect 16301 11163 16359 11169
rect 16574 11160 16580 11172
rect 16632 11160 16638 11212
rect 16942 11160 16948 11212
rect 17000 11200 17006 11212
rect 18892 11209 18920 11240
rect 19518 11228 19524 11240
rect 19576 11228 19582 11280
rect 24688 11277 24716 11308
rect 26694 11296 26700 11348
rect 26752 11296 26758 11348
rect 22465 11271 22523 11277
rect 22465 11237 22477 11271
rect 22511 11268 22523 11271
rect 24673 11271 24731 11277
rect 22511 11240 23704 11268
rect 22511 11237 22523 11240
rect 22465 11231 22523 11237
rect 18877 11203 18935 11209
rect 18877 11200 18889 11203
rect 17000 11172 18889 11200
rect 17000 11160 17006 11172
rect 18877 11169 18889 11172
rect 18923 11169 18935 11203
rect 19981 11203 20039 11209
rect 19981 11200 19993 11203
rect 18877 11163 18935 11169
rect 19260 11172 19993 11200
rect 19260 11144 19288 11172
rect 19981 11169 19993 11172
rect 20027 11200 20039 11203
rect 22480 11200 22508 11231
rect 23676 11212 23704 11240
rect 24673 11237 24685 11271
rect 24719 11237 24731 11271
rect 24673 11231 24731 11237
rect 20027 11172 21773 11200
rect 20027 11169 20039 11172
rect 19981 11163 20039 11169
rect 17862 11132 17868 11144
rect 17710 11104 17868 11132
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 18414 11092 18420 11144
rect 18472 11132 18478 11144
rect 18509 11135 18567 11141
rect 18509 11132 18521 11135
rect 18472 11104 18521 11132
rect 18472 11092 18478 11104
rect 18509 11101 18521 11104
rect 18555 11101 18567 11135
rect 18509 11095 18567 11101
rect 18690 11092 18696 11144
rect 18748 11092 18754 11144
rect 19242 11092 19248 11144
rect 19300 11092 19306 11144
rect 19426 11092 19432 11144
rect 19484 11092 19490 11144
rect 19610 11092 19616 11144
rect 19668 11132 19674 11144
rect 19705 11135 19763 11141
rect 19705 11132 19717 11135
rect 19668 11104 19717 11132
rect 19668 11092 19674 11104
rect 19705 11101 19717 11104
rect 19751 11101 19763 11135
rect 21542 11132 21548 11144
rect 21390 11104 21548 11132
rect 19705 11095 19763 11101
rect 21542 11092 21548 11104
rect 21600 11092 21606 11144
rect 16577 11067 16635 11073
rect 16577 11064 16589 11067
rect 16224 11036 16589 11064
rect 16577 11033 16589 11036
rect 16623 11033 16635 11067
rect 16577 11027 16635 11033
rect 16666 11024 16672 11076
rect 16724 11064 16730 11076
rect 16850 11064 16856 11076
rect 16724 11036 16856 11064
rect 16724 11024 16730 11036
rect 16850 11024 16856 11036
rect 16908 11024 16914 11076
rect 18708 11064 18736 11092
rect 19978 11064 19984 11076
rect 18708 11036 19984 11064
rect 19978 11024 19984 11036
rect 20036 11024 20042 11076
rect 16684 10996 16712 11024
rect 15856 10968 16712 10996
rect 17862 10956 17868 11008
rect 17920 10996 17926 11008
rect 19334 10996 19340 11008
rect 17920 10968 19340 10996
rect 17920 10956 17926 10968
rect 19334 10956 19340 10968
rect 19392 10996 19398 11008
rect 20530 10996 20536 11008
rect 19392 10968 20536 10996
rect 19392 10956 19398 10968
rect 20530 10956 20536 10968
rect 20588 10956 20594 11008
rect 21745 10996 21773 11172
rect 22158 11172 22508 11200
rect 22158 11144 22186 11172
rect 23658 11160 23664 11212
rect 23716 11160 23722 11212
rect 24394 11160 24400 11212
rect 24452 11200 24458 11212
rect 26712 11200 26740 11296
rect 26881 11203 26939 11209
rect 26881 11200 26893 11203
rect 24452 11172 26372 11200
rect 26712 11172 26893 11200
rect 24452 11160 24458 11172
rect 26344 11144 26372 11172
rect 26881 11169 26893 11172
rect 26927 11169 26939 11203
rect 26881 11163 26939 11169
rect 22094 11092 22100 11144
rect 22152 11135 22186 11144
rect 22167 11104 22186 11135
rect 22281 11135 22339 11141
rect 22167 11101 22179 11104
rect 22152 11095 22179 11101
rect 22281 11101 22293 11135
rect 22327 11101 22339 11135
rect 22281 11095 22339 11101
rect 22373 11135 22431 11141
rect 22373 11101 22385 11135
rect 22419 11132 22431 11135
rect 22554 11132 22560 11144
rect 22419 11104 22560 11132
rect 22419 11101 22431 11104
rect 22373 11095 22431 11101
rect 22152 11092 22158 11095
rect 22002 11024 22008 11076
rect 22060 11064 22066 11076
rect 22296 11064 22324 11095
rect 22554 11092 22560 11104
rect 22612 11092 22618 11144
rect 22649 11135 22707 11141
rect 22649 11101 22661 11135
rect 22695 11132 22707 11135
rect 23290 11132 23296 11144
rect 22695 11104 23296 11132
rect 22695 11101 22707 11104
rect 22649 11095 22707 11101
rect 22664 11064 22692 11095
rect 23290 11092 23296 11104
rect 23348 11092 23354 11144
rect 23385 11135 23443 11141
rect 23385 11101 23397 11135
rect 23431 11132 23443 11135
rect 23431 11104 24900 11132
rect 23431 11101 23443 11104
rect 23385 11095 23443 11101
rect 22060 11036 22692 11064
rect 22060 11024 22066 11036
rect 22738 11024 22744 11076
rect 22796 11024 22802 11076
rect 22830 11024 22836 11076
rect 22888 11064 22894 11076
rect 23109 11067 23167 11073
rect 23109 11064 23121 11067
rect 22888 11036 23121 11064
rect 22888 11024 22894 11036
rect 23109 11033 23121 11036
rect 23155 11064 23167 11067
rect 23566 11064 23572 11076
rect 23155 11036 23572 11064
rect 23155 11033 23167 11036
rect 23109 11027 23167 11033
rect 23566 11024 23572 11036
rect 23624 11024 23630 11076
rect 24029 11067 24087 11073
rect 24029 11033 24041 11067
rect 24075 11033 24087 11067
rect 24029 11027 24087 11033
rect 22756 10996 22784 11024
rect 21745 10968 22784 10996
rect 23474 10956 23480 11008
rect 23532 10996 23538 11008
rect 24044 10996 24072 11027
rect 24118 11024 24124 11076
rect 24176 11064 24182 11076
rect 24397 11067 24455 11073
rect 24397 11064 24409 11067
rect 24176 11036 24409 11064
rect 24176 11024 24182 11036
rect 24397 11033 24409 11036
rect 24443 11033 24455 11067
rect 24397 11027 24455 11033
rect 24762 11024 24768 11076
rect 24820 11024 24826 11076
rect 24780 10996 24808 11024
rect 24872 11005 24900 11104
rect 24946 11092 24952 11144
rect 25004 11092 25010 11144
rect 26326 11092 26332 11144
rect 26384 11132 26390 11144
rect 27062 11132 27068 11144
rect 26384 11104 27068 11132
rect 26384 11092 26390 11104
rect 27062 11092 27068 11104
rect 27120 11092 27126 11144
rect 28718 11092 28724 11144
rect 28776 11092 28782 11144
rect 25222 11024 25228 11076
rect 25280 11024 25286 11076
rect 26620 11036 27568 11064
rect 23532 10968 24808 10996
rect 24857 10999 24915 11005
rect 23532 10956 23538 10968
rect 24857 10965 24869 10999
rect 24903 10965 24915 10999
rect 24857 10959 24915 10965
rect 26050 10956 26056 11008
rect 26108 10996 26114 11008
rect 26620 10996 26648 11036
rect 27540 11005 27568 11036
rect 29086 11024 29092 11076
rect 29144 11024 29150 11076
rect 26108 10968 26648 10996
rect 27525 10999 27583 11005
rect 26108 10956 26114 10968
rect 27525 10965 27537 10999
rect 27571 10965 27583 10999
rect 27525 10959 27583 10965
rect 1104 10906 29595 10928
rect 1104 10854 8032 10906
rect 8084 10854 8096 10906
rect 8148 10854 8160 10906
rect 8212 10854 8224 10906
rect 8276 10854 8288 10906
rect 8340 10854 15115 10906
rect 15167 10854 15179 10906
rect 15231 10854 15243 10906
rect 15295 10854 15307 10906
rect 15359 10854 15371 10906
rect 15423 10854 22198 10906
rect 22250 10854 22262 10906
rect 22314 10854 22326 10906
rect 22378 10854 22390 10906
rect 22442 10854 22454 10906
rect 22506 10854 29281 10906
rect 29333 10854 29345 10906
rect 29397 10854 29409 10906
rect 29461 10854 29473 10906
rect 29525 10854 29537 10906
rect 29589 10854 29595 10906
rect 1104 10832 29595 10854
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 5169 10795 5227 10801
rect 5169 10792 5181 10795
rect 4212 10764 5181 10792
rect 4212 10752 4218 10764
rect 5169 10761 5181 10764
rect 5215 10761 5227 10795
rect 5169 10755 5227 10761
rect 5902 10752 5908 10804
rect 5960 10752 5966 10804
rect 5997 10795 6055 10801
rect 5997 10761 6009 10795
rect 6043 10792 6055 10795
rect 6454 10792 6460 10804
rect 6043 10764 6460 10792
rect 6043 10761 6055 10764
rect 5997 10755 6055 10761
rect 6454 10752 6460 10764
rect 6512 10752 6518 10804
rect 6825 10795 6883 10801
rect 6825 10761 6837 10795
rect 6871 10792 6883 10795
rect 9677 10795 9735 10801
rect 6871 10764 9628 10792
rect 6871 10761 6883 10764
rect 6825 10755 6883 10761
rect 3973 10727 4031 10733
rect 3973 10693 3985 10727
rect 4019 10724 4031 10727
rect 4798 10724 4804 10736
rect 4019 10696 4804 10724
rect 4019 10693 4031 10696
rect 3973 10687 4031 10693
rect 4798 10684 4804 10696
rect 4856 10684 4862 10736
rect 4893 10727 4951 10733
rect 4893 10693 4905 10727
rect 4939 10724 4951 10727
rect 4939 10696 5212 10724
rect 4939 10693 4951 10696
rect 4893 10687 4951 10693
rect 3789 10659 3847 10665
rect 3789 10625 3801 10659
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 4065 10659 4123 10665
rect 4065 10625 4077 10659
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10656 4215 10659
rect 4617 10659 4675 10665
rect 4203 10628 4568 10656
rect 4203 10625 4215 10628
rect 4157 10619 4215 10625
rect 3804 10452 3832 10619
rect 3970 10548 3976 10600
rect 4028 10588 4034 10600
rect 4080 10588 4108 10619
rect 4028 10560 4108 10588
rect 4028 10548 4034 10560
rect 4062 10452 4068 10464
rect 3804 10424 4068 10452
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 4154 10412 4160 10464
rect 4212 10452 4218 10464
rect 4341 10455 4399 10461
rect 4341 10452 4353 10455
rect 4212 10424 4353 10452
rect 4212 10412 4218 10424
rect 4341 10421 4353 10424
rect 4387 10421 4399 10455
rect 4540 10452 4568 10628
rect 4617 10625 4629 10659
rect 4663 10656 4675 10659
rect 4706 10656 4712 10668
rect 4663 10628 4712 10656
rect 4663 10625 4675 10628
rect 4617 10619 4675 10625
rect 4706 10616 4712 10628
rect 4764 10616 4770 10668
rect 4908 10656 4936 10687
rect 4816 10628 4936 10656
rect 4985 10659 5043 10665
rect 4614 10480 4620 10532
rect 4672 10520 4678 10532
rect 4816 10520 4844 10628
rect 4985 10625 4997 10659
rect 5031 10625 5043 10659
rect 5184 10656 5212 10696
rect 5350 10684 5356 10736
rect 5408 10724 5414 10736
rect 5445 10727 5503 10733
rect 5445 10724 5457 10727
rect 5408 10696 5457 10724
rect 5408 10684 5414 10696
rect 5445 10693 5457 10696
rect 5491 10693 5503 10727
rect 5445 10687 5503 10693
rect 5534 10684 5540 10736
rect 5592 10724 5598 10736
rect 6365 10727 6423 10733
rect 6365 10724 6377 10727
rect 5592 10696 6377 10724
rect 5592 10684 5598 10696
rect 6365 10693 6377 10696
rect 6411 10693 6423 10727
rect 7650 10724 7656 10736
rect 6365 10687 6423 10693
rect 6472 10696 7656 10724
rect 6472 10656 6500 10696
rect 7650 10684 7656 10696
rect 7708 10684 7714 10736
rect 9600 10724 9628 10764
rect 9677 10761 9689 10795
rect 9723 10792 9735 10795
rect 9766 10792 9772 10804
rect 9723 10764 9772 10792
rect 9723 10761 9735 10764
rect 9677 10755 9735 10761
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10008 10764 11192 10792
rect 10008 10752 10014 10764
rect 11164 10736 11192 10764
rect 14090 10752 14096 10804
rect 14148 10792 14154 10804
rect 14461 10795 14519 10801
rect 14461 10792 14473 10795
rect 14148 10764 14473 10792
rect 14148 10752 14154 10764
rect 14461 10761 14473 10764
rect 14507 10761 14519 10795
rect 14461 10755 14519 10761
rect 14553 10795 14611 10801
rect 14553 10761 14565 10795
rect 14599 10792 14611 10795
rect 14734 10792 14740 10804
rect 14599 10764 14740 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 14734 10752 14740 10764
rect 14792 10752 14798 10804
rect 17865 10795 17923 10801
rect 17865 10761 17877 10795
rect 17911 10792 17923 10795
rect 18506 10792 18512 10804
rect 17911 10764 18512 10792
rect 17911 10761 17923 10764
rect 17865 10755 17923 10761
rect 18506 10752 18512 10764
rect 18564 10792 18570 10804
rect 19981 10795 20039 10801
rect 19981 10792 19993 10795
rect 18564 10764 19993 10792
rect 18564 10752 18570 10764
rect 19981 10761 19993 10764
rect 20027 10761 20039 10795
rect 19981 10755 20039 10761
rect 21450 10752 21456 10804
rect 21508 10752 21514 10804
rect 22002 10752 22008 10804
rect 22060 10752 22066 10804
rect 22741 10795 22799 10801
rect 22741 10761 22753 10795
rect 22787 10792 22799 10795
rect 23014 10792 23020 10804
rect 22787 10764 23020 10792
rect 22787 10761 22799 10764
rect 22741 10755 22799 10761
rect 23014 10752 23020 10764
rect 23072 10752 23078 10804
rect 23842 10792 23848 10804
rect 23124 10764 23848 10792
rect 9600 10696 10456 10724
rect 5184 10628 6500 10656
rect 6641 10659 6699 10665
rect 4985 10619 5043 10625
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 7190 10656 7196 10668
rect 6687 10628 7196 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 5000 10588 5028 10619
rect 7190 10616 7196 10628
rect 7248 10616 7254 10668
rect 9766 10616 9772 10668
rect 9824 10656 9830 10668
rect 9861 10659 9919 10665
rect 9861 10656 9873 10659
rect 9824 10628 9873 10656
rect 9824 10616 9830 10628
rect 9861 10625 9873 10628
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 5258 10588 5264 10600
rect 4672 10492 4844 10520
rect 4904 10560 5264 10588
rect 4672 10480 4678 10492
rect 4904 10452 4932 10560
rect 5258 10548 5264 10560
rect 5316 10548 5322 10600
rect 6181 10591 6239 10597
rect 6181 10557 6193 10591
rect 6227 10588 6239 10591
rect 6457 10591 6515 10597
rect 6457 10588 6469 10591
rect 6227 10560 6469 10588
rect 6227 10557 6239 10560
rect 6181 10551 6239 10557
rect 6457 10557 6469 10560
rect 6503 10557 6515 10591
rect 7006 10588 7012 10600
rect 6457 10551 6515 10557
rect 6564 10560 7012 10588
rect 4982 10480 4988 10532
rect 5040 10520 5046 10532
rect 5445 10523 5503 10529
rect 5445 10520 5457 10523
rect 5040 10492 5457 10520
rect 5040 10480 5046 10492
rect 5445 10489 5457 10492
rect 5491 10489 5503 10523
rect 5445 10483 5503 10489
rect 6564 10461 6592 10560
rect 7006 10548 7012 10560
rect 7064 10548 7070 10600
rect 4540 10424 4932 10452
rect 6549 10455 6607 10461
rect 4341 10415 4399 10421
rect 6549 10421 6561 10455
rect 6595 10421 6607 10455
rect 9968 10452 9996 10619
rect 10134 10616 10140 10668
rect 10192 10616 10198 10668
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10625 10287 10659
rect 10229 10619 10287 10625
rect 10244 10520 10272 10619
rect 10318 10616 10324 10668
rect 10376 10665 10382 10668
rect 10376 10659 10397 10665
rect 10385 10625 10397 10659
rect 10428 10656 10456 10696
rect 10502 10684 10508 10736
rect 10560 10724 10566 10736
rect 10560 10696 10603 10724
rect 10560 10684 10566 10696
rect 11146 10684 11152 10736
rect 11204 10684 11210 10736
rect 17129 10727 17187 10733
rect 17129 10724 17141 10727
rect 13372 10696 17141 10724
rect 13372 10656 13400 10696
rect 17129 10693 17141 10696
rect 17175 10693 17187 10727
rect 17129 10687 17187 10693
rect 17221 10727 17279 10733
rect 17221 10693 17233 10727
rect 17267 10724 17279 10727
rect 19886 10724 19892 10736
rect 17267 10696 19892 10724
rect 17267 10693 17279 10696
rect 17221 10687 17279 10693
rect 19886 10684 19892 10696
rect 19944 10684 19950 10736
rect 20070 10724 20076 10736
rect 19996 10696 20076 10724
rect 10428 10628 13400 10656
rect 10376 10619 10397 10625
rect 10376 10616 10382 10619
rect 13630 10616 13636 10668
rect 13688 10616 13694 10668
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10656 13783 10659
rect 14274 10656 14280 10668
rect 13771 10628 14280 10656
rect 13771 10625 13783 10628
rect 13725 10619 13783 10625
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 14366 10616 14372 10668
rect 14424 10616 14430 10668
rect 16301 10659 16359 10665
rect 16301 10625 16313 10659
rect 16347 10656 16359 10659
rect 16390 10656 16396 10668
rect 16347 10628 16396 10656
rect 16347 10625 16359 10628
rect 16301 10619 16359 10625
rect 16390 10616 16396 10628
rect 16448 10616 16454 10668
rect 16485 10659 16543 10665
rect 16485 10625 16497 10659
rect 16531 10656 16543 10659
rect 16853 10659 16911 10665
rect 16853 10656 16865 10659
rect 16531 10628 16865 10656
rect 16531 10625 16543 10628
rect 16485 10619 16543 10625
rect 16853 10625 16865 10628
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 17001 10659 17059 10665
rect 17001 10625 17013 10659
rect 17047 10656 17059 10659
rect 17047 10625 17080 10656
rect 17001 10619 17080 10625
rect 10502 10548 10508 10600
rect 10560 10588 10566 10600
rect 11422 10588 11428 10600
rect 10560 10560 11428 10588
rect 10560 10548 10566 10560
rect 11422 10548 11428 10560
rect 11480 10548 11486 10600
rect 12434 10548 12440 10600
rect 12492 10548 12498 10600
rect 13648 10588 13676 10616
rect 13817 10591 13875 10597
rect 13817 10588 13829 10591
rect 13648 10560 13829 10588
rect 13817 10557 13829 10560
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 13909 10591 13967 10597
rect 13909 10557 13921 10591
rect 13955 10557 13967 10591
rect 13909 10551 13967 10557
rect 14001 10591 14059 10597
rect 14001 10557 14013 10591
rect 14047 10588 14059 10591
rect 14090 10588 14096 10600
rect 14047 10560 14096 10588
rect 14047 10557 14059 10560
rect 14001 10551 14059 10557
rect 10594 10520 10600 10532
rect 10244 10492 10600 10520
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 12452 10520 12480 10548
rect 13924 10520 13952 10551
rect 14090 10548 14096 10560
rect 14148 10548 14154 10600
rect 15930 10588 15936 10600
rect 14200 10560 15936 10588
rect 14200 10529 14228 10560
rect 15930 10548 15936 10560
rect 15988 10588 15994 10600
rect 16117 10591 16175 10597
rect 16117 10588 16129 10591
rect 15988 10560 16129 10588
rect 15988 10548 15994 10560
rect 16117 10557 16129 10560
rect 16163 10557 16175 10591
rect 17052 10588 17080 10619
rect 17310 10616 17316 10668
rect 17368 10665 17374 10668
rect 17368 10656 17376 10665
rect 17678 10656 17684 10668
rect 17368 10628 17684 10656
rect 17368 10619 17376 10628
rect 17368 10616 17374 10619
rect 17678 10616 17684 10628
rect 17736 10616 17742 10668
rect 17862 10616 17868 10668
rect 17920 10656 17926 10668
rect 17920 10628 17962 10656
rect 17920 10616 17926 10628
rect 18046 10616 18052 10668
rect 18104 10656 18110 10668
rect 18233 10659 18291 10665
rect 18233 10656 18245 10659
rect 18104 10628 18245 10656
rect 18104 10616 18110 10628
rect 18233 10625 18245 10628
rect 18279 10625 18291 10659
rect 18233 10619 18291 10625
rect 18322 10616 18328 10668
rect 18380 10616 18386 10668
rect 18601 10659 18659 10665
rect 18601 10625 18613 10659
rect 18647 10656 18659 10659
rect 18690 10656 18696 10668
rect 18647 10628 18696 10656
rect 18647 10625 18659 10628
rect 18601 10619 18659 10625
rect 18690 10616 18696 10628
rect 18748 10616 18754 10668
rect 18793 10659 18851 10665
rect 18793 10625 18805 10659
rect 18839 10656 18851 10659
rect 18839 10628 19104 10656
rect 18839 10625 18851 10628
rect 18793 10619 18851 10625
rect 19076 10588 19104 10628
rect 19150 10616 19156 10668
rect 19208 10616 19214 10668
rect 19245 10659 19303 10665
rect 19245 10625 19257 10659
rect 19291 10656 19303 10659
rect 19996 10656 20024 10696
rect 20070 10684 20076 10696
rect 20128 10724 20134 10736
rect 22020 10724 22048 10752
rect 23124 10733 23152 10764
rect 23842 10752 23848 10764
rect 23900 10752 23906 10804
rect 25222 10752 25228 10804
rect 25280 10792 25286 10804
rect 25409 10795 25467 10801
rect 25409 10792 25421 10795
rect 25280 10764 25421 10792
rect 25280 10752 25286 10764
rect 25409 10761 25421 10764
rect 25455 10761 25467 10795
rect 25409 10755 25467 10761
rect 26145 10795 26203 10801
rect 26145 10761 26157 10795
rect 26191 10761 26203 10795
rect 26145 10755 26203 10761
rect 23109 10727 23167 10733
rect 20128 10696 22600 10724
rect 20128 10684 20134 10696
rect 19291 10628 20024 10656
rect 20165 10659 20223 10665
rect 19291 10625 19303 10628
rect 19245 10619 19303 10625
rect 20165 10625 20177 10659
rect 20211 10656 20223 10659
rect 20254 10656 20260 10668
rect 20211 10628 20260 10656
rect 20211 10625 20223 10628
rect 20165 10619 20223 10625
rect 20254 10616 20260 10628
rect 20312 10616 20318 10668
rect 20640 10665 20668 10696
rect 20625 10659 20683 10665
rect 20625 10625 20637 10659
rect 20671 10625 20683 10659
rect 20625 10619 20683 10625
rect 20901 10659 20959 10665
rect 20901 10625 20913 10659
rect 20947 10656 20959 10659
rect 22094 10656 22100 10668
rect 20947 10628 22100 10656
rect 20947 10625 20959 10628
rect 20901 10619 20959 10625
rect 19705 10591 19763 10597
rect 19705 10588 19717 10591
rect 17052 10560 17724 10588
rect 19076 10560 19717 10588
rect 16117 10551 16175 10557
rect 14185 10523 14243 10529
rect 14185 10520 14197 10523
rect 12452 10492 13768 10520
rect 10226 10452 10232 10464
rect 9968 10424 10232 10452
rect 6549 10415 6607 10421
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 10689 10455 10747 10461
rect 10689 10452 10701 10455
rect 10560 10424 10701 10452
rect 10560 10412 10566 10424
rect 10689 10421 10701 10424
rect 10735 10421 10747 10455
rect 10689 10415 10747 10421
rect 13538 10412 13544 10464
rect 13596 10412 13602 10464
rect 13740 10452 13768 10492
rect 13924 10492 14197 10520
rect 13924 10452 13952 10492
rect 14185 10489 14197 10492
rect 14231 10489 14243 10523
rect 14185 10483 14243 10489
rect 15286 10480 15292 10532
rect 15344 10520 15350 10532
rect 17696 10529 17724 10560
rect 19705 10557 19717 10560
rect 19751 10588 19763 10591
rect 20346 10588 20352 10600
rect 19751 10560 20352 10588
rect 19751 10557 19763 10560
rect 19705 10551 19763 10557
rect 20346 10548 20352 10560
rect 20404 10588 20410 10600
rect 20916 10588 20944 10619
rect 22094 10616 22100 10628
rect 22152 10616 22158 10668
rect 22572 10665 22600 10696
rect 23109 10693 23121 10727
rect 23155 10693 23167 10727
rect 24394 10724 24400 10736
rect 24334 10696 24400 10724
rect 23109 10687 23167 10693
rect 24394 10684 24400 10696
rect 24452 10684 24458 10736
rect 26050 10684 26056 10736
rect 26108 10684 26114 10736
rect 22557 10659 22615 10665
rect 22557 10625 22569 10659
rect 22603 10625 22615 10659
rect 22557 10619 22615 10625
rect 22833 10659 22891 10665
rect 22833 10625 22845 10659
rect 22879 10625 22891 10659
rect 22833 10619 22891 10625
rect 25685 10659 25743 10665
rect 25685 10625 25697 10659
rect 25731 10656 25743 10659
rect 26160 10656 26188 10755
rect 26234 10684 26240 10736
rect 26292 10684 26298 10736
rect 25731 10628 26188 10656
rect 26252 10656 26280 10684
rect 26329 10659 26387 10665
rect 26329 10656 26341 10659
rect 26252 10628 26341 10656
rect 25731 10625 25743 10628
rect 25685 10619 25743 10625
rect 26329 10625 26341 10628
rect 26375 10625 26387 10659
rect 26329 10619 26387 10625
rect 20404 10560 20944 10588
rect 22373 10591 22431 10597
rect 20404 10548 20410 10560
rect 22373 10557 22385 10591
rect 22419 10588 22431 10591
rect 22646 10588 22652 10600
rect 22419 10560 22652 10588
rect 22419 10557 22431 10560
rect 22373 10551 22431 10557
rect 17681 10523 17739 10529
rect 15344 10492 17632 10520
rect 15344 10480 15350 10492
rect 13740 10424 13952 10452
rect 14458 10412 14464 10464
rect 14516 10452 14522 10464
rect 14737 10455 14795 10461
rect 14737 10452 14749 10455
rect 14516 10424 14749 10452
rect 14516 10412 14522 10424
rect 14737 10421 14749 10424
rect 14783 10421 14795 10455
rect 14737 10415 14795 10421
rect 15654 10412 15660 10464
rect 15712 10452 15718 10464
rect 16390 10452 16396 10464
rect 15712 10424 16396 10452
rect 15712 10412 15718 10424
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 16942 10412 16948 10464
rect 17000 10452 17006 10464
rect 17497 10455 17555 10461
rect 17497 10452 17509 10455
rect 17000 10424 17509 10452
rect 17000 10412 17006 10424
rect 17497 10421 17509 10424
rect 17543 10421 17555 10455
rect 17604 10452 17632 10492
rect 17681 10489 17693 10523
rect 17727 10489 17739 10523
rect 17681 10483 17739 10489
rect 17785 10492 22094 10520
rect 17785 10452 17813 10492
rect 22066 10464 22094 10492
rect 22388 10464 22416 10551
rect 22646 10548 22652 10560
rect 22704 10548 22710 10600
rect 22848 10588 22876 10619
rect 26418 10616 26424 10668
rect 26476 10616 26482 10668
rect 26510 10616 26516 10668
rect 26568 10616 26574 10668
rect 26697 10659 26755 10665
rect 26697 10625 26709 10659
rect 26743 10625 26755 10659
rect 26697 10619 26755 10625
rect 26789 10659 26847 10665
rect 26789 10625 26801 10659
rect 26835 10625 26847 10659
rect 26789 10619 26847 10625
rect 22848 10560 22968 10588
rect 22830 10480 22836 10532
rect 22888 10480 22894 10532
rect 17604 10424 17813 10452
rect 17497 10415 17555 10421
rect 18046 10412 18052 10464
rect 18104 10452 18110 10464
rect 18969 10455 19027 10461
rect 18969 10452 18981 10455
rect 18104 10424 18981 10452
rect 18104 10412 18110 10424
rect 18969 10421 18981 10424
rect 19015 10421 19027 10455
rect 18969 10415 19027 10421
rect 19058 10412 19064 10464
rect 19116 10452 19122 10464
rect 19613 10455 19671 10461
rect 19613 10452 19625 10455
rect 19116 10424 19625 10452
rect 19116 10412 19122 10424
rect 19613 10421 19625 10424
rect 19659 10452 19671 10455
rect 20254 10452 20260 10464
rect 19659 10424 20260 10452
rect 19659 10421 19671 10424
rect 19613 10415 19671 10421
rect 20254 10412 20260 10424
rect 20312 10412 20318 10464
rect 22066 10424 22100 10464
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 22370 10412 22376 10464
rect 22428 10412 22434 10464
rect 22554 10412 22560 10464
rect 22612 10412 22618 10464
rect 22646 10412 22652 10464
rect 22704 10452 22710 10464
rect 22848 10452 22876 10480
rect 22940 10464 22968 10560
rect 23658 10548 23664 10600
rect 23716 10588 23722 10600
rect 24857 10591 24915 10597
rect 24857 10588 24869 10591
rect 23716 10560 24869 10588
rect 23716 10548 23722 10560
rect 24857 10557 24869 10560
rect 24903 10557 24915 10591
rect 24857 10551 24915 10557
rect 25590 10548 25596 10600
rect 25648 10548 25654 10600
rect 25866 10548 25872 10600
rect 25924 10588 25930 10600
rect 25961 10591 26019 10597
rect 25961 10588 25973 10591
rect 25924 10560 25973 10588
rect 25924 10548 25930 10560
rect 25961 10557 25973 10560
rect 26007 10588 26019 10591
rect 26142 10588 26148 10600
rect 26007 10560 26148 10588
rect 26007 10557 26019 10560
rect 25961 10551 26019 10557
rect 26142 10548 26148 10560
rect 26200 10588 26206 10600
rect 26712 10588 26740 10619
rect 26200 10560 26740 10588
rect 26200 10548 26206 10560
rect 24762 10480 24768 10532
rect 24820 10520 24826 10532
rect 26804 10520 26832 10619
rect 24820 10492 26832 10520
rect 24820 10480 24826 10492
rect 22704 10424 22876 10452
rect 22704 10412 22710 10424
rect 22922 10412 22928 10464
rect 22980 10452 22986 10464
rect 24946 10452 24952 10464
rect 22980 10424 24952 10452
rect 22980 10412 22986 10424
rect 24946 10412 24952 10424
rect 25004 10412 25010 10464
rect 1104 10362 29440 10384
rect 1104 10310 4491 10362
rect 4543 10310 4555 10362
rect 4607 10310 4619 10362
rect 4671 10310 4683 10362
rect 4735 10310 4747 10362
rect 4799 10310 11574 10362
rect 11626 10310 11638 10362
rect 11690 10310 11702 10362
rect 11754 10310 11766 10362
rect 11818 10310 11830 10362
rect 11882 10310 18657 10362
rect 18709 10310 18721 10362
rect 18773 10310 18785 10362
rect 18837 10310 18849 10362
rect 18901 10310 18913 10362
rect 18965 10310 25740 10362
rect 25792 10310 25804 10362
rect 25856 10310 25868 10362
rect 25920 10310 25932 10362
rect 25984 10310 25996 10362
rect 26048 10310 29440 10362
rect 1104 10288 29440 10310
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 4709 10251 4767 10257
rect 4709 10248 4721 10251
rect 4120 10220 4721 10248
rect 4120 10208 4126 10220
rect 4709 10217 4721 10220
rect 4755 10217 4767 10251
rect 4709 10211 4767 10217
rect 9766 10208 9772 10260
rect 9824 10208 9830 10260
rect 10134 10208 10140 10260
rect 10192 10248 10198 10260
rect 10597 10251 10655 10257
rect 10597 10248 10609 10251
rect 10192 10220 10609 10248
rect 10192 10208 10198 10220
rect 10597 10217 10609 10220
rect 10643 10217 10655 10251
rect 10597 10211 10655 10217
rect 12161 10251 12219 10257
rect 12161 10217 12173 10251
rect 12207 10248 12219 10251
rect 12342 10248 12348 10260
rect 12207 10220 12348 10248
rect 12207 10217 12219 10220
rect 12161 10211 12219 10217
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 13538 10208 13544 10260
rect 13596 10208 13602 10260
rect 13725 10251 13783 10257
rect 13725 10217 13737 10251
rect 13771 10248 13783 10251
rect 13906 10248 13912 10260
rect 13771 10220 13912 10248
rect 13771 10217 13783 10220
rect 13725 10211 13783 10217
rect 13906 10208 13912 10220
rect 13964 10208 13970 10260
rect 18046 10248 18052 10260
rect 14016 10220 18052 10248
rect 3970 10140 3976 10192
rect 4028 10180 4034 10192
rect 5258 10180 5264 10192
rect 4028 10152 5264 10180
rect 4028 10140 4034 10152
rect 5258 10140 5264 10152
rect 5316 10140 5322 10192
rect 9784 10180 9812 10208
rect 10962 10180 10968 10192
rect 9416 10152 10968 10180
rect 9416 10112 9444 10152
rect 10962 10140 10968 10152
rect 11020 10180 11026 10192
rect 14016 10180 14044 10220
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 20530 10208 20536 10260
rect 20588 10208 20594 10260
rect 22094 10208 22100 10260
rect 22152 10248 22158 10260
rect 22646 10248 22652 10260
rect 22152 10220 22652 10248
rect 22152 10208 22158 10220
rect 22646 10208 22652 10220
rect 22704 10208 22710 10260
rect 22833 10251 22891 10257
rect 22833 10217 22845 10251
rect 22879 10217 22891 10251
rect 22833 10211 22891 10217
rect 11020 10152 14044 10180
rect 16500 10152 16712 10180
rect 11020 10140 11026 10152
rect 9493 10115 9551 10121
rect 9493 10112 9505 10115
rect 9416 10084 9505 10112
rect 9493 10081 9505 10084
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 9582 10072 9588 10124
rect 9640 10072 9646 10124
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 9824 10084 10088 10112
rect 9824 10072 9830 10084
rect 4062 10004 4068 10056
rect 4120 10004 4126 10056
rect 9861 10047 9919 10053
rect 9861 10013 9873 10047
rect 9907 10044 9919 10047
rect 9950 10044 9956 10056
rect 9907 10016 9956 10044
rect 9907 10013 9919 10016
rect 9861 10007 9919 10013
rect 9950 10004 9956 10016
rect 10008 10004 10014 10056
rect 10060 10053 10088 10084
rect 10226 10072 10232 10124
rect 10284 10112 10290 10124
rect 11333 10115 11391 10121
rect 11333 10112 11345 10115
rect 10284 10084 11345 10112
rect 10284 10072 10290 10084
rect 11333 10081 11345 10084
rect 11379 10081 11391 10115
rect 16500 10112 16528 10152
rect 11333 10075 11391 10081
rect 12360 10084 16528 10112
rect 10045 10047 10103 10053
rect 10045 10013 10057 10047
rect 10091 10013 10103 10047
rect 10045 10007 10103 10013
rect 10137 10047 10195 10053
rect 10137 10013 10149 10047
rect 10183 10044 10195 10047
rect 10318 10044 10324 10056
rect 10183 10016 10324 10044
rect 10183 10013 10195 10016
rect 10137 10007 10195 10013
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 10413 10047 10471 10053
rect 10413 10013 10425 10047
rect 10459 10044 10471 10047
rect 10778 10044 10784 10056
rect 10459 10016 10784 10044
rect 10459 10013 10471 10016
rect 10413 10007 10471 10013
rect 10778 10004 10784 10016
rect 10836 10004 10842 10056
rect 10873 10047 10931 10053
rect 10873 10013 10885 10047
rect 10919 10044 10931 10047
rect 10962 10044 10968 10056
rect 10919 10016 10968 10044
rect 10919 10013 10931 10016
rect 10873 10007 10931 10013
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11149 10047 11207 10053
rect 11149 10044 11161 10047
rect 11112 10016 11161 10044
rect 11112 10004 11118 10016
rect 11149 10013 11161 10016
rect 11195 10013 11207 10047
rect 11149 10007 11207 10013
rect 11238 10004 11244 10056
rect 11296 10004 11302 10056
rect 11422 10004 11428 10056
rect 11480 10004 11486 10056
rect 11701 10047 11759 10053
rect 11701 10013 11713 10047
rect 11747 10044 11759 10047
rect 12360 10044 12388 10084
rect 12820 10053 12848 10084
rect 16574 10072 16580 10124
rect 16632 10072 16638 10124
rect 16684 10112 16712 10152
rect 18414 10140 18420 10192
rect 18472 10140 18478 10192
rect 20349 10183 20407 10189
rect 20349 10180 20361 10183
rect 19812 10152 20361 10180
rect 18432 10112 18460 10140
rect 19150 10112 19156 10124
rect 16684 10084 19156 10112
rect 19150 10072 19156 10084
rect 19208 10112 19214 10124
rect 19812 10112 19840 10152
rect 20349 10149 20361 10152
rect 20395 10180 20407 10183
rect 22370 10180 22376 10192
rect 20395 10152 22376 10180
rect 20395 10149 20407 10152
rect 20349 10143 20407 10149
rect 22370 10140 22376 10152
rect 22428 10140 22434 10192
rect 22554 10140 22560 10192
rect 22612 10180 22618 10192
rect 22848 10180 22876 10211
rect 23106 10208 23112 10260
rect 23164 10208 23170 10260
rect 23198 10208 23204 10260
rect 23256 10248 23262 10260
rect 23293 10251 23351 10257
rect 23293 10248 23305 10251
rect 23256 10220 23305 10248
rect 23256 10208 23262 10220
rect 23293 10217 23305 10220
rect 23339 10217 23351 10251
rect 23293 10211 23351 10217
rect 25590 10208 25596 10260
rect 25648 10248 25654 10260
rect 25869 10251 25927 10257
rect 25869 10248 25881 10251
rect 25648 10220 25881 10248
rect 25648 10208 25654 10220
rect 25869 10217 25881 10220
rect 25915 10217 25927 10251
rect 25869 10211 25927 10217
rect 22612 10152 22876 10180
rect 22612 10140 22618 10152
rect 19208 10084 19840 10112
rect 19889 10115 19947 10121
rect 19208 10072 19214 10084
rect 19889 10081 19901 10115
rect 19935 10112 19947 10115
rect 20254 10112 20260 10124
rect 19935 10084 20260 10112
rect 19935 10081 19947 10084
rect 19889 10075 19947 10081
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 20441 10115 20499 10121
rect 20441 10081 20453 10115
rect 20487 10081 20499 10115
rect 20441 10075 20499 10081
rect 23017 10115 23075 10121
rect 23017 10081 23029 10115
rect 23063 10112 23075 10115
rect 23124 10112 23152 10208
rect 23063 10084 23152 10112
rect 23063 10081 23075 10084
rect 23017 10075 23075 10081
rect 11747 10016 12388 10044
rect 12529 10047 12587 10053
rect 11747 10013 11759 10016
rect 11701 10007 11759 10013
rect 12529 10013 12541 10047
rect 12575 10013 12587 10047
rect 12529 10007 12587 10013
rect 12805 10047 12863 10053
rect 12805 10013 12817 10047
rect 12851 10013 12863 10047
rect 12805 10007 12863 10013
rect 9401 9979 9459 9985
rect 9401 9945 9413 9979
rect 9447 9976 9459 9979
rect 12544 9976 12572 10007
rect 13262 10004 13268 10056
rect 13320 10004 13326 10056
rect 13906 10004 13912 10056
rect 13964 10044 13970 10056
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 13964 10016 14289 10044
rect 13964 10004 13970 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 15378 10004 15384 10056
rect 15436 10004 15442 10056
rect 15474 10047 15532 10053
rect 15474 10013 15486 10047
rect 15520 10013 15532 10047
rect 15474 10007 15532 10013
rect 13280 9976 13308 10004
rect 9447 9948 13308 9976
rect 9447 9945 9459 9948
rect 9401 9939 9459 9945
rect 13354 9936 13360 9988
rect 13412 9976 13418 9988
rect 15286 9976 15292 9988
rect 13412 9948 15292 9976
rect 13412 9936 13418 9948
rect 15286 9936 15292 9948
rect 15344 9936 15350 9988
rect 9030 9868 9036 9920
rect 9088 9868 9094 9920
rect 9858 9868 9864 9920
rect 9916 9908 9922 9920
rect 10410 9908 10416 9920
rect 9916 9880 10416 9908
rect 9916 9868 9922 9880
rect 10410 9868 10416 9880
rect 10468 9868 10474 9920
rect 10686 9868 10692 9920
rect 10744 9868 10750 9920
rect 11057 9911 11115 9917
rect 11057 9877 11069 9911
rect 11103 9908 11115 9911
rect 11146 9908 11152 9920
rect 11103 9880 11152 9908
rect 11103 9877 11115 9880
rect 11057 9871 11115 9877
rect 11146 9868 11152 9880
rect 11204 9868 11210 9920
rect 11974 9868 11980 9920
rect 12032 9908 12038 9920
rect 12805 9911 12863 9917
rect 12805 9908 12817 9911
rect 12032 9880 12817 9908
rect 12032 9868 12038 9880
rect 12805 9877 12817 9880
rect 12851 9877 12863 9911
rect 12805 9871 12863 9877
rect 13078 9868 13084 9920
rect 13136 9908 13142 9920
rect 13557 9911 13615 9917
rect 13557 9908 13569 9911
rect 13136 9880 13569 9908
rect 13136 9868 13142 9880
rect 13557 9877 13569 9880
rect 13603 9877 13615 9911
rect 13557 9871 13615 9877
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 14093 9911 14151 9917
rect 14093 9908 14105 9911
rect 13872 9880 14105 9908
rect 13872 9868 13878 9880
rect 14093 9877 14105 9880
rect 14139 9877 14151 9911
rect 14093 9871 14151 9877
rect 14366 9868 14372 9920
rect 14424 9908 14430 9920
rect 15488 9908 15516 10007
rect 15654 10004 15660 10056
rect 15712 10004 15718 10056
rect 15887 10047 15945 10053
rect 15887 10013 15899 10047
rect 15933 10044 15945 10047
rect 16298 10044 16304 10056
rect 15933 10016 16304 10044
rect 15933 10013 15945 10016
rect 15887 10007 15945 10013
rect 16298 10004 16304 10016
rect 16356 10004 16362 10056
rect 17954 10004 17960 10056
rect 18012 10004 18018 10056
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 18417 10047 18475 10053
rect 18417 10044 18429 10047
rect 18380 10016 18429 10044
rect 18380 10004 18386 10016
rect 18417 10013 18429 10016
rect 18463 10013 18475 10047
rect 18417 10007 18475 10013
rect 19981 10047 20039 10053
rect 19981 10013 19993 10047
rect 20027 10044 20039 10047
rect 20070 10044 20076 10056
rect 20027 10016 20076 10044
rect 20027 10013 20039 10016
rect 19981 10007 20039 10013
rect 20070 10004 20076 10016
rect 20128 10004 20134 10056
rect 20346 10004 20352 10056
rect 20404 10044 20410 10056
rect 20456 10044 20484 10075
rect 20404 10016 20484 10044
rect 20404 10004 20410 10016
rect 21634 10004 21640 10056
rect 21692 10044 21698 10056
rect 22281 10047 22339 10053
rect 22281 10044 22293 10047
rect 21692 10016 22293 10044
rect 21692 10004 21698 10016
rect 22281 10013 22293 10016
rect 22327 10013 22339 10047
rect 22281 10007 22339 10013
rect 22465 10047 22523 10053
rect 22465 10013 22477 10047
rect 22511 10013 22523 10047
rect 22465 10007 22523 10013
rect 15749 9979 15807 9985
rect 15749 9945 15761 9979
rect 15795 9976 15807 9979
rect 15795 9948 16804 9976
rect 15795 9945 15807 9948
rect 15749 9939 15807 9945
rect 14424 9880 15516 9908
rect 14424 9868 14430 9880
rect 15562 9868 15568 9920
rect 15620 9908 15626 9920
rect 16025 9911 16083 9917
rect 16025 9908 16037 9911
rect 15620 9880 16037 9908
rect 15620 9868 15626 9880
rect 16025 9877 16037 9880
rect 16071 9877 16083 9911
rect 16776 9908 16804 9948
rect 16850 9936 16856 9988
rect 16908 9936 16914 9988
rect 22480 9976 22508 10007
rect 22646 10004 22652 10056
rect 22704 10044 22710 10056
rect 23106 10044 23112 10056
rect 22704 10016 23112 10044
rect 22704 10004 22710 10016
rect 23106 10004 23112 10016
rect 23164 10004 23170 10056
rect 26145 10047 26203 10053
rect 26145 10013 26157 10047
rect 26191 10044 26203 10047
rect 26418 10044 26424 10056
rect 26191 10016 26424 10044
rect 26191 10013 26203 10016
rect 26145 10007 26203 10013
rect 26418 10004 26424 10016
rect 26476 10004 26482 10056
rect 22554 9976 22560 9988
rect 18248 9948 22560 9976
rect 18248 9908 18276 9948
rect 22554 9936 22560 9948
rect 22612 9936 22618 9988
rect 22830 9936 22836 9988
rect 22888 9936 22894 9988
rect 25869 9979 25927 9985
rect 25869 9945 25881 9979
rect 25915 9976 25927 9979
rect 26234 9976 26240 9988
rect 25915 9948 26240 9976
rect 25915 9945 25927 9948
rect 25869 9939 25927 9945
rect 26234 9936 26240 9948
rect 26292 9936 26298 9988
rect 16776 9880 18276 9908
rect 16025 9871 16083 9877
rect 18322 9868 18328 9920
rect 18380 9868 18386 9920
rect 19058 9868 19064 9920
rect 19116 9868 19122 9920
rect 22094 9868 22100 9920
rect 22152 9908 22158 9920
rect 22373 9911 22431 9917
rect 22373 9908 22385 9911
rect 22152 9880 22385 9908
rect 22152 9868 22158 9880
rect 22373 9877 22385 9880
rect 22419 9877 22431 9911
rect 22373 9871 22431 9877
rect 26053 9911 26111 9917
rect 26053 9877 26065 9911
rect 26099 9908 26111 9911
rect 26510 9908 26516 9920
rect 26099 9880 26516 9908
rect 26099 9877 26111 9880
rect 26053 9871 26111 9877
rect 26510 9868 26516 9880
rect 26568 9868 26574 9920
rect 1104 9818 29595 9840
rect 1104 9766 8032 9818
rect 8084 9766 8096 9818
rect 8148 9766 8160 9818
rect 8212 9766 8224 9818
rect 8276 9766 8288 9818
rect 8340 9766 15115 9818
rect 15167 9766 15179 9818
rect 15231 9766 15243 9818
rect 15295 9766 15307 9818
rect 15359 9766 15371 9818
rect 15423 9766 22198 9818
rect 22250 9766 22262 9818
rect 22314 9766 22326 9818
rect 22378 9766 22390 9818
rect 22442 9766 22454 9818
rect 22506 9766 29281 9818
rect 29333 9766 29345 9818
rect 29397 9766 29409 9818
rect 29461 9766 29473 9818
rect 29525 9766 29537 9818
rect 29589 9766 29595 9818
rect 1104 9744 29595 9766
rect 3697 9707 3755 9713
rect 3697 9673 3709 9707
rect 3743 9704 3755 9707
rect 3743 9676 4108 9704
rect 3743 9673 3755 9676
rect 3697 9667 3755 9673
rect 4080 9648 4108 9676
rect 6546 9664 6552 9716
rect 6604 9664 6610 9716
rect 9677 9707 9735 9713
rect 9677 9673 9689 9707
rect 9723 9704 9735 9707
rect 9950 9704 9956 9716
rect 9723 9676 9956 9704
rect 9723 9673 9735 9676
rect 9677 9667 9735 9673
rect 2222 9636 2228 9648
rect 1964 9608 2228 9636
rect 1964 9577 1992 9608
rect 2222 9596 2228 9608
rect 2280 9596 2286 9648
rect 4062 9596 4068 9648
rect 4120 9596 4126 9648
rect 5261 9639 5319 9645
rect 5261 9636 5273 9639
rect 5184 9608 5273 9636
rect 5184 9580 5212 9608
rect 5261 9605 5273 9608
rect 5307 9605 5319 9639
rect 5261 9599 5319 9605
rect 6270 9596 6276 9648
rect 6328 9636 6334 9648
rect 6457 9639 6515 9645
rect 6457 9636 6469 9639
rect 6328 9608 6469 9636
rect 6328 9596 6334 9608
rect 6457 9605 6469 9608
rect 6503 9605 6515 9639
rect 6564 9636 6592 9664
rect 7009 9639 7067 9645
rect 7009 9636 7021 9639
rect 6564 9608 7021 9636
rect 6457 9599 6515 9605
rect 7009 9605 7021 9608
rect 7055 9605 7067 9639
rect 9692 9636 9720 9667
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 10502 9704 10508 9716
rect 10152 9676 10508 9704
rect 10152 9645 10180 9676
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 10594 9664 10600 9716
rect 10652 9664 10658 9716
rect 10962 9704 10968 9716
rect 10888 9676 10968 9704
rect 7009 9599 7067 9605
rect 8772 9608 9720 9636
rect 10137 9639 10195 9645
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 3326 9528 3332 9580
rect 3384 9568 3390 9580
rect 3786 9568 3792 9580
rect 3384 9540 3792 9568
rect 3384 9528 3390 9540
rect 3786 9528 3792 9540
rect 3844 9528 3850 9580
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5077 9571 5135 9577
rect 5077 9568 5089 9571
rect 5031 9540 5089 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5077 9537 5089 9540
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 5166 9528 5172 9580
rect 5224 9528 5230 9580
rect 5345 9571 5403 9577
rect 5345 9568 5357 9571
rect 5276 9540 5357 9568
rect 2225 9503 2283 9509
rect 2225 9469 2237 9503
rect 2271 9500 2283 9503
rect 4154 9500 4160 9512
rect 2271 9472 4160 9500
rect 2271 9469 2283 9472
rect 2225 9463 2283 9469
rect 4154 9460 4160 9472
rect 4212 9460 4218 9512
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9469 4399 9503
rect 5276 9500 5304 9540
rect 5345 9537 5357 9540
rect 5391 9537 5403 9571
rect 5345 9531 5403 9537
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9568 5503 9571
rect 5534 9568 5540 9580
rect 5491 9540 5540 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 6914 9528 6920 9580
rect 6972 9528 6978 9580
rect 8772 9577 8800 9608
rect 10137 9605 10149 9639
rect 10183 9605 10195 9639
rect 10137 9599 10195 9605
rect 10226 9596 10232 9648
rect 10284 9596 10290 9648
rect 10367 9639 10425 9645
rect 10367 9605 10379 9639
rect 10413 9636 10425 9639
rect 10686 9636 10692 9648
rect 10413 9608 10692 9636
rect 10413 9605 10425 9608
rect 10367 9599 10425 9605
rect 10686 9596 10692 9608
rect 10744 9596 10750 9648
rect 10888 9645 10916 9676
rect 10962 9664 10968 9676
rect 11020 9664 11026 9716
rect 16850 9664 16856 9716
rect 16908 9704 16914 9716
rect 17221 9707 17279 9713
rect 17221 9704 17233 9707
rect 16908 9676 17233 9704
rect 16908 9664 16914 9676
rect 17221 9673 17233 9676
rect 17267 9673 17279 9707
rect 17221 9667 17279 9673
rect 17773 9707 17831 9713
rect 17773 9673 17785 9707
rect 17819 9704 17831 9707
rect 18506 9704 18512 9716
rect 17819 9676 18512 9704
rect 17819 9673 17831 9676
rect 17773 9667 17831 9673
rect 18506 9664 18512 9676
rect 18564 9664 18570 9716
rect 21726 9664 21732 9716
rect 21784 9704 21790 9716
rect 21784 9676 22094 9704
rect 21784 9664 21790 9676
rect 10873 9639 10931 9645
rect 10873 9605 10885 9639
rect 10919 9636 10931 9639
rect 11149 9639 11207 9645
rect 10919 9608 11100 9636
rect 10919 9605 10931 9608
rect 10873 9599 10931 9605
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 9030 9528 9036 9580
rect 9088 9568 9094 9580
rect 9309 9571 9367 9577
rect 9309 9568 9321 9571
rect 9088 9540 9321 9568
rect 9088 9528 9094 9540
rect 9309 9537 9321 9540
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 9539 9571 9597 9577
rect 9539 9537 9551 9571
rect 9585 9568 9597 9571
rect 9858 9568 9864 9580
rect 9585 9540 9864 9568
rect 9585 9537 9597 9540
rect 9539 9531 9597 9537
rect 9858 9528 9864 9540
rect 9916 9528 9922 9580
rect 10045 9571 10103 9577
rect 10045 9537 10057 9571
rect 10091 9568 10103 9571
rect 10505 9571 10563 9577
rect 10091 9540 10272 9568
rect 10091 9537 10103 9540
rect 10045 9531 10103 9537
rect 4341 9463 4399 9469
rect 4908 9472 5304 9500
rect 8665 9503 8723 9509
rect 4356 9376 4384 9463
rect 4338 9324 4344 9376
rect 4396 9324 4402 9376
rect 4908 9364 4936 9472
rect 8665 9469 8677 9503
rect 8711 9469 8723 9503
rect 8665 9463 8723 9469
rect 4982 9392 4988 9444
rect 5040 9432 5046 9444
rect 5902 9432 5908 9444
rect 5040 9404 5908 9432
rect 5040 9392 5046 9404
rect 5902 9392 5908 9404
rect 5960 9432 5966 9444
rect 6457 9435 6515 9441
rect 6457 9432 6469 9435
rect 5960 9404 6469 9432
rect 5960 9392 5966 9404
rect 6457 9401 6469 9404
rect 6503 9401 6515 9435
rect 6457 9395 6515 9401
rect 5074 9364 5080 9376
rect 4908 9336 5080 9364
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 5626 9324 5632 9376
rect 5684 9324 5690 9376
rect 6472 9364 6500 9395
rect 6546 9392 6552 9444
rect 6604 9432 6610 9444
rect 8481 9435 8539 9441
rect 8481 9432 8493 9435
rect 6604 9404 8493 9432
rect 6604 9392 6610 9404
rect 8481 9401 8493 9404
rect 8527 9401 8539 9435
rect 8481 9395 8539 9401
rect 6638 9364 6644 9376
rect 6472 9336 6644 9364
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 7190 9324 7196 9376
rect 7248 9324 7254 9376
rect 8680 9364 8708 9463
rect 8846 9460 8852 9512
rect 8904 9460 8910 9512
rect 8941 9503 8999 9509
rect 8941 9469 8953 9503
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 8956 9432 8984 9463
rect 9122 9460 9128 9512
rect 9180 9460 9186 9512
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9500 9459 9503
rect 9674 9500 9680 9512
rect 9447 9472 9680 9500
rect 9447 9469 9459 9472
rect 9401 9463 9459 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 9766 9460 9772 9512
rect 9824 9460 9830 9512
rect 10244 9444 10272 9540
rect 10505 9537 10517 9571
rect 10551 9537 10563 9571
rect 10505 9531 10563 9537
rect 10597 9571 10655 9577
rect 10597 9537 10609 9571
rect 10643 9537 10655 9571
rect 10965 9571 11023 9577
rect 10965 9568 10977 9571
rect 10597 9531 10655 9537
rect 10704 9540 10977 9568
rect 10410 9460 10416 9512
rect 10468 9460 10474 9512
rect 9861 9435 9919 9441
rect 9861 9432 9873 9435
rect 8956 9404 9873 9432
rect 9861 9401 9873 9404
rect 9907 9401 9919 9435
rect 9861 9395 9919 9401
rect 10226 9392 10232 9444
rect 10284 9392 10290 9444
rect 10428 9364 10456 9460
rect 10520 9376 10548 9531
rect 10612 9432 10640 9531
rect 10704 9512 10732 9540
rect 10965 9537 10977 9540
rect 11011 9537 11023 9571
rect 11072 9568 11100 9608
rect 11149 9605 11161 9639
rect 11195 9636 11207 9639
rect 11330 9636 11336 9648
rect 11195 9608 11336 9636
rect 11195 9605 11207 9608
rect 11149 9599 11207 9605
rect 11330 9596 11336 9608
rect 11388 9636 11394 9648
rect 11388 9608 11928 9636
rect 11388 9596 11394 9608
rect 11900 9577 11928 9608
rect 13170 9596 13176 9648
rect 13228 9596 13234 9648
rect 13446 9636 13452 9648
rect 13280 9608 13452 9636
rect 11241 9571 11299 9577
rect 11241 9568 11253 9571
rect 11072 9540 11253 9568
rect 10965 9531 11023 9537
rect 11241 9537 11253 9540
rect 11287 9537 11299 9571
rect 11241 9531 11299 9537
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 12342 9528 12348 9580
rect 12400 9568 12406 9580
rect 13280 9577 13308 9608
rect 13446 9596 13452 9608
rect 13504 9596 13510 9648
rect 13541 9639 13599 9645
rect 13541 9605 13553 9639
rect 13587 9636 13599 9639
rect 13814 9636 13820 9648
rect 13587 9608 13820 9636
rect 13587 9605 13599 9608
rect 13541 9599 13599 9605
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 14274 9596 14280 9648
rect 14332 9596 14338 9648
rect 16684 9608 19104 9636
rect 16684 9577 16712 9608
rect 19076 9580 19104 9608
rect 12529 9571 12587 9577
rect 12529 9568 12541 9571
rect 12400 9540 12541 9568
rect 12400 9528 12434 9540
rect 12529 9537 12541 9540
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 13265 9571 13323 9577
rect 13265 9537 13277 9571
rect 13311 9537 13323 9571
rect 13265 9531 13323 9537
rect 16669 9571 16727 9577
rect 16669 9537 16681 9571
rect 16715 9537 16727 9571
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16669 9531 16727 9537
rect 16776 9540 16865 9568
rect 10686 9460 10692 9512
rect 10744 9460 10750 9512
rect 11054 9460 11060 9512
rect 11112 9460 11118 9512
rect 10965 9435 11023 9441
rect 10612 9404 10732 9432
rect 8680 9336 10456 9364
rect 10502 9324 10508 9376
rect 10560 9324 10566 9376
rect 10704 9364 10732 9404
rect 10965 9401 10977 9435
rect 11011 9432 11023 9435
rect 11072 9432 11100 9460
rect 11011 9404 11100 9432
rect 11011 9401 11023 9404
rect 10965 9395 11023 9401
rect 11422 9364 11428 9376
rect 10704 9336 11428 9364
rect 11422 9324 11428 9336
rect 11480 9364 11486 9376
rect 12406 9364 12434 9528
rect 16776 9512 16804 9540
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 16945 9571 17003 9577
rect 16945 9537 16957 9571
rect 16991 9537 17003 9571
rect 16945 9531 17003 9537
rect 14090 9460 14096 9512
rect 14148 9500 14154 9512
rect 15289 9503 15347 9509
rect 15289 9500 15301 9503
rect 14148 9472 15301 9500
rect 14148 9460 14154 9472
rect 15289 9469 15301 9472
rect 15335 9469 15347 9503
rect 15289 9463 15347 9469
rect 15304 9432 15332 9463
rect 16758 9460 16764 9512
rect 16816 9460 16822 9512
rect 16960 9432 16988 9531
rect 17034 9528 17040 9580
rect 17092 9528 17098 9580
rect 17770 9571 17828 9577
rect 17770 9537 17782 9571
rect 17816 9568 17828 9571
rect 17862 9568 17868 9580
rect 17816 9540 17868 9568
rect 17816 9537 17828 9540
rect 17770 9531 17828 9537
rect 17862 9528 17868 9540
rect 17920 9528 17926 9580
rect 18046 9528 18052 9580
rect 18104 9528 18110 9580
rect 18141 9571 18199 9577
rect 18141 9537 18153 9571
rect 18187 9568 18199 9571
rect 18322 9568 18328 9580
rect 18187 9540 18328 9568
rect 18187 9537 18199 9540
rect 18141 9531 18199 9537
rect 18322 9528 18328 9540
rect 18380 9528 18386 9580
rect 18414 9528 18420 9580
rect 18472 9577 18478 9580
rect 18472 9571 18508 9577
rect 18496 9537 18508 9571
rect 18472 9531 18508 9537
rect 18472 9528 18478 9531
rect 19058 9528 19064 9580
rect 19116 9528 19122 9580
rect 22066 9568 22094 9676
rect 25590 9596 25596 9648
rect 25648 9636 25654 9648
rect 27709 9639 27767 9645
rect 27709 9636 27721 9639
rect 25648 9608 27721 9636
rect 25648 9596 25654 9608
rect 27709 9605 27721 9608
rect 27755 9605 27767 9639
rect 27709 9599 27767 9605
rect 22646 9568 22652 9580
rect 22066 9540 22652 9568
rect 22646 9528 22652 9540
rect 22704 9528 22710 9580
rect 23382 9528 23388 9580
rect 23440 9528 23446 9580
rect 25498 9528 25504 9580
rect 25556 9568 25562 9580
rect 26237 9571 26295 9577
rect 26237 9568 26249 9571
rect 25556 9540 26249 9568
rect 25556 9528 25562 9540
rect 26237 9537 26249 9540
rect 26283 9537 26295 9571
rect 26237 9531 26295 9537
rect 26467 9571 26525 9577
rect 26467 9537 26479 9571
rect 26513 9568 26525 9571
rect 27893 9571 27951 9577
rect 26513 9540 26648 9568
rect 26513 9537 26525 9540
rect 26467 9531 26525 9537
rect 17052 9500 17080 9528
rect 18064 9500 18092 9528
rect 17052 9472 18092 9500
rect 18233 9503 18291 9509
rect 18233 9469 18245 9503
rect 18279 9469 18291 9503
rect 18233 9463 18291 9469
rect 18969 9503 19027 9509
rect 18969 9469 18981 9503
rect 19015 9469 19027 9503
rect 23400 9500 23428 9528
rect 26620 9500 26648 9540
rect 27893 9537 27905 9571
rect 27939 9537 27951 9571
rect 27893 9531 27951 9537
rect 27985 9571 28043 9577
rect 27985 9537 27997 9571
rect 28031 9537 28043 9571
rect 27985 9531 28043 9537
rect 26878 9500 26884 9512
rect 23400 9472 26884 9500
rect 18969 9463 19027 9469
rect 15304 9404 16988 9432
rect 17126 9392 17132 9444
rect 17184 9432 17190 9444
rect 18248 9432 18276 9463
rect 18984 9432 19012 9463
rect 26878 9460 26884 9472
rect 26936 9500 26942 9512
rect 26973 9503 27031 9509
rect 26973 9500 26985 9503
rect 26936 9472 26985 9500
rect 26936 9460 26942 9472
rect 26973 9469 26985 9472
rect 27019 9469 27031 9503
rect 26973 9463 27031 9469
rect 27908 9444 27936 9531
rect 17184 9404 19012 9432
rect 17184 9392 17190 9404
rect 26142 9392 26148 9444
rect 26200 9432 26206 9444
rect 27617 9435 27675 9441
rect 27617 9432 27629 9435
rect 26200 9404 27629 9432
rect 26200 9392 26206 9404
rect 27617 9401 27629 9404
rect 27663 9401 27675 9435
rect 27617 9395 27675 9401
rect 27890 9392 27896 9444
rect 27948 9392 27954 9444
rect 11480 9336 12434 9364
rect 11480 9324 11486 9336
rect 13722 9324 13728 9376
rect 13780 9364 13786 9376
rect 14274 9364 14280 9376
rect 13780 9336 14280 9364
rect 13780 9324 13786 9336
rect 14274 9324 14280 9336
rect 14332 9324 14338 9376
rect 17586 9324 17592 9376
rect 17644 9324 17650 9376
rect 17954 9324 17960 9376
rect 18012 9364 18018 9376
rect 18325 9367 18383 9373
rect 18325 9364 18337 9367
rect 18012 9336 18337 9364
rect 18012 9324 18018 9336
rect 18325 9333 18337 9336
rect 18371 9333 18383 9367
rect 18325 9327 18383 9333
rect 18877 9367 18935 9373
rect 18877 9333 18889 9367
rect 18923 9364 18935 9367
rect 19334 9364 19340 9376
rect 18923 9336 19340 9364
rect 18923 9333 18935 9336
rect 18877 9327 18935 9333
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 26329 9367 26387 9373
rect 26329 9333 26341 9367
rect 26375 9364 26387 9367
rect 26602 9364 26608 9376
rect 26375 9336 26608 9364
rect 26375 9333 26387 9336
rect 26329 9327 26387 9333
rect 26602 9324 26608 9336
rect 26660 9364 26666 9376
rect 28000 9364 28028 9531
rect 28166 9528 28172 9580
rect 28224 9528 28230 9580
rect 28261 9571 28319 9577
rect 28261 9537 28273 9571
rect 28307 9537 28319 9571
rect 28261 9531 28319 9537
rect 28074 9460 28080 9512
rect 28132 9500 28138 9512
rect 28276 9500 28304 9531
rect 28132 9472 28304 9500
rect 28132 9460 28138 9472
rect 26660 9336 28028 9364
rect 26660 9324 26666 9336
rect 1104 9274 29440 9296
rect 1104 9222 4491 9274
rect 4543 9222 4555 9274
rect 4607 9222 4619 9274
rect 4671 9222 4683 9274
rect 4735 9222 4747 9274
rect 4799 9222 11574 9274
rect 11626 9222 11638 9274
rect 11690 9222 11702 9274
rect 11754 9222 11766 9274
rect 11818 9222 11830 9274
rect 11882 9222 18657 9274
rect 18709 9222 18721 9274
rect 18773 9222 18785 9274
rect 18837 9222 18849 9274
rect 18901 9222 18913 9274
rect 18965 9222 25740 9274
rect 25792 9222 25804 9274
rect 25856 9222 25868 9274
rect 25920 9222 25932 9274
rect 25984 9222 25996 9274
rect 26048 9222 29440 9274
rect 1104 9200 29440 9222
rect 2120 9163 2178 9169
rect 2120 9129 2132 9163
rect 2166 9160 2178 9163
rect 5626 9160 5632 9172
rect 2166 9132 5632 9160
rect 2166 9129 2178 9132
rect 2120 9123 2178 9129
rect 5626 9120 5632 9132
rect 5684 9120 5690 9172
rect 5736 9132 13032 9160
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 4893 9095 4951 9101
rect 4893 9092 4905 9095
rect 4212 9064 4905 9092
rect 4212 9052 4218 9064
rect 4893 9061 4905 9064
rect 4939 9061 4951 9095
rect 4893 9055 4951 9061
rect 4982 9052 4988 9104
rect 5040 9092 5046 9104
rect 5353 9095 5411 9101
rect 5353 9092 5365 9095
rect 5040 9064 5365 9092
rect 5040 9052 5046 9064
rect 5353 9061 5365 9064
rect 5399 9061 5411 9095
rect 5353 9055 5411 9061
rect 5442 9052 5448 9104
rect 5500 9092 5506 9104
rect 5736 9092 5764 9132
rect 5500 9064 5764 9092
rect 5500 9052 5506 9064
rect 10226 9052 10232 9104
rect 10284 9092 10290 9104
rect 13004 9092 13032 9132
rect 13078 9120 13084 9172
rect 13136 9120 13142 9172
rect 17494 9120 17500 9172
rect 17552 9160 17558 9172
rect 22557 9163 22615 9169
rect 22557 9160 22569 9163
rect 17552 9132 22569 9160
rect 17552 9120 17558 9132
rect 22557 9129 22569 9132
rect 22603 9129 22615 9163
rect 22557 9123 22615 9129
rect 17310 9092 17316 9104
rect 10284 9064 11401 9092
rect 13004 9064 17316 9092
rect 10284 9052 10290 9064
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 9024 1915 9027
rect 2222 9024 2228 9036
rect 1903 8996 2228 9024
rect 1903 8993 1915 8996
rect 1857 8987 1915 8993
rect 2222 8984 2228 8996
rect 2280 8984 2286 9036
rect 3605 9027 3663 9033
rect 3605 8993 3617 9027
rect 3651 9024 3663 9027
rect 4338 9024 4344 9036
rect 3651 8996 4344 9024
rect 3651 8993 3663 8996
rect 3605 8987 3663 8993
rect 4338 8984 4344 8996
rect 4396 9024 4402 9036
rect 5813 9027 5871 9033
rect 5813 9024 5825 9027
rect 4396 8996 5825 9024
rect 4396 8984 4402 8996
rect 5813 8993 5825 8996
rect 5859 8993 5871 9027
rect 5813 8987 5871 8993
rect 6181 9027 6239 9033
rect 6181 8993 6193 9027
rect 6227 9024 6239 9027
rect 6227 8996 8984 9024
rect 6227 8993 6239 8996
rect 6181 8987 6239 8993
rect 8956 8968 8984 8996
rect 9122 8984 9128 9036
rect 9180 9024 9186 9036
rect 9309 9027 9367 9033
rect 9309 9024 9321 9027
rect 9180 8996 9321 9024
rect 9180 8984 9186 8996
rect 9309 8993 9321 8996
rect 9355 8993 9367 9027
rect 9309 8987 9367 8993
rect 9858 8984 9864 9036
rect 9916 9024 9922 9036
rect 10134 9024 10140 9036
rect 9916 8996 10140 9024
rect 9916 8984 9922 8996
rect 10134 8984 10140 8996
rect 10192 9024 10198 9036
rect 10192 8996 10732 9024
rect 10192 8984 10198 8996
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 5905 8959 5963 8965
rect 4295 8928 4384 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 3786 8888 3792 8900
rect 3358 8860 3792 8888
rect 3786 8848 3792 8860
rect 3844 8848 3850 8900
rect 4356 8832 4384 8928
rect 5905 8925 5917 8959
rect 5951 8956 5963 8959
rect 5994 8956 6000 8968
rect 5951 8928 6000 8956
rect 5951 8925 5963 8928
rect 5905 8919 5963 8925
rect 5994 8916 6000 8928
rect 6052 8956 6058 8968
rect 6454 8956 6460 8968
rect 6052 8928 6460 8956
rect 6052 8916 6058 8928
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 6546 8916 6552 8968
rect 6604 8916 6610 8968
rect 8938 8916 8944 8968
rect 8996 8916 9002 8968
rect 10704 8956 10732 8996
rect 10778 8984 10784 9036
rect 10836 9024 10842 9036
rect 11146 9024 11152 9036
rect 10836 8996 11152 9024
rect 10836 8984 10842 8996
rect 11146 8984 11152 8996
rect 11204 8984 11210 9036
rect 11373 9033 11401 9064
rect 17310 9052 17316 9064
rect 17368 9052 17374 9104
rect 22572 9092 22600 9123
rect 22830 9120 22836 9172
rect 22888 9160 22894 9172
rect 23017 9163 23075 9169
rect 23017 9160 23029 9163
rect 22888 9132 23029 9160
rect 22888 9120 22894 9132
rect 23017 9129 23029 9132
rect 23063 9129 23075 9163
rect 23017 9123 23075 9129
rect 26878 9120 26884 9172
rect 26936 9160 26942 9172
rect 27985 9163 28043 9169
rect 27985 9160 27997 9163
rect 26936 9132 27997 9160
rect 26936 9120 26942 9132
rect 27985 9129 27997 9132
rect 28031 9160 28043 9163
rect 28031 9132 28488 9160
rect 28031 9129 28043 9132
rect 27985 9123 28043 9129
rect 24026 9092 24032 9104
rect 22572 9064 24032 9092
rect 24026 9052 24032 9064
rect 24084 9052 24090 9104
rect 11358 9027 11416 9033
rect 11358 8993 11370 9027
rect 11404 9024 11416 9027
rect 11974 9024 11980 9036
rect 11404 8996 11980 9024
rect 11404 8993 11416 8996
rect 11358 8987 11416 8993
rect 11974 8984 11980 8996
rect 12032 8984 12038 9036
rect 14645 9027 14703 9033
rect 14645 8993 14657 9027
rect 14691 9024 14703 9027
rect 15746 9024 15752 9036
rect 14691 8996 15752 9024
rect 14691 8993 14703 8996
rect 14645 8987 14703 8993
rect 15746 8984 15752 8996
rect 15804 8984 15810 9036
rect 16666 8984 16672 9036
rect 16724 9024 16730 9036
rect 16724 8996 18184 9024
rect 16724 8984 16730 8996
rect 10873 8959 10931 8965
rect 10873 8956 10885 8959
rect 10704 8928 10885 8956
rect 10873 8925 10885 8928
rect 10919 8925 10931 8959
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 10873 8919 10931 8925
rect 11532 8928 11621 8956
rect 5353 8891 5411 8897
rect 5353 8857 5365 8891
rect 5399 8888 5411 8891
rect 6270 8888 6276 8900
rect 5399 8860 6276 8888
rect 5399 8857 5411 8860
rect 5353 8851 5411 8857
rect 6270 8848 6276 8860
rect 6328 8848 6334 8900
rect 7098 8848 7104 8900
rect 7156 8848 7162 8900
rect 10042 8848 10048 8900
rect 10100 8848 10106 8900
rect 11241 8891 11299 8897
rect 11241 8857 11253 8891
rect 11287 8888 11299 8891
rect 11330 8888 11336 8900
rect 11287 8860 11336 8888
rect 11287 8857 11299 8860
rect 11241 8851 11299 8857
rect 11330 8848 11336 8860
rect 11388 8848 11394 8900
rect 4338 8780 4344 8832
rect 4396 8780 4402 8832
rect 6086 8780 6092 8832
rect 6144 8780 6150 8832
rect 6288 8820 6316 8848
rect 7975 8823 8033 8829
rect 7975 8820 7987 8823
rect 6288 8792 7987 8820
rect 7975 8789 7987 8792
rect 8021 8789 8033 8823
rect 7975 8783 8033 8789
rect 9950 8780 9956 8832
rect 10008 8820 10014 8832
rect 11532 8829 11560 8928
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8956 11943 8959
rect 12250 8956 12256 8968
rect 11931 8928 12256 8956
rect 11931 8925 11943 8928
rect 11885 8919 11943 8925
rect 12250 8916 12256 8928
rect 12308 8916 12314 8968
rect 12989 8959 13047 8965
rect 12989 8925 13001 8959
rect 13035 8956 13047 8959
rect 13722 8956 13728 8968
rect 13035 8928 13728 8956
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 18156 8965 18184 8996
rect 22370 8984 22376 9036
rect 22428 8984 22434 9036
rect 22554 8984 22560 9036
rect 22612 8984 22618 9036
rect 22646 8984 22652 9036
rect 22704 8984 22710 9036
rect 26237 9027 26295 9033
rect 26237 9024 26249 9027
rect 24964 8996 26249 9024
rect 13817 8959 13875 8965
rect 13817 8925 13829 8959
rect 13863 8925 13875 8959
rect 13817 8919 13875 8925
rect 17957 8959 18015 8965
rect 17957 8925 17969 8959
rect 18003 8925 18015 8959
rect 17957 8919 18015 8925
rect 18141 8959 18199 8965
rect 18141 8925 18153 8959
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 13541 8891 13599 8897
rect 13541 8888 13553 8891
rect 13320 8860 13553 8888
rect 13320 8848 13326 8860
rect 13541 8857 13553 8860
rect 13587 8857 13599 8891
rect 13832 8888 13860 8919
rect 13906 8888 13912 8900
rect 13832 8860 13912 8888
rect 13541 8851 13599 8857
rect 13906 8848 13912 8860
rect 13964 8848 13970 8900
rect 10735 8823 10793 8829
rect 10735 8820 10747 8823
rect 10008 8792 10747 8820
rect 10008 8780 10014 8792
rect 10735 8789 10747 8792
rect 10781 8789 10793 8823
rect 10735 8783 10793 8789
rect 11517 8823 11575 8829
rect 11517 8789 11529 8823
rect 11563 8789 11575 8823
rect 13630 8820 13636 8832
rect 13688 8829 13694 8832
rect 13597 8792 13636 8820
rect 11517 8783 11575 8789
rect 13630 8780 13636 8792
rect 13688 8783 13697 8829
rect 13725 8823 13783 8829
rect 13725 8789 13737 8823
rect 13771 8820 13783 8823
rect 15197 8823 15255 8829
rect 15197 8820 15209 8823
rect 13771 8792 15209 8820
rect 13771 8789 13783 8792
rect 13725 8783 13783 8789
rect 15197 8789 15209 8792
rect 15243 8789 15255 8823
rect 17972 8820 18000 8919
rect 18322 8916 18328 8968
rect 18380 8916 18386 8968
rect 19334 8916 19340 8968
rect 19392 8956 19398 8968
rect 19392 8928 20668 8956
rect 19392 8916 19398 8928
rect 18230 8897 18236 8900
rect 18229 8888 18236 8897
rect 18191 8860 18236 8888
rect 18229 8851 18236 8860
rect 18230 8848 18236 8851
rect 18288 8848 18294 8900
rect 19889 8891 19947 8897
rect 19889 8888 19901 8891
rect 18340 8860 19901 8888
rect 18340 8820 18368 8860
rect 19889 8857 19901 8860
rect 19935 8857 19947 8891
rect 19889 8851 19947 8857
rect 20640 8832 20668 8928
rect 22094 8916 22100 8968
rect 22152 8916 22158 8968
rect 22189 8959 22247 8965
rect 22189 8925 22201 8959
rect 22235 8956 22247 8959
rect 22572 8956 22600 8984
rect 24964 8968 24992 8996
rect 26237 8993 26249 8996
rect 26283 8993 26295 9027
rect 26237 8987 26295 8993
rect 27246 8984 27252 9036
rect 27304 9024 27310 9036
rect 27304 8996 27752 9024
rect 27304 8984 27310 8996
rect 22235 8928 22600 8956
rect 22235 8925 22247 8928
rect 22189 8919 22247 8925
rect 22830 8916 22836 8968
rect 22888 8916 22894 8968
rect 24946 8916 24952 8968
rect 25004 8916 25010 8968
rect 25590 8916 25596 8968
rect 25648 8956 25654 8968
rect 25685 8959 25743 8965
rect 25685 8956 25697 8959
rect 25648 8928 25697 8956
rect 25648 8916 25654 8928
rect 25685 8925 25697 8928
rect 25731 8925 25743 8959
rect 25685 8919 25743 8925
rect 26142 8916 26148 8968
rect 26200 8916 26206 8968
rect 27724 8956 27752 8996
rect 27890 8956 27896 8968
rect 27724 8928 27896 8956
rect 27890 8916 27896 8928
rect 27948 8956 27954 8968
rect 28353 8959 28411 8965
rect 27948 8928 28304 8956
rect 27948 8916 27954 8928
rect 22557 8891 22615 8897
rect 22557 8888 22569 8891
rect 22112 8860 22569 8888
rect 22112 8832 22140 8860
rect 22557 8857 22569 8860
rect 22603 8888 22615 8891
rect 23382 8888 23388 8900
rect 22603 8860 23388 8888
rect 22603 8857 22615 8860
rect 22557 8851 22615 8857
rect 23382 8848 23388 8860
rect 23440 8848 23446 8900
rect 25774 8848 25780 8900
rect 25832 8848 25838 8900
rect 25866 8848 25872 8900
rect 25924 8848 25930 8900
rect 26007 8891 26065 8897
rect 26007 8857 26019 8891
rect 26053 8888 26065 8891
rect 26234 8888 26240 8900
rect 26053 8860 26240 8888
rect 26053 8857 26065 8860
rect 26007 8851 26065 8857
rect 26234 8848 26240 8860
rect 26292 8888 26298 8900
rect 26418 8888 26424 8900
rect 26292 8860 26424 8888
rect 26292 8848 26298 8860
rect 26418 8848 26424 8860
rect 26476 8848 26482 8900
rect 26513 8891 26571 8897
rect 26513 8857 26525 8891
rect 26559 8857 26571 8891
rect 26513 8851 26571 8857
rect 17972 8792 18368 8820
rect 15197 8783 15255 8789
rect 13688 8780 13694 8783
rect 18506 8780 18512 8832
rect 18564 8780 18570 8832
rect 20622 8780 20628 8832
rect 20680 8780 20686 8832
rect 21726 8780 21732 8832
rect 21784 8780 21790 8832
rect 22094 8780 22100 8832
rect 22152 8780 22158 8832
rect 22370 8780 22376 8832
rect 22428 8820 22434 8832
rect 24302 8820 24308 8832
rect 22428 8792 24308 8820
rect 22428 8780 22434 8792
rect 24302 8780 24308 8792
rect 24360 8780 24366 8832
rect 25501 8823 25559 8829
rect 25501 8789 25513 8823
rect 25547 8820 25559 8823
rect 26528 8820 26556 8851
rect 27062 8848 27068 8900
rect 27120 8848 27126 8900
rect 27798 8848 27804 8900
rect 27856 8888 27862 8900
rect 28169 8891 28227 8897
rect 28169 8888 28181 8891
rect 27856 8860 28181 8888
rect 27856 8848 27862 8860
rect 28169 8857 28181 8860
rect 28215 8857 28227 8891
rect 28276 8888 28304 8928
rect 28353 8925 28365 8959
rect 28399 8956 28411 8959
rect 28460 8956 28488 9132
rect 28399 8928 28488 8956
rect 28399 8925 28411 8928
rect 28353 8919 28411 8925
rect 28537 8891 28595 8897
rect 28537 8888 28549 8891
rect 28276 8860 28549 8888
rect 28169 8851 28227 8857
rect 28537 8857 28549 8860
rect 28583 8857 28595 8891
rect 28537 8851 28595 8857
rect 25547 8792 26556 8820
rect 25547 8789 25559 8792
rect 25501 8783 25559 8789
rect 1104 8730 29595 8752
rect 1104 8678 8032 8730
rect 8084 8678 8096 8730
rect 8148 8678 8160 8730
rect 8212 8678 8224 8730
rect 8276 8678 8288 8730
rect 8340 8678 15115 8730
rect 15167 8678 15179 8730
rect 15231 8678 15243 8730
rect 15295 8678 15307 8730
rect 15359 8678 15371 8730
rect 15423 8678 22198 8730
rect 22250 8678 22262 8730
rect 22314 8678 22326 8730
rect 22378 8678 22390 8730
rect 22442 8678 22454 8730
rect 22506 8678 29281 8730
rect 29333 8678 29345 8730
rect 29397 8678 29409 8730
rect 29461 8678 29473 8730
rect 29525 8678 29537 8730
rect 29589 8678 29595 8730
rect 1104 8656 29595 8678
rect 2222 8576 2228 8628
rect 2280 8576 2286 8628
rect 4154 8576 4160 8628
rect 4212 8576 4218 8628
rect 5442 8576 5448 8628
rect 5500 8576 5506 8628
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8585 5687 8619
rect 5629 8579 5687 8585
rect 2240 8548 2268 8576
rect 2682 8548 2688 8560
rect 2148 8520 2688 8548
rect 1670 8440 1676 8492
rect 1728 8480 1734 8492
rect 2148 8489 2176 8520
rect 2682 8508 2688 8520
rect 2740 8508 2746 8560
rect 4172 8548 4200 8576
rect 3988 8520 4200 8548
rect 4249 8551 4307 8557
rect 2133 8483 2191 8489
rect 2133 8480 2145 8483
rect 1728 8452 2145 8480
rect 1728 8440 1734 8452
rect 2133 8449 2145 8452
rect 2179 8449 2191 8483
rect 3786 8480 3792 8492
rect 3542 8452 3792 8480
rect 2133 8443 2191 8449
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 3988 8489 4016 8520
rect 4249 8517 4261 8551
rect 4295 8548 4307 8551
rect 4985 8551 5043 8557
rect 4295 8520 4936 8548
rect 4295 8517 4307 8520
rect 4249 8511 4307 8517
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 4154 8440 4160 8492
rect 4212 8440 4218 8492
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4798 8480 4804 8492
rect 4387 8452 4804 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 4908 8480 4936 8520
rect 4985 8517 4997 8551
rect 5031 8548 5043 8551
rect 5644 8548 5672 8579
rect 6086 8576 6092 8628
rect 6144 8576 6150 8628
rect 6454 8576 6460 8628
rect 6512 8616 6518 8628
rect 6730 8616 6736 8628
rect 6512 8588 6736 8616
rect 6512 8576 6518 8588
rect 6730 8576 6736 8588
rect 6788 8576 6794 8628
rect 9950 8616 9956 8628
rect 7668 8588 9168 8616
rect 5031 8520 5672 8548
rect 5031 8517 5043 8520
rect 4985 8511 5043 8517
rect 5810 8508 5816 8560
rect 5868 8548 5874 8560
rect 5994 8548 6000 8560
rect 5868 8520 6000 8548
rect 5868 8508 5874 8520
rect 5994 8508 6000 8520
rect 6052 8508 6058 8560
rect 5261 8483 5319 8489
rect 4908 8452 5120 8480
rect 5092 8424 5120 8452
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5442 8480 5448 8492
rect 5307 8452 5448 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 6104 8480 6132 8576
rect 7668 8557 7696 8588
rect 7653 8551 7711 8557
rect 7653 8548 7665 8551
rect 5552 8452 6132 8480
rect 6196 8520 7665 8548
rect 2409 8415 2467 8421
rect 2409 8381 2421 8415
rect 2455 8412 2467 8415
rect 2455 8384 4568 8412
rect 2455 8381 2467 8384
rect 2409 8375 2467 8381
rect 3881 8347 3939 8353
rect 3881 8313 3893 8347
rect 3927 8344 3939 8347
rect 4338 8344 4344 8356
rect 3927 8316 4344 8344
rect 3927 8313 3939 8316
rect 3881 8307 3939 8313
rect 4338 8304 4344 8316
rect 4396 8344 4402 8356
rect 4540 8353 4568 8384
rect 5074 8372 5080 8424
rect 5132 8372 5138 8424
rect 5169 8415 5227 8421
rect 5169 8381 5181 8415
rect 5215 8412 5227 8415
rect 5552 8412 5580 8452
rect 5215 8384 5580 8412
rect 5813 8415 5871 8421
rect 5215 8381 5227 8384
rect 5169 8375 5227 8381
rect 5813 8381 5825 8415
rect 5859 8381 5871 8415
rect 5813 8375 5871 8381
rect 4525 8347 4583 8353
rect 4396 8316 4476 8344
rect 4396 8304 4402 8316
rect 4448 8276 4476 8316
rect 4525 8313 4537 8347
rect 4571 8313 4583 8347
rect 5828 8344 5856 8375
rect 5902 8372 5908 8424
rect 5960 8372 5966 8424
rect 5994 8372 6000 8424
rect 6052 8372 6058 8424
rect 6089 8415 6147 8421
rect 6089 8381 6101 8415
rect 6135 8412 6147 8415
rect 6196 8412 6224 8520
rect 7653 8517 7665 8520
rect 7699 8517 7711 8551
rect 7653 8511 7711 8517
rect 8297 8551 8355 8557
rect 8297 8517 8309 8551
rect 8343 8517 8355 8551
rect 8297 8511 8355 8517
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 6822 8480 6828 8492
rect 6328 8452 6828 8480
rect 6328 8440 6334 8452
rect 6822 8440 6828 8452
rect 6880 8480 6886 8492
rect 7285 8483 7343 8489
rect 7285 8480 7297 8483
rect 6880 8452 7297 8480
rect 6880 8440 6886 8452
rect 7285 8449 7297 8452
rect 7331 8480 7343 8483
rect 8312 8480 8340 8511
rect 9030 8508 9036 8560
rect 9088 8508 9094 8560
rect 7331 8452 8340 8480
rect 9140 8480 9168 8588
rect 9232 8588 9956 8616
rect 9232 8557 9260 8588
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 13262 8576 13268 8628
rect 13320 8616 13326 8628
rect 13357 8619 13415 8625
rect 13357 8616 13369 8619
rect 13320 8588 13369 8616
rect 13320 8576 13326 8588
rect 13357 8585 13369 8588
rect 13403 8585 13415 8619
rect 13357 8579 13415 8585
rect 13556 8588 15516 8616
rect 9217 8551 9275 8557
rect 9217 8517 9229 8551
rect 9263 8517 9275 8551
rect 13556 8548 13584 8588
rect 9217 8511 9275 8517
rect 13096 8520 13584 8548
rect 9674 8480 9680 8492
rect 9140 8452 9680 8480
rect 7331 8449 7343 8452
rect 7285 8443 7343 8449
rect 9674 8440 9680 8452
rect 9732 8480 9738 8492
rect 10502 8480 10508 8492
rect 9732 8452 10508 8480
rect 9732 8440 9738 8452
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 13096 8489 13124 8520
rect 13630 8508 13636 8560
rect 13688 8548 13694 8560
rect 13725 8551 13783 8557
rect 13725 8548 13737 8551
rect 13688 8520 13737 8548
rect 13688 8508 13694 8520
rect 13725 8517 13737 8520
rect 13771 8517 13783 8551
rect 13725 8511 13783 8517
rect 14274 8508 14280 8560
rect 14332 8508 14338 8560
rect 15488 8557 15516 8588
rect 16574 8576 16580 8628
rect 16632 8576 16638 8628
rect 17586 8576 17592 8628
rect 17644 8576 17650 8628
rect 18506 8576 18512 8628
rect 18564 8576 18570 8628
rect 20622 8576 20628 8628
rect 20680 8576 20686 8628
rect 21726 8576 21732 8628
rect 21784 8576 21790 8628
rect 22830 8576 22836 8628
rect 22888 8616 22894 8628
rect 26234 8616 26240 8628
rect 22888 8588 26240 8616
rect 22888 8576 22894 8588
rect 26234 8576 26240 8588
rect 26292 8576 26298 8628
rect 26789 8619 26847 8625
rect 26789 8585 26801 8619
rect 26835 8616 26847 8619
rect 28166 8616 28172 8628
rect 26835 8588 28172 8616
rect 26835 8585 26847 8588
rect 26789 8579 26847 8585
rect 15473 8551 15531 8557
rect 15473 8517 15485 8551
rect 15519 8548 15531 8551
rect 15746 8548 15752 8560
rect 15519 8520 15752 8548
rect 15519 8517 15531 8520
rect 15473 8511 15531 8517
rect 15746 8508 15752 8520
rect 15804 8508 15810 8560
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8449 13139 8483
rect 16592 8480 16620 8576
rect 17604 8548 17632 8576
rect 17328 8520 17632 8548
rect 17328 8489 17356 8520
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16592 8452 16865 8480
rect 13081 8443 13139 8449
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8480 17095 8483
rect 17129 8483 17187 8489
rect 17129 8480 17141 8483
rect 17083 8452 17141 8480
rect 17083 8449 17095 8452
rect 17037 8443 17095 8449
rect 17129 8449 17141 8452
rect 17175 8449 17187 8483
rect 17129 8443 17187 8449
rect 17277 8483 17356 8489
rect 17277 8449 17289 8483
rect 17323 8452 17356 8483
rect 17323 8449 17335 8452
rect 17277 8443 17335 8449
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 17494 8440 17500 8492
rect 17552 8440 17558 8492
rect 17678 8489 17684 8492
rect 17635 8483 17684 8489
rect 17635 8449 17647 8483
rect 17681 8449 17684 8483
rect 17635 8443 17684 8449
rect 17678 8440 17684 8443
rect 17736 8440 17742 8492
rect 6135 8384 6224 8412
rect 6549 8415 6607 8421
rect 6135 8381 6147 8384
rect 6089 8375 6147 8381
rect 6549 8381 6561 8415
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 6564 8344 6592 8375
rect 6638 8372 6644 8424
rect 6696 8372 6702 8424
rect 6730 8372 6736 8424
rect 6788 8372 6794 8424
rect 7926 8372 7932 8424
rect 7984 8412 7990 8424
rect 8757 8415 8815 8421
rect 8757 8412 8769 8415
rect 7984 8384 8769 8412
rect 7984 8372 7990 8384
rect 8757 8381 8769 8384
rect 8803 8381 8815 8415
rect 8757 8375 8815 8381
rect 8849 8415 8907 8421
rect 8849 8381 8861 8415
rect 8895 8412 8907 8415
rect 9582 8412 9588 8424
rect 8895 8384 9588 8412
rect 8895 8381 8907 8384
rect 8849 8375 8907 8381
rect 4525 8307 4583 8313
rect 4632 8316 5856 8344
rect 5920 8316 6592 8344
rect 4632 8276 4660 8316
rect 4448 8248 4660 8276
rect 5258 8236 5264 8288
rect 5316 8236 5322 8288
rect 5534 8236 5540 8288
rect 5592 8276 5598 8288
rect 5920 8276 5948 8316
rect 5592 8248 5948 8276
rect 5592 8236 5598 8248
rect 6178 8236 6184 8288
rect 6236 8276 6242 8288
rect 6365 8279 6423 8285
rect 6365 8276 6377 8279
rect 6236 8248 6377 8276
rect 6236 8236 6242 8248
rect 6365 8245 6377 8248
rect 6411 8245 6423 8279
rect 6656 8276 6684 8372
rect 6748 8344 6776 8372
rect 8297 8347 8355 8353
rect 8297 8344 8309 8347
rect 6748 8316 8309 8344
rect 8297 8313 8309 8316
rect 8343 8313 8355 8347
rect 8864 8344 8892 8375
rect 9582 8372 9588 8384
rect 9640 8412 9646 8424
rect 9953 8415 10011 8421
rect 9953 8412 9965 8415
rect 9640 8384 9965 8412
rect 9640 8372 9646 8384
rect 9953 8381 9965 8384
rect 9999 8381 10011 8415
rect 13354 8412 13360 8424
rect 9953 8375 10011 8381
rect 12728 8384 13360 8412
rect 12728 8356 12756 8384
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 13446 8372 13452 8424
rect 13504 8372 13510 8424
rect 14090 8372 14096 8424
rect 14148 8412 14154 8424
rect 16669 8415 16727 8421
rect 16669 8412 16681 8415
rect 14148 8384 16681 8412
rect 14148 8372 14154 8384
rect 16669 8381 16681 8384
rect 16715 8381 16727 8415
rect 18524 8412 18552 8576
rect 19242 8548 19248 8560
rect 18892 8520 19248 8548
rect 18892 8489 18920 8520
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8449 18935 8483
rect 21085 8483 21143 8489
rect 18877 8443 18935 8449
rect 19153 8415 19211 8421
rect 19153 8412 19165 8415
rect 18524 8384 19165 8412
rect 16669 8375 16727 8381
rect 19153 8381 19165 8384
rect 19199 8381 19211 8415
rect 19153 8375 19211 8381
rect 8297 8307 8355 8313
rect 8404 8316 8892 8344
rect 8404 8276 8432 8316
rect 12710 8304 12716 8356
rect 12768 8304 12774 8356
rect 13173 8347 13231 8353
rect 13173 8313 13185 8347
rect 13219 8344 13231 8347
rect 18230 8344 18236 8356
rect 13219 8316 13584 8344
rect 13219 8313 13231 8316
rect 13173 8307 13231 8313
rect 6656 8248 8432 8276
rect 13556 8276 13584 8316
rect 16408 8316 18236 8344
rect 16408 8288 16436 8316
rect 18230 8304 18236 8316
rect 18288 8304 18294 8356
rect 20272 8344 20300 8466
rect 21085 8449 21097 8483
rect 21131 8480 21143 8483
rect 21744 8480 21772 8576
rect 23385 8551 23443 8557
rect 23385 8548 23397 8551
rect 22572 8520 23397 8548
rect 22572 8492 22600 8520
rect 23385 8517 23397 8520
rect 23431 8548 23443 8551
rect 23566 8548 23572 8560
rect 23431 8520 23572 8548
rect 23431 8517 23443 8520
rect 23385 8511 23443 8517
rect 23566 8508 23572 8520
rect 23624 8508 23630 8560
rect 25774 8508 25780 8560
rect 25832 8548 25838 8560
rect 26326 8548 26332 8560
rect 25832 8520 26332 8548
rect 25832 8508 25838 8520
rect 26326 8508 26332 8520
rect 26384 8548 26390 8560
rect 27065 8551 27123 8557
rect 27065 8548 27077 8551
rect 26384 8520 27077 8548
rect 26384 8508 26390 8520
rect 27065 8517 27077 8520
rect 27111 8517 27123 8551
rect 27065 8511 27123 8517
rect 21131 8452 21772 8480
rect 21131 8449 21143 8452
rect 21085 8443 21143 8449
rect 22554 8440 22560 8492
rect 22612 8440 22618 8492
rect 22833 8483 22891 8489
rect 22833 8449 22845 8483
rect 22879 8449 22891 8483
rect 22833 8443 22891 8449
rect 22848 8412 22876 8443
rect 23014 8440 23020 8492
rect 23072 8480 23078 8492
rect 23290 8480 23296 8492
rect 23072 8452 23296 8480
rect 23072 8440 23078 8452
rect 23290 8440 23296 8452
rect 23348 8440 23354 8492
rect 23474 8440 23480 8492
rect 23532 8440 23538 8492
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 23676 8452 23949 8480
rect 23106 8412 23112 8424
rect 22848 8384 23112 8412
rect 23106 8372 23112 8384
rect 23164 8412 23170 8424
rect 23382 8412 23388 8424
rect 23164 8384 23388 8412
rect 23164 8372 23170 8384
rect 23382 8372 23388 8384
rect 23440 8412 23446 8424
rect 23676 8412 23704 8452
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 23440 8384 23704 8412
rect 23440 8372 23446 8384
rect 23750 8372 23756 8424
rect 23808 8372 23814 8424
rect 23952 8412 23980 8443
rect 24026 8440 24032 8492
rect 24084 8480 24090 8492
rect 24121 8483 24179 8489
rect 24121 8480 24133 8483
rect 24084 8452 24133 8480
rect 24084 8440 24090 8452
rect 24121 8449 24133 8452
rect 24167 8449 24179 8483
rect 25498 8480 25504 8492
rect 24121 8443 24179 8449
rect 24826 8452 25504 8480
rect 24578 8412 24584 8424
rect 23952 8384 24584 8412
rect 24578 8372 24584 8384
rect 24636 8372 24642 8424
rect 20272 8316 20760 8344
rect 13906 8276 13912 8288
rect 13556 8248 13912 8276
rect 6365 8239 6423 8245
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 16390 8236 16396 8288
rect 16448 8236 16454 8288
rect 17770 8236 17776 8288
rect 17828 8236 17834 8288
rect 20732 8276 20760 8316
rect 23658 8304 23664 8356
rect 23716 8344 23722 8356
rect 23937 8347 23995 8353
rect 23937 8344 23949 8347
rect 23716 8316 23949 8344
rect 23716 8304 23722 8316
rect 23937 8313 23949 8316
rect 23983 8313 23995 8347
rect 24596 8344 24624 8372
rect 24826 8344 24854 8452
rect 25498 8440 25504 8452
rect 25556 8480 25562 8492
rect 26053 8483 26111 8489
rect 26053 8480 26065 8483
rect 25556 8478 25820 8480
rect 25884 8478 26065 8480
rect 25556 8452 26065 8478
rect 25556 8440 25562 8452
rect 25792 8450 25912 8452
rect 26053 8449 26065 8452
rect 26099 8480 26111 8483
rect 26142 8480 26148 8492
rect 26099 8452 26148 8480
rect 26099 8449 26111 8452
rect 26053 8443 26111 8449
rect 26142 8440 26148 8452
rect 26200 8440 26206 8492
rect 26602 8440 26608 8492
rect 26660 8480 26666 8492
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 26660 8452 26985 8480
rect 26660 8440 26666 8452
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 27246 8440 27252 8492
rect 27304 8440 27310 8492
rect 27448 8489 27476 8588
rect 28166 8576 28172 8588
rect 28224 8576 28230 8628
rect 27801 8551 27859 8557
rect 27801 8517 27813 8551
rect 27847 8548 27859 8551
rect 28074 8548 28080 8560
rect 27847 8520 28080 8548
rect 27847 8517 27859 8520
rect 27801 8511 27859 8517
rect 28074 8508 28080 8520
rect 28132 8508 28138 8560
rect 27433 8483 27491 8489
rect 27433 8449 27445 8483
rect 27479 8449 27491 8483
rect 27433 8443 27491 8449
rect 25869 8415 25927 8421
rect 25869 8381 25881 8415
rect 25915 8412 25927 8415
rect 26234 8412 26240 8424
rect 25915 8384 26240 8412
rect 25915 8381 25927 8384
rect 25869 8375 25927 8381
rect 26234 8372 26240 8384
rect 26292 8372 26298 8424
rect 26329 8415 26387 8421
rect 26329 8381 26341 8415
rect 26375 8412 26387 8415
rect 27522 8412 27528 8424
rect 26375 8384 27528 8412
rect 26375 8381 26387 8384
rect 26329 8375 26387 8381
rect 27522 8372 27528 8384
rect 27580 8372 27586 8424
rect 24596 8316 24854 8344
rect 23937 8307 23995 8313
rect 25222 8304 25228 8356
rect 25280 8344 25286 8356
rect 26602 8344 26608 8356
rect 25280 8316 26608 8344
rect 25280 8304 25286 8316
rect 26602 8304 26608 8316
rect 26660 8304 26666 8356
rect 20806 8276 20812 8288
rect 20732 8248 20812 8276
rect 20806 8236 20812 8248
rect 20864 8236 20870 8288
rect 20898 8236 20904 8288
rect 20956 8236 20962 8288
rect 22462 8236 22468 8288
rect 22520 8276 22526 8288
rect 22922 8276 22928 8288
rect 22520 8248 22928 8276
rect 22520 8236 22526 8248
rect 22922 8236 22928 8248
rect 22980 8276 22986 8288
rect 23201 8279 23259 8285
rect 23201 8276 23213 8279
rect 22980 8248 23213 8276
rect 22980 8236 22986 8248
rect 23201 8245 23213 8248
rect 23247 8245 23259 8279
rect 23201 8239 23259 8245
rect 23845 8279 23903 8285
rect 23845 8245 23857 8279
rect 23891 8276 23903 8279
rect 24670 8276 24676 8288
rect 23891 8248 24676 8276
rect 23891 8245 23903 8248
rect 23845 8239 23903 8245
rect 24670 8236 24676 8248
rect 24728 8236 24734 8288
rect 26237 8279 26295 8285
rect 26237 8245 26249 8279
rect 26283 8276 26295 8279
rect 27338 8276 27344 8288
rect 26283 8248 27344 8276
rect 26283 8245 26295 8248
rect 26237 8239 26295 8245
rect 27338 8236 27344 8248
rect 27396 8236 27402 8288
rect 1104 8186 29440 8208
rect 1104 8134 4491 8186
rect 4543 8134 4555 8186
rect 4607 8134 4619 8186
rect 4671 8134 4683 8186
rect 4735 8134 4747 8186
rect 4799 8134 11574 8186
rect 11626 8134 11638 8186
rect 11690 8134 11702 8186
rect 11754 8134 11766 8186
rect 11818 8134 11830 8186
rect 11882 8134 18657 8186
rect 18709 8134 18721 8186
rect 18773 8134 18785 8186
rect 18837 8134 18849 8186
rect 18901 8134 18913 8186
rect 18965 8134 25740 8186
rect 25792 8134 25804 8186
rect 25856 8134 25868 8186
rect 25920 8134 25932 8186
rect 25984 8134 25996 8186
rect 26048 8134 29440 8186
rect 1104 8112 29440 8134
rect 5169 8075 5227 8081
rect 5169 8072 5181 8075
rect 3988 8044 5181 8072
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7936 2007 7939
rect 3988 7936 4016 8044
rect 5169 8041 5181 8044
rect 5215 8041 5227 8075
rect 5169 8035 5227 8041
rect 5537 8075 5595 8081
rect 5537 8041 5549 8075
rect 5583 8072 5595 8075
rect 6089 8075 6147 8081
rect 6089 8072 6101 8075
rect 5583 8044 6101 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 6089 8041 6101 8044
rect 6135 8041 6147 8075
rect 13725 8075 13783 8081
rect 6089 8035 6147 8041
rect 6196 8044 12434 8072
rect 4062 7964 4068 8016
rect 4120 8004 4126 8016
rect 6196 8004 6224 8044
rect 4120 7976 6224 8004
rect 4120 7964 4126 7976
rect 6730 7964 6736 8016
rect 6788 7964 6794 8016
rect 12406 8004 12434 8044
rect 13725 8041 13737 8075
rect 13771 8072 13783 8075
rect 13998 8072 14004 8084
rect 13771 8044 14004 8072
rect 13771 8041 13783 8044
rect 13725 8035 13783 8041
rect 13998 8032 14004 8044
rect 14056 8032 14062 8084
rect 17402 8072 17408 8084
rect 14292 8044 17408 8072
rect 14182 8004 14188 8016
rect 12406 7976 14188 8004
rect 14182 7964 14188 7976
rect 14240 7964 14246 8016
rect 5442 7936 5448 7948
rect 1995 7908 4016 7936
rect 4448 7908 5448 7936
rect 1995 7905 2007 7908
rect 1949 7899 2007 7905
rect 1670 7828 1676 7880
rect 1728 7828 1734 7880
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4448 7868 4476 7908
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 5721 7939 5779 7945
rect 5721 7905 5733 7939
rect 5767 7936 5779 7939
rect 5994 7936 6000 7948
rect 5767 7908 6000 7936
rect 5767 7905 5779 7908
rect 5721 7899 5779 7905
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 6273 7939 6331 7945
rect 6273 7905 6285 7939
rect 6319 7936 6331 7939
rect 7190 7936 7196 7948
rect 6319 7908 7196 7936
rect 6319 7905 6331 7908
rect 6273 7899 6331 7905
rect 7190 7896 7196 7908
rect 7248 7896 7254 7948
rect 12802 7896 12808 7948
rect 12860 7936 12866 7948
rect 14292 7936 14320 8044
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 17678 8072 17684 8084
rect 17512 8044 17684 8072
rect 16574 7964 16580 8016
rect 16632 8004 16638 8016
rect 16632 7976 17080 8004
rect 16632 7964 16638 7976
rect 12860 7908 14320 7936
rect 12860 7896 12866 7908
rect 4019 7840 4476 7868
rect 4525 7871 4583 7877
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4525 7837 4537 7871
rect 4571 7868 4583 7871
rect 4617 7871 4675 7877
rect 4617 7868 4629 7871
rect 4571 7840 4629 7868
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 4617 7837 4629 7840
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 3786 7800 3792 7812
rect 3174 7772 3792 7800
rect 3786 7760 3792 7772
rect 3844 7760 3850 7812
rect 3421 7735 3479 7741
rect 3421 7701 3433 7735
rect 3467 7732 3479 7735
rect 3988 7732 4016 7831
rect 4982 7828 4988 7880
rect 5040 7828 5046 7880
rect 5810 7828 5816 7880
rect 5868 7828 5874 7880
rect 5902 7828 5908 7880
rect 5960 7828 5966 7880
rect 6012 7868 6040 7896
rect 6365 7871 6423 7877
rect 6012 7840 6316 7868
rect 4246 7760 4252 7812
rect 4304 7800 4310 7812
rect 4801 7803 4859 7809
rect 4801 7800 4813 7803
rect 4304 7772 4813 7800
rect 4304 7760 4310 7772
rect 4801 7769 4813 7772
rect 4847 7769 4859 7803
rect 4801 7763 4859 7769
rect 4890 7760 4896 7812
rect 4948 7800 4954 7812
rect 5166 7800 5172 7812
rect 4948 7772 5172 7800
rect 4948 7760 4954 7772
rect 5166 7760 5172 7772
rect 5224 7760 5230 7812
rect 6089 7803 6147 7809
rect 6089 7769 6101 7803
rect 6135 7800 6147 7803
rect 6178 7800 6184 7812
rect 6135 7772 6184 7800
rect 6135 7769 6147 7772
rect 6089 7763 6147 7769
rect 6178 7760 6184 7772
rect 6236 7760 6242 7812
rect 6288 7800 6316 7840
rect 6365 7837 6377 7871
rect 6411 7868 6423 7871
rect 7469 7871 7527 7877
rect 7469 7868 7481 7871
rect 6411 7840 7481 7868
rect 6411 7837 6423 7840
rect 6365 7831 6423 7837
rect 7469 7837 7481 7840
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 13998 7828 14004 7880
rect 14056 7868 14062 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 14056 7840 14105 7868
rect 14056 7828 14062 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7868 14335 7871
rect 14366 7868 14372 7880
rect 14323 7840 14372 7868
rect 14323 7837 14335 7840
rect 14277 7831 14335 7837
rect 6733 7803 6791 7809
rect 6288 7772 6684 7800
rect 3467 7704 4016 7732
rect 3467 7701 3479 7704
rect 3421 7695 3479 7701
rect 6546 7692 6552 7744
rect 6604 7692 6610 7744
rect 6656 7732 6684 7772
rect 6733 7769 6745 7803
rect 6779 7800 6791 7803
rect 6822 7800 6828 7812
rect 6779 7772 6828 7800
rect 6779 7769 6791 7772
rect 6733 7763 6791 7769
rect 6822 7760 6828 7772
rect 6880 7760 6886 7812
rect 7285 7803 7343 7809
rect 7285 7800 7297 7803
rect 6932 7772 7297 7800
rect 6932 7732 6960 7772
rect 7285 7769 7297 7772
rect 7331 7769 7343 7803
rect 7285 7763 7343 7769
rect 13541 7803 13599 7809
rect 13541 7769 13553 7803
rect 13587 7800 13599 7803
rect 13630 7800 13636 7812
rect 13587 7772 13636 7800
rect 13587 7769 13599 7772
rect 13541 7763 13599 7769
rect 13630 7760 13636 7772
rect 13688 7760 13694 7812
rect 13722 7760 13728 7812
rect 13780 7809 13786 7812
rect 13780 7803 13815 7809
rect 13803 7800 13815 7803
rect 14292 7800 14320 7831
rect 14366 7828 14372 7840
rect 14424 7828 14430 7880
rect 14553 7871 14611 7877
rect 14553 7868 14565 7871
rect 14476 7840 14565 7868
rect 13803 7772 14320 7800
rect 13803 7769 13815 7772
rect 13780 7763 13815 7769
rect 13780 7760 13786 7763
rect 6656 7704 6960 7732
rect 7190 7692 7196 7744
rect 7248 7692 7254 7744
rect 13354 7692 13360 7744
rect 13412 7732 13418 7744
rect 13740 7732 13768 7760
rect 14476 7744 14504 7840
rect 14553 7837 14565 7840
rect 14599 7837 14611 7871
rect 14553 7831 14611 7837
rect 14642 7828 14648 7880
rect 14700 7868 14706 7880
rect 14737 7871 14795 7877
rect 14737 7868 14749 7871
rect 14700 7840 14749 7868
rect 14700 7828 14706 7840
rect 14737 7837 14749 7840
rect 14783 7837 14795 7871
rect 14737 7831 14795 7837
rect 15010 7828 15016 7880
rect 15068 7828 15074 7880
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 16390 7868 16396 7880
rect 15528 7840 16396 7868
rect 15528 7828 15534 7840
rect 16390 7828 16396 7840
rect 16448 7828 16454 7880
rect 16574 7828 16580 7880
rect 16632 7828 16638 7880
rect 17052 7877 17080 7976
rect 16853 7871 16911 7877
rect 16853 7837 16865 7871
rect 16899 7837 16911 7871
rect 16853 7831 16911 7837
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 15028 7800 15056 7828
rect 16868 7800 16896 7831
rect 17310 7828 17316 7880
rect 17368 7828 17374 7880
rect 17402 7828 17408 7880
rect 17460 7828 17466 7880
rect 17512 7877 17540 8044
rect 17678 8032 17684 8044
rect 17736 8072 17742 8084
rect 22094 8072 22100 8084
rect 17736 8044 18281 8072
rect 17736 8032 17742 8044
rect 17586 7964 17592 8016
rect 17644 8004 17650 8016
rect 17644 7976 18184 8004
rect 17644 7964 17650 7976
rect 17604 7908 18092 7936
rect 17497 7871 17555 7877
rect 17497 7837 17509 7871
rect 17543 7837 17555 7871
rect 17497 7831 17555 7837
rect 15028 7772 16896 7800
rect 17218 7760 17224 7812
rect 17276 7760 17282 7812
rect 17328 7800 17356 7828
rect 17604 7800 17632 7908
rect 17954 7877 17960 7880
rect 17773 7871 17831 7877
rect 17773 7868 17785 7871
rect 17328 7772 17632 7800
rect 17696 7840 17785 7868
rect 13412 7704 13768 7732
rect 13412 7692 13418 7704
rect 13906 7692 13912 7744
rect 13964 7692 13970 7744
rect 14458 7692 14464 7744
rect 14516 7692 14522 7744
rect 14642 7692 14648 7744
rect 14700 7692 14706 7744
rect 16758 7692 16764 7744
rect 16816 7732 16822 7744
rect 17696 7732 17724 7840
rect 17773 7837 17785 7840
rect 17819 7837 17831 7871
rect 17773 7831 17831 7837
rect 17921 7871 17960 7877
rect 17921 7837 17933 7871
rect 17921 7831 17960 7837
rect 17954 7828 17960 7831
rect 18012 7828 18018 7880
rect 18064 7877 18092 7908
rect 18156 7877 18184 7976
rect 18253 7877 18281 8044
rect 19260 8044 22100 8072
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 18238 7871 18296 7877
rect 18238 7837 18250 7871
rect 18284 7837 18296 7871
rect 18238 7831 18296 7837
rect 18156 7800 18184 7831
rect 19260 7800 19288 8044
rect 22094 8032 22100 8044
rect 22152 8032 22158 8084
rect 22186 8032 22192 8084
rect 22244 8072 22250 8084
rect 22373 8075 22431 8081
rect 22373 8072 22385 8075
rect 22244 8044 22385 8072
rect 22244 8032 22250 8044
rect 22373 8041 22385 8044
rect 22419 8041 22431 8075
rect 23201 8075 23259 8081
rect 23201 8072 23213 8075
rect 22373 8035 22431 8041
rect 22480 8044 22692 8072
rect 22480 8004 22508 8044
rect 22020 7976 22508 8004
rect 22664 8004 22692 8044
rect 22940 8044 23213 8072
rect 22940 8004 22968 8044
rect 23201 8041 23213 8044
rect 23247 8072 23259 8075
rect 23474 8072 23480 8084
rect 23247 8044 23480 8072
rect 23247 8041 23259 8044
rect 23201 8035 23259 8041
rect 23474 8032 23480 8044
rect 23532 8032 23538 8084
rect 25222 8032 25228 8084
rect 25280 8032 25286 8084
rect 26142 8072 26148 8084
rect 25516 8044 26148 8072
rect 23566 8004 23572 8016
rect 22664 7976 22968 8004
rect 23492 7976 23572 8004
rect 20349 7939 20407 7945
rect 20349 7905 20361 7939
rect 20395 7936 20407 7939
rect 20898 7936 20904 7948
rect 20395 7908 20904 7936
rect 20395 7905 20407 7908
rect 20349 7899 20407 7905
rect 20898 7896 20904 7908
rect 20956 7896 20962 7948
rect 20070 7828 20076 7880
rect 20128 7828 20134 7880
rect 22020 7877 22048 7976
rect 22462 7936 22468 7948
rect 22388 7908 22468 7936
rect 22005 7871 22063 7877
rect 22005 7837 22017 7871
rect 22051 7837 22063 7871
rect 22278 7868 22284 7880
rect 22005 7831 22063 7837
rect 22112 7840 22284 7868
rect 18156 7772 19288 7800
rect 20806 7760 20812 7812
rect 20864 7760 20870 7812
rect 22112 7744 22140 7840
rect 22278 7828 22284 7840
rect 22336 7828 22342 7880
rect 22189 7803 22247 7809
rect 22189 7769 22201 7803
rect 22235 7800 22247 7803
rect 22388 7800 22416 7908
rect 22462 7896 22468 7908
rect 22520 7896 22526 7948
rect 22554 7828 22560 7880
rect 22612 7828 22618 7880
rect 22830 7828 22836 7880
rect 22888 7877 22894 7880
rect 23014 7877 23020 7882
rect 22888 7871 22937 7877
rect 22888 7837 22891 7871
rect 22925 7837 22937 7871
rect 22888 7831 22937 7837
rect 22971 7871 23020 7877
rect 22971 7837 22983 7871
rect 23017 7837 23020 7871
rect 22971 7831 23020 7837
rect 22888 7828 22894 7831
rect 23014 7830 23020 7831
rect 23072 7830 23078 7882
rect 23106 7828 23112 7880
rect 23164 7877 23170 7880
rect 23164 7868 23173 7877
rect 23164 7840 23209 7868
rect 23164 7831 23173 7840
rect 23164 7828 23170 7831
rect 23290 7828 23296 7880
rect 23348 7828 23354 7880
rect 22235 7772 22416 7800
rect 22235 7769 22247 7772
rect 22189 7763 22247 7769
rect 22646 7760 22652 7812
rect 22704 7760 22710 7812
rect 22741 7803 22799 7809
rect 22741 7769 22753 7803
rect 22787 7769 22799 7803
rect 22741 7763 22799 7769
rect 16816 7704 17724 7732
rect 16816 7692 16822 7704
rect 18322 7692 18328 7744
rect 18380 7732 18386 7744
rect 18417 7735 18475 7741
rect 18417 7732 18429 7735
rect 18380 7704 18429 7732
rect 18380 7692 18386 7704
rect 18417 7701 18429 7704
rect 18463 7701 18475 7735
rect 18417 7695 18475 7701
rect 21821 7735 21879 7741
rect 21821 7701 21833 7735
rect 21867 7732 21879 7735
rect 22094 7732 22100 7744
rect 21867 7704 22100 7732
rect 21867 7701 21879 7704
rect 21821 7695 21879 7701
rect 22094 7692 22100 7704
rect 22152 7692 22158 7744
rect 22281 7735 22339 7741
rect 22281 7701 22293 7735
rect 22327 7732 22339 7735
rect 22462 7732 22468 7744
rect 22327 7704 22468 7732
rect 22327 7701 22339 7704
rect 22281 7695 22339 7701
rect 22462 7692 22468 7704
rect 22520 7692 22526 7744
rect 22756 7732 22784 7763
rect 23382 7760 23388 7812
rect 23440 7760 23446 7812
rect 23492 7800 23520 7976
rect 23566 7964 23572 7976
rect 23624 7964 23630 8016
rect 24026 7964 24032 8016
rect 24084 8004 24090 8016
rect 25516 8004 25544 8044
rect 26142 8032 26148 8044
rect 26200 8032 26206 8084
rect 27338 8032 27344 8084
rect 27396 8072 27402 8084
rect 27617 8075 27675 8081
rect 27617 8072 27629 8075
rect 27396 8044 27629 8072
rect 27396 8032 27402 8044
rect 27617 8041 27629 8044
rect 27663 8072 27675 8075
rect 28074 8072 28080 8084
rect 27663 8044 28080 8072
rect 27663 8041 27675 8044
rect 27617 8035 27675 8041
rect 28074 8032 28080 8044
rect 28132 8032 28138 8084
rect 27801 8007 27859 8013
rect 27801 8004 27813 8007
rect 24084 7976 25544 8004
rect 25884 7976 27813 8004
rect 24084 7964 24090 7976
rect 23584 7908 23888 7936
rect 23584 7880 23612 7908
rect 23566 7828 23572 7880
rect 23624 7828 23630 7880
rect 23658 7828 23664 7880
rect 23716 7828 23722 7880
rect 23750 7828 23756 7880
rect 23808 7828 23814 7880
rect 23860 7877 23888 7908
rect 23934 7896 23940 7948
rect 23992 7936 23998 7948
rect 24765 7939 24823 7945
rect 24765 7936 24777 7939
rect 23992 7908 24777 7936
rect 23992 7896 23998 7908
rect 24765 7905 24777 7908
rect 24811 7936 24823 7939
rect 24811 7908 25084 7936
rect 24811 7905 24823 7908
rect 24765 7899 24823 7905
rect 23845 7871 23903 7877
rect 23845 7837 23857 7871
rect 23891 7837 23903 7871
rect 23845 7831 23903 7837
rect 24029 7871 24087 7877
rect 24029 7837 24041 7871
rect 24075 7837 24087 7871
rect 24029 7831 24087 7837
rect 24044 7800 24072 7831
rect 24118 7828 24124 7880
rect 24176 7868 24182 7880
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 24176 7840 24409 7868
rect 24176 7828 24182 7840
rect 24397 7837 24409 7840
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 24578 7828 24584 7880
rect 24636 7828 24642 7880
rect 24670 7828 24676 7880
rect 24728 7868 24734 7880
rect 25056 7877 25084 7908
rect 24857 7871 24915 7877
rect 24857 7868 24869 7871
rect 24728 7840 24869 7868
rect 24728 7828 24734 7840
rect 24857 7837 24869 7840
rect 24903 7837 24915 7871
rect 24857 7831 24915 7837
rect 25041 7871 25099 7877
rect 25041 7837 25053 7871
rect 25087 7837 25099 7871
rect 25041 7831 25099 7837
rect 25777 7871 25835 7877
rect 25777 7837 25789 7871
rect 25823 7868 25835 7871
rect 25884 7868 25912 7976
rect 27801 7973 27813 7976
rect 27847 7973 27859 8007
rect 27801 7967 27859 7973
rect 26142 7896 26148 7948
rect 26200 7896 26206 7948
rect 26237 7939 26295 7945
rect 26237 7905 26249 7939
rect 26283 7936 26295 7939
rect 27157 7939 27215 7945
rect 27157 7936 27169 7939
rect 26283 7908 27169 7936
rect 26283 7905 26295 7908
rect 26237 7899 26295 7905
rect 27157 7905 27169 7908
rect 27203 7905 27215 7939
rect 27157 7899 27215 7905
rect 27522 7896 27528 7948
rect 27580 7896 27586 7948
rect 25823 7840 25912 7868
rect 25961 7871 26019 7877
rect 25823 7837 25835 7840
rect 25777 7831 25835 7837
rect 25961 7837 25973 7871
rect 26007 7868 26019 7871
rect 26160 7868 26188 7896
rect 26007 7840 26188 7868
rect 26513 7871 26571 7877
rect 26007 7837 26019 7840
rect 25961 7831 26019 7837
rect 26513 7837 26525 7871
rect 26559 7837 26571 7871
rect 26513 7831 26571 7837
rect 23492 7772 24072 7800
rect 24302 7760 24308 7812
rect 24360 7800 24366 7812
rect 24360 7772 25820 7800
rect 24360 7760 24366 7772
rect 24026 7732 24032 7744
rect 22756 7704 24032 7732
rect 24026 7692 24032 7704
rect 24084 7692 24090 7744
rect 25590 7692 25596 7744
rect 25648 7692 25654 7744
rect 25792 7732 25820 7772
rect 25866 7760 25872 7812
rect 25924 7760 25930 7812
rect 26079 7803 26137 7809
rect 26079 7800 26091 7803
rect 25976 7772 26091 7800
rect 25976 7732 26004 7772
rect 26079 7769 26091 7772
rect 26125 7769 26137 7803
rect 26079 7763 26137 7769
rect 26234 7760 26240 7812
rect 26292 7800 26298 7812
rect 26528 7800 26556 7831
rect 26602 7828 26608 7880
rect 26660 7868 26666 7880
rect 27249 7871 27307 7877
rect 27249 7868 27261 7871
rect 26660 7840 27261 7868
rect 26660 7828 26666 7840
rect 27249 7837 27261 7840
rect 27295 7837 27307 7871
rect 27249 7831 27307 7837
rect 26292 7772 26556 7800
rect 26292 7760 26298 7772
rect 26418 7732 26424 7744
rect 25792 7704 26424 7732
rect 26418 7692 26424 7704
rect 26476 7692 26482 7744
rect 1104 7642 29595 7664
rect 1104 7590 8032 7642
rect 8084 7590 8096 7642
rect 8148 7590 8160 7642
rect 8212 7590 8224 7642
rect 8276 7590 8288 7642
rect 8340 7590 15115 7642
rect 15167 7590 15179 7642
rect 15231 7590 15243 7642
rect 15295 7590 15307 7642
rect 15359 7590 15371 7642
rect 15423 7590 22198 7642
rect 22250 7590 22262 7642
rect 22314 7590 22326 7642
rect 22378 7590 22390 7642
rect 22442 7590 22454 7642
rect 22506 7590 29281 7642
rect 29333 7590 29345 7642
rect 29397 7590 29409 7642
rect 29461 7590 29473 7642
rect 29525 7590 29537 7642
rect 29589 7590 29595 7642
rect 1104 7568 29595 7590
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 5629 7531 5687 7537
rect 5629 7528 5641 7531
rect 5316 7500 5641 7528
rect 5316 7488 5322 7500
rect 5629 7497 5641 7500
rect 5675 7497 5687 7531
rect 5629 7491 5687 7497
rect 5810 7488 5816 7540
rect 5868 7488 5874 7540
rect 6546 7488 6552 7540
rect 6604 7528 6610 7540
rect 12802 7528 12808 7540
rect 6604 7500 12808 7528
rect 6604 7488 6610 7500
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 14642 7528 14648 7540
rect 12912 7500 14648 7528
rect 5828 7460 5856 7488
rect 11517 7463 11575 7469
rect 11517 7460 11529 7463
rect 5828 7432 6132 7460
rect 5997 7395 6055 7401
rect 5997 7392 6009 7395
rect 5736 7364 6009 7392
rect 5736 7336 5764 7364
rect 5997 7361 6009 7364
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 5718 7284 5724 7336
rect 5776 7284 5782 7336
rect 5813 7327 5871 7333
rect 5813 7293 5825 7327
rect 5859 7293 5871 7327
rect 5813 7287 5871 7293
rect 5905 7327 5963 7333
rect 5905 7293 5917 7327
rect 5951 7324 5963 7327
rect 6104 7324 6132 7432
rect 10336 7432 11529 7460
rect 10336 7401 10364 7432
rect 11517 7429 11529 7432
rect 11563 7429 11575 7463
rect 12710 7460 12716 7472
rect 11517 7423 11575 7429
rect 11808 7432 12716 7460
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 10502 7352 10508 7404
rect 10560 7392 10566 7404
rect 10597 7395 10655 7401
rect 10597 7392 10609 7395
rect 10560 7364 10609 7392
rect 10560 7352 10566 7364
rect 10597 7361 10609 7364
rect 10643 7361 10655 7395
rect 10597 7355 10655 7361
rect 10873 7395 10931 7401
rect 10873 7361 10885 7395
rect 10919 7392 10931 7395
rect 11330 7392 11336 7404
rect 10919 7364 11336 7392
rect 10919 7361 10931 7364
rect 10873 7355 10931 7361
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 11808 7401 11836 7432
rect 12710 7420 12716 7432
rect 12768 7420 12774 7472
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7361 11851 7395
rect 11793 7355 11851 7361
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 12253 7395 12311 7401
rect 12253 7392 12265 7395
rect 12124 7364 12265 7392
rect 12124 7352 12130 7364
rect 12253 7361 12265 7364
rect 12299 7361 12311 7395
rect 12912 7392 12940 7500
rect 14642 7488 14648 7500
rect 14700 7488 14706 7540
rect 16758 7488 16764 7540
rect 16816 7488 16822 7540
rect 16850 7488 16856 7540
rect 16908 7528 16914 7540
rect 16945 7531 17003 7537
rect 16945 7528 16957 7531
rect 16908 7500 16957 7528
rect 16908 7488 16914 7500
rect 16945 7497 16957 7500
rect 16991 7497 17003 7531
rect 17954 7528 17960 7540
rect 16945 7491 17003 7497
rect 17292 7500 17960 7528
rect 12989 7463 13047 7469
rect 12989 7429 13001 7463
rect 13035 7460 13047 7463
rect 13817 7463 13875 7469
rect 13817 7460 13829 7463
rect 13035 7432 13829 7460
rect 13035 7429 13047 7432
rect 12989 7423 13047 7429
rect 13817 7429 13829 7432
rect 13863 7429 13875 7463
rect 13817 7423 13875 7429
rect 14274 7420 14280 7472
rect 14332 7420 14338 7472
rect 16776 7460 16804 7488
rect 16776 7432 17172 7460
rect 13173 7395 13231 7401
rect 13173 7392 13185 7395
rect 12912 7364 13185 7392
rect 12253 7355 12311 7361
rect 13173 7361 13185 7364
rect 13219 7361 13231 7395
rect 13173 7355 13231 7361
rect 13354 7352 13360 7404
rect 13412 7352 13418 7404
rect 13538 7352 13544 7404
rect 13596 7352 13602 7404
rect 16761 7395 16819 7401
rect 16761 7361 16773 7395
rect 16807 7361 16819 7395
rect 16761 7355 16819 7361
rect 5951 7296 6132 7324
rect 11057 7327 11115 7333
rect 5951 7293 5963 7296
rect 5905 7287 5963 7293
rect 11057 7293 11069 7327
rect 11103 7293 11115 7327
rect 11057 7287 11115 7293
rect 4982 7216 4988 7268
rect 5040 7216 5046 7268
rect 5828 7256 5856 7287
rect 5994 7256 6000 7268
rect 5828 7228 6000 7256
rect 5994 7216 6000 7228
rect 6052 7216 6058 7268
rect 5000 7188 5028 7216
rect 11072 7188 11100 7287
rect 11146 7284 11152 7336
rect 11204 7284 11210 7336
rect 13449 7327 13507 7333
rect 13449 7293 13461 7327
rect 13495 7293 13507 7327
rect 15010 7324 15016 7336
rect 13449 7287 13507 7293
rect 14844 7296 15016 7324
rect 11164 7256 11192 7284
rect 12069 7259 12127 7265
rect 12069 7256 12081 7259
rect 11164 7228 12081 7256
rect 12069 7225 12081 7228
rect 12115 7225 12127 7259
rect 12069 7219 12127 7225
rect 5000 7160 11100 7188
rect 11422 7148 11428 7200
rect 11480 7188 11486 7200
rect 11885 7191 11943 7197
rect 11885 7188 11897 7191
rect 11480 7160 11897 7188
rect 11480 7148 11486 7160
rect 11885 7157 11897 7160
rect 11931 7157 11943 7191
rect 11885 7151 11943 7157
rect 11974 7148 11980 7200
rect 12032 7148 12038 7200
rect 13464 7188 13492 7287
rect 13998 7188 14004 7200
rect 13464 7160 14004 7188
rect 13998 7148 14004 7160
rect 14056 7188 14062 7200
rect 14844 7188 14872 7296
rect 15010 7284 15016 7296
rect 15068 7324 15074 7336
rect 15565 7327 15623 7333
rect 15565 7324 15577 7327
rect 15068 7296 15577 7324
rect 15068 7284 15074 7296
rect 15565 7293 15577 7296
rect 15611 7293 15623 7327
rect 16776 7324 16804 7355
rect 17034 7352 17040 7404
rect 17092 7352 17098 7404
rect 17144 7401 17172 7432
rect 17292 7401 17320 7500
rect 17954 7488 17960 7500
rect 18012 7488 18018 7540
rect 22557 7531 22615 7537
rect 22557 7497 22569 7531
rect 22603 7528 22615 7531
rect 22646 7528 22652 7540
rect 22603 7500 22652 7528
rect 22603 7497 22615 7500
rect 22557 7491 22615 7497
rect 22646 7488 22652 7500
rect 22704 7488 22710 7540
rect 22922 7488 22928 7540
rect 22980 7488 22986 7540
rect 23014 7488 23020 7540
rect 23072 7488 23078 7540
rect 23382 7488 23388 7540
rect 23440 7528 23446 7540
rect 23440 7500 24716 7528
rect 23440 7488 23446 7500
rect 18325 7463 18383 7469
rect 18325 7460 18337 7463
rect 18156 7432 18337 7460
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7361 17187 7395
rect 17129 7355 17187 7361
rect 17277 7395 17335 7401
rect 17277 7361 17289 7395
rect 17323 7361 17335 7395
rect 17277 7355 17335 7361
rect 17402 7352 17408 7404
rect 17460 7352 17466 7404
rect 17494 7352 17500 7404
rect 17552 7352 17558 7404
rect 17589 7395 17647 7401
rect 17589 7361 17601 7395
rect 17635 7392 17647 7395
rect 17678 7392 17684 7404
rect 17635 7364 17684 7392
rect 17635 7361 17647 7364
rect 17589 7355 17647 7361
rect 17678 7352 17684 7364
rect 17736 7352 17742 7404
rect 17862 7352 17868 7404
rect 17920 7352 17926 7404
rect 18046 7352 18052 7404
rect 18104 7352 18110 7404
rect 18156 7324 18184 7432
rect 18325 7429 18337 7432
rect 18371 7429 18383 7463
rect 18325 7423 18383 7429
rect 22465 7463 22523 7469
rect 22465 7429 22477 7463
rect 22511 7460 22523 7463
rect 23032 7460 23060 7488
rect 22511 7432 23060 7460
rect 22511 7429 22523 7432
rect 22465 7423 22523 7429
rect 23474 7420 23480 7472
rect 23532 7420 23538 7472
rect 23753 7463 23811 7469
rect 23753 7429 23765 7463
rect 23799 7460 23811 7463
rect 24121 7463 24179 7469
rect 24121 7460 24133 7463
rect 23799 7432 24133 7460
rect 23799 7429 23811 7432
rect 23753 7423 23811 7429
rect 24121 7429 24133 7432
rect 24167 7429 24179 7463
rect 24121 7423 24179 7429
rect 24578 7420 24584 7472
rect 24636 7420 24642 7472
rect 18233 7395 18291 7401
rect 18233 7361 18245 7395
rect 18279 7361 18291 7395
rect 18233 7355 18291 7361
rect 18417 7395 18475 7401
rect 18417 7361 18429 7395
rect 18463 7361 18475 7395
rect 18417 7355 18475 7361
rect 16776 7296 18184 7324
rect 15565 7287 15623 7293
rect 17034 7216 17040 7268
rect 17092 7256 17098 7268
rect 17770 7256 17776 7268
rect 17092 7228 17776 7256
rect 17092 7216 17098 7228
rect 17770 7216 17776 7228
rect 17828 7256 17834 7268
rect 18248 7256 18276 7355
rect 18432 7256 18460 7355
rect 22094 7352 22100 7404
rect 22152 7392 22158 7404
rect 22741 7395 22799 7401
rect 22741 7392 22753 7395
rect 22152 7364 22753 7392
rect 22152 7352 22158 7364
rect 22741 7361 22753 7364
rect 22787 7361 22799 7395
rect 22741 7355 22799 7361
rect 23017 7395 23075 7401
rect 23017 7361 23029 7395
rect 23063 7392 23075 7395
rect 23492 7392 23520 7420
rect 23063 7364 23520 7392
rect 23845 7395 23903 7401
rect 23063 7361 23075 7364
rect 23017 7355 23075 7361
rect 23845 7361 23857 7395
rect 23891 7361 23903 7395
rect 23845 7355 23903 7361
rect 21913 7327 21971 7333
rect 21913 7293 21925 7327
rect 21959 7324 21971 7327
rect 22278 7324 22284 7336
rect 21959 7296 22284 7324
rect 21959 7293 21971 7296
rect 21913 7287 21971 7293
rect 22278 7284 22284 7296
rect 22336 7324 22342 7336
rect 23106 7324 23112 7336
rect 22336 7296 23112 7324
rect 22336 7284 22342 7296
rect 23106 7284 23112 7296
rect 23164 7284 23170 7336
rect 23201 7327 23259 7333
rect 23201 7293 23213 7327
rect 23247 7293 23259 7327
rect 23860 7324 23888 7355
rect 24026 7352 24032 7404
rect 24084 7352 24090 7404
rect 24213 7398 24271 7401
rect 24302 7398 24308 7404
rect 24213 7395 24308 7398
rect 24213 7361 24225 7395
rect 24259 7370 24308 7395
rect 24259 7361 24271 7370
rect 24213 7355 24271 7361
rect 24302 7352 24308 7370
rect 24360 7352 24366 7404
rect 24489 7395 24547 7401
rect 24489 7361 24501 7395
rect 24535 7392 24547 7395
rect 24596 7392 24624 7420
rect 24688 7401 24716 7500
rect 25590 7488 25596 7540
rect 25648 7488 25654 7540
rect 25866 7488 25872 7540
rect 25924 7528 25930 7540
rect 27157 7531 27215 7537
rect 27157 7528 27169 7531
rect 25924 7500 27169 7528
rect 25924 7488 25930 7500
rect 27157 7497 27169 7500
rect 27203 7497 27215 7531
rect 27157 7491 27215 7497
rect 27522 7488 27528 7540
rect 27580 7528 27586 7540
rect 27617 7531 27675 7537
rect 27617 7528 27629 7531
rect 27580 7500 27629 7528
rect 27580 7488 27586 7500
rect 27617 7497 27629 7500
rect 27663 7497 27675 7531
rect 27617 7491 27675 7497
rect 25225 7463 25283 7469
rect 25225 7429 25237 7463
rect 25271 7460 25283 7463
rect 25608 7460 25636 7488
rect 26510 7460 26516 7472
rect 25271 7432 25636 7460
rect 26450 7432 26516 7460
rect 25271 7429 25283 7432
rect 25225 7423 25283 7429
rect 26510 7420 26516 7432
rect 26568 7460 26574 7472
rect 27062 7460 27068 7472
rect 26568 7432 27068 7460
rect 26568 7420 26574 7432
rect 27062 7420 27068 7432
rect 27120 7420 27126 7472
rect 27540 7460 27568 7488
rect 27448 7432 27568 7460
rect 27632 7432 27844 7460
rect 24535 7364 24624 7392
rect 24673 7395 24731 7401
rect 24535 7361 24547 7364
rect 24489 7355 24547 7361
rect 24673 7361 24685 7395
rect 24719 7361 24731 7395
rect 24673 7355 24731 7361
rect 24946 7352 24952 7404
rect 25004 7352 25010 7404
rect 26234 7352 26240 7404
rect 26292 7352 26298 7404
rect 26602 7352 26608 7404
rect 26660 7392 26666 7404
rect 26973 7395 27031 7401
rect 26973 7392 26985 7395
rect 26660 7364 26985 7392
rect 26660 7352 26666 7364
rect 26973 7361 26985 7364
rect 27019 7361 27031 7395
rect 26973 7355 27031 7361
rect 27249 7395 27307 7401
rect 27249 7361 27261 7395
rect 27295 7392 27307 7395
rect 27338 7392 27344 7404
rect 27295 7364 27344 7392
rect 27295 7361 27307 7364
rect 27249 7355 27307 7361
rect 27338 7352 27344 7364
rect 27396 7352 27402 7404
rect 27448 7401 27476 7432
rect 27433 7395 27491 7401
rect 27433 7361 27445 7395
rect 27479 7361 27491 7395
rect 27433 7355 27491 7361
rect 27525 7395 27583 7401
rect 27525 7361 27537 7395
rect 27571 7392 27583 7395
rect 27632 7392 27660 7432
rect 27816 7404 27844 7432
rect 27571 7364 27660 7392
rect 27709 7395 27767 7401
rect 27571 7361 27583 7364
rect 27525 7355 27583 7361
rect 27709 7361 27721 7395
rect 27755 7361 27767 7395
rect 27709 7355 27767 7361
rect 26252 7324 26280 7352
rect 26697 7327 26755 7333
rect 26697 7324 26709 7327
rect 23860 7296 24164 7324
rect 26252 7296 26709 7324
rect 23201 7287 23259 7293
rect 17828 7228 18276 7256
rect 18340 7228 18460 7256
rect 17828 7216 17834 7228
rect 18340 7200 18368 7228
rect 14056 7160 14872 7188
rect 14056 7148 14062 7160
rect 16758 7148 16764 7200
rect 16816 7148 16822 7200
rect 17129 7191 17187 7197
rect 17129 7157 17141 7191
rect 17175 7188 17187 7191
rect 17402 7188 17408 7200
rect 17175 7160 17408 7188
rect 17175 7157 17187 7160
rect 17129 7151 17187 7157
rect 17402 7148 17408 7160
rect 17460 7148 17466 7200
rect 17862 7148 17868 7200
rect 17920 7148 17926 7200
rect 18322 7148 18328 7200
rect 18380 7148 18386 7200
rect 23216 7188 23244 7287
rect 24136 7256 24164 7296
rect 26697 7293 26709 7296
rect 26743 7324 26755 7327
rect 26743 7296 27614 7324
rect 26743 7293 26755 7296
rect 26697 7287 26755 7293
rect 24489 7259 24547 7265
rect 24489 7256 24501 7259
rect 24136 7228 24501 7256
rect 24489 7225 24501 7228
rect 24535 7225 24547 7259
rect 27586 7256 27614 7296
rect 27724 7256 27752 7355
rect 27798 7352 27804 7404
rect 27856 7352 27862 7404
rect 28718 7352 28724 7404
rect 28776 7352 28782 7404
rect 27586 7228 27752 7256
rect 24489 7219 24547 7225
rect 24118 7188 24124 7200
rect 23216 7160 24124 7188
rect 24118 7148 24124 7160
rect 24176 7148 24182 7200
rect 24394 7148 24400 7200
rect 24452 7148 24458 7200
rect 28994 7148 29000 7200
rect 29052 7148 29058 7200
rect 1104 7098 29440 7120
rect 1104 7046 4491 7098
rect 4543 7046 4555 7098
rect 4607 7046 4619 7098
rect 4671 7046 4683 7098
rect 4735 7046 4747 7098
rect 4799 7046 11574 7098
rect 11626 7046 11638 7098
rect 11690 7046 11702 7098
rect 11754 7046 11766 7098
rect 11818 7046 11830 7098
rect 11882 7046 18657 7098
rect 18709 7046 18721 7098
rect 18773 7046 18785 7098
rect 18837 7046 18849 7098
rect 18901 7046 18913 7098
rect 18965 7046 25740 7098
rect 25792 7046 25804 7098
rect 25856 7046 25868 7098
rect 25920 7046 25932 7098
rect 25984 7046 25996 7098
rect 26048 7046 29440 7098
rect 1104 7024 29440 7046
rect 4982 6944 4988 6996
rect 5040 6984 5046 6996
rect 5040 6956 8156 6984
rect 5040 6944 5046 6956
rect 4816 6888 6224 6916
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6780 4583 6783
rect 4614 6780 4620 6792
rect 4571 6752 4620 6780
rect 4571 6749 4583 6752
rect 4525 6743 4583 6749
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6780 4767 6783
rect 4816 6780 4844 6888
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6848 5411 6851
rect 5902 6848 5908 6860
rect 5399 6820 5908 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 6196 6792 6224 6888
rect 4755 6752 4844 6780
rect 4893 6783 4951 6789
rect 4755 6749 4767 6752
rect 4709 6743 4767 6749
rect 4893 6749 4905 6783
rect 4939 6780 4951 6783
rect 4982 6780 4988 6792
rect 4939 6752 4988 6780
rect 4939 6749 4951 6752
rect 4893 6743 4951 6749
rect 4982 6740 4988 6752
rect 5040 6740 5046 6792
rect 5074 6740 5080 6792
rect 5132 6780 5138 6792
rect 5994 6780 6000 6792
rect 5132 6752 6000 6780
rect 5132 6740 5138 6752
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 6178 6740 6184 6792
rect 6236 6740 6242 6792
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6780 6423 6783
rect 6748 6780 6776 6956
rect 7558 6916 7564 6928
rect 7024 6888 7564 6916
rect 6411 6752 6776 6780
rect 6411 6749 6423 6752
rect 6365 6743 6423 6749
rect 6822 6740 6828 6792
rect 6880 6740 6886 6792
rect 7024 6789 7052 6888
rect 7558 6876 7564 6888
rect 7616 6876 7622 6928
rect 8021 6919 8079 6925
rect 8021 6885 8033 6919
rect 8067 6885 8079 6919
rect 8021 6879 8079 6885
rect 7282 6808 7288 6860
rect 7340 6848 7346 6860
rect 8036 6848 8064 6879
rect 7340 6820 8064 6848
rect 8128 6848 8156 6956
rect 10502 6944 10508 6996
rect 10560 6944 10566 6996
rect 10594 6944 10600 6996
rect 10652 6984 10658 6996
rect 11149 6987 11207 6993
rect 11149 6984 11161 6987
rect 10652 6956 11161 6984
rect 10652 6944 10658 6956
rect 11149 6953 11161 6956
rect 11195 6984 11207 6987
rect 11238 6984 11244 6996
rect 11195 6956 11244 6984
rect 11195 6953 11207 6956
rect 11149 6947 11207 6953
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 11330 6944 11336 6996
rect 11388 6944 11394 6996
rect 11514 6944 11520 6996
rect 11572 6984 11578 6996
rect 12066 6984 12072 6996
rect 11572 6956 12072 6984
rect 11572 6944 11578 6956
rect 12066 6944 12072 6956
rect 12124 6944 12130 6996
rect 13630 6944 13636 6996
rect 13688 6984 13694 6996
rect 13688 6956 14136 6984
rect 13688 6944 13694 6956
rect 10520 6916 10548 6944
rect 9692 6888 10548 6916
rect 11256 6916 11284 6944
rect 12161 6919 12219 6925
rect 12161 6916 12173 6919
rect 11256 6888 12173 6916
rect 9692 6848 9720 6888
rect 12161 6885 12173 6888
rect 12207 6885 12219 6919
rect 12161 6879 12219 6885
rect 11422 6848 11428 6860
rect 8128 6820 9720 6848
rect 9968 6820 11428 6848
rect 7340 6808 7346 6820
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6749 7067 6783
rect 7009 6743 7067 6749
rect 7193 6783 7251 6789
rect 7193 6749 7205 6783
rect 7239 6780 7251 6783
rect 7374 6780 7380 6792
rect 7239 6752 7380 6780
rect 7239 6749 7251 6752
rect 7193 6743 7251 6749
rect 7374 6740 7380 6752
rect 7432 6740 7438 6792
rect 7466 6740 7472 6792
rect 7524 6740 7530 6792
rect 7558 6740 7564 6792
rect 7616 6780 7622 6792
rect 7653 6783 7711 6789
rect 7653 6780 7665 6783
rect 7616 6752 7665 6780
rect 7616 6740 7622 6752
rect 7653 6749 7665 6752
rect 7699 6749 7711 6783
rect 7653 6743 7711 6749
rect 7834 6740 7840 6792
rect 7892 6740 7898 6792
rect 9968 6789 9996 6820
rect 11422 6808 11428 6820
rect 11480 6808 11486 6860
rect 11698 6848 11704 6860
rect 11624 6820 11704 6848
rect 9953 6783 10011 6789
rect 9953 6749 9965 6783
rect 9999 6749 10011 6783
rect 9953 6743 10011 6749
rect 10042 6740 10048 6792
rect 10100 6740 10106 6792
rect 10134 6740 10140 6792
rect 10192 6740 10198 6792
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6780 10839 6783
rect 10962 6780 10968 6792
rect 10827 6752 10968 6780
rect 10827 6749 10839 6752
rect 10781 6743 10839 6749
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 11624 6789 11652 6820
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 11790 6808 11796 6860
rect 11848 6848 11854 6860
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 11848 6820 11989 6848
rect 11848 6808 11854 6820
rect 11977 6817 11989 6820
rect 12023 6817 12035 6851
rect 11977 6811 12035 6817
rect 11609 6783 11667 6789
rect 11609 6749 11621 6783
rect 11655 6749 11667 6783
rect 11609 6743 11667 6749
rect 12066 6740 12072 6792
rect 12124 6740 12130 6792
rect 4801 6715 4859 6721
rect 4801 6681 4813 6715
rect 4847 6712 4859 6715
rect 4847 6684 5304 6712
rect 4847 6681 4859 6684
rect 4801 6675 4859 6681
rect 5074 6604 5080 6656
rect 5132 6604 5138 6656
rect 5276 6644 5304 6684
rect 6270 6672 6276 6724
rect 6328 6672 6334 6724
rect 7101 6715 7159 6721
rect 7101 6681 7113 6715
rect 7147 6712 7159 6715
rect 7147 6684 7604 6712
rect 7147 6681 7159 6684
rect 7101 6675 7159 6681
rect 7576 6656 7604 6684
rect 7742 6672 7748 6724
rect 7800 6672 7806 6724
rect 10410 6672 10416 6724
rect 10468 6712 10474 6724
rect 10505 6715 10563 6721
rect 10505 6712 10517 6715
rect 10468 6684 10517 6712
rect 10468 6672 10474 6684
rect 10505 6681 10517 6684
rect 10551 6681 10563 6715
rect 10505 6675 10563 6681
rect 11330 6672 11336 6724
rect 11388 6712 11394 6724
rect 11425 6715 11483 6721
rect 11425 6712 11437 6715
rect 11388 6684 11437 6712
rect 11388 6672 11394 6684
rect 11425 6681 11437 6684
rect 11471 6712 11483 6715
rect 11514 6712 11520 6724
rect 11471 6684 11520 6712
rect 11471 6681 11483 6684
rect 11425 6675 11483 6681
rect 11514 6672 11520 6684
rect 11572 6672 11578 6724
rect 11701 6715 11759 6721
rect 11701 6681 11713 6715
rect 11747 6712 11759 6715
rect 12176 6712 12204 6879
rect 13906 6876 13912 6928
rect 13964 6876 13970 6928
rect 14108 6916 14136 6956
rect 14458 6944 14464 6996
rect 14516 6944 14522 6996
rect 16758 6944 16764 6996
rect 16816 6944 16822 6996
rect 17586 6984 17592 6996
rect 16868 6956 17592 6984
rect 14108 6888 14596 6916
rect 13924 6848 13952 6876
rect 14108 6860 14136 6888
rect 13740 6820 13952 6848
rect 13740 6789 13768 6820
rect 14090 6808 14096 6860
rect 14148 6808 14154 6860
rect 14568 6857 14596 6888
rect 14553 6851 14611 6857
rect 14200 6820 14504 6848
rect 13725 6783 13783 6789
rect 13725 6749 13737 6783
rect 13771 6749 13783 6783
rect 13725 6743 13783 6749
rect 13906 6740 13912 6792
rect 13964 6780 13970 6792
rect 14200 6780 14228 6820
rect 13964 6752 14228 6780
rect 14277 6783 14335 6789
rect 13964 6740 13970 6752
rect 14277 6749 14289 6783
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 11747 6684 12204 6712
rect 13817 6715 13875 6721
rect 11747 6681 11759 6684
rect 11701 6675 11759 6681
rect 13817 6681 13829 6715
rect 13863 6712 13875 6715
rect 14292 6712 14320 6743
rect 13863 6684 14320 6712
rect 14476 6712 14504 6820
rect 14553 6817 14565 6851
rect 14599 6848 14611 6851
rect 15470 6848 15476 6860
rect 14599 6820 15476 6848
rect 14599 6817 14611 6820
rect 14553 6811 14611 6817
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 16776 6848 16804 6944
rect 16868 6928 16896 6956
rect 17586 6944 17592 6956
rect 17644 6944 17650 6996
rect 20796 6987 20854 6993
rect 20796 6953 20808 6987
rect 20842 6984 20854 6987
rect 22002 6984 22008 6996
rect 20842 6956 22008 6984
rect 20842 6953 20854 6956
rect 20796 6947 20854 6953
rect 22002 6944 22008 6956
rect 22060 6944 22066 6996
rect 22278 6944 22284 6996
rect 22336 6944 22342 6996
rect 22728 6987 22786 6993
rect 22728 6953 22740 6987
rect 22774 6984 22786 6987
rect 24394 6984 24400 6996
rect 22774 6956 24400 6984
rect 22774 6953 22786 6956
rect 22728 6947 22786 6953
rect 24394 6944 24400 6956
rect 24452 6944 24458 6996
rect 16850 6876 16856 6928
rect 16908 6876 16914 6928
rect 16942 6876 16948 6928
rect 17000 6916 17006 6928
rect 17494 6916 17500 6928
rect 17000 6888 17500 6916
rect 17000 6876 17006 6888
rect 17494 6876 17500 6888
rect 17552 6916 17558 6928
rect 17552 6888 18000 6916
rect 17552 6876 17558 6888
rect 16776 6820 17908 6848
rect 17037 6783 17095 6789
rect 17037 6749 17049 6783
rect 17083 6749 17095 6783
rect 17037 6743 17095 6749
rect 14734 6712 14740 6724
rect 14476 6684 14740 6712
rect 13863 6681 13875 6684
rect 13817 6675 13875 6681
rect 14734 6672 14740 6684
rect 14792 6672 14798 6724
rect 17052 6712 17080 6743
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 17313 6783 17371 6789
rect 17313 6780 17325 6783
rect 17276 6752 17325 6780
rect 17276 6740 17282 6752
rect 17313 6749 17325 6752
rect 17359 6749 17371 6783
rect 17313 6743 17371 6749
rect 17402 6740 17408 6792
rect 17460 6740 17466 6792
rect 17880 6789 17908 6820
rect 17865 6783 17923 6789
rect 17865 6749 17877 6783
rect 17911 6749 17923 6783
rect 17972 6780 18000 6888
rect 24026 6876 24032 6928
rect 24084 6876 24090 6928
rect 24118 6876 24124 6928
rect 24176 6916 24182 6928
rect 24213 6919 24271 6925
rect 24213 6916 24225 6919
rect 24176 6888 24225 6916
rect 24176 6876 24182 6888
rect 24213 6885 24225 6888
rect 24259 6885 24271 6919
rect 24213 6879 24271 6885
rect 20070 6808 20076 6860
rect 20128 6848 20134 6860
rect 20533 6851 20591 6857
rect 20533 6848 20545 6851
rect 20128 6820 20545 6848
rect 20128 6808 20134 6820
rect 20533 6817 20545 6820
rect 20579 6848 20591 6851
rect 22465 6851 22523 6857
rect 22465 6848 22477 6851
rect 20579 6820 22477 6848
rect 20579 6817 20591 6820
rect 20533 6811 20591 6817
rect 22465 6817 22477 6820
rect 22511 6848 22523 6851
rect 22738 6848 22744 6860
rect 22511 6820 22744 6848
rect 22511 6817 22523 6820
rect 22465 6811 22523 6817
rect 22738 6808 22744 6820
rect 22796 6808 22802 6860
rect 22830 6808 22836 6860
rect 22888 6848 22894 6860
rect 24044 6848 24072 6876
rect 24489 6851 24547 6857
rect 24489 6848 24501 6851
rect 22888 6820 23980 6848
rect 24044 6820 24501 6848
rect 22888 6808 22894 6820
rect 18049 6783 18107 6789
rect 18049 6780 18061 6783
rect 17972 6752 18061 6780
rect 17865 6743 17923 6749
rect 18049 6749 18061 6752
rect 18095 6749 18107 6783
rect 23952 6780 23980 6820
rect 24489 6817 24501 6820
rect 24535 6817 24547 6851
rect 24489 6811 24547 6817
rect 24302 6780 24308 6792
rect 23952 6752 24308 6780
rect 18049 6743 18107 6749
rect 24302 6740 24308 6752
rect 24360 6780 24366 6792
rect 24397 6783 24455 6789
rect 24397 6780 24409 6783
rect 24360 6752 24409 6780
rect 24360 6740 24366 6752
rect 24397 6749 24409 6752
rect 24443 6749 24455 6783
rect 24397 6743 24455 6749
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6780 24639 6783
rect 24762 6780 24768 6792
rect 24627 6752 24768 6780
rect 24627 6749 24639 6752
rect 24581 6743 24639 6749
rect 24762 6740 24768 6752
rect 24820 6740 24826 6792
rect 17420 6712 17448 6740
rect 17052 6684 17448 6712
rect 17586 6672 17592 6724
rect 17644 6672 17650 6724
rect 17696 6684 18092 6712
rect 5905 6647 5963 6653
rect 5905 6644 5917 6647
rect 5276 6616 5917 6644
rect 5905 6613 5917 6616
rect 5951 6613 5963 6647
rect 5905 6607 5963 6613
rect 6546 6604 6552 6656
rect 6604 6604 6610 6656
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 7377 6647 7435 6653
rect 7377 6644 7389 6647
rect 6972 6616 7389 6644
rect 6972 6604 6978 6616
rect 7377 6613 7389 6616
rect 7423 6613 7435 6647
rect 7377 6607 7435 6613
rect 7558 6604 7564 6656
rect 7616 6604 7622 6656
rect 7760 6644 7788 6672
rect 10778 6644 10784 6656
rect 7760 6616 10784 6644
rect 10778 6604 10784 6616
rect 10836 6604 10842 6656
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 11793 6647 11851 6653
rect 11793 6644 11805 6647
rect 11204 6616 11805 6644
rect 11204 6604 11210 6616
rect 11793 6613 11805 6616
rect 11839 6644 11851 6647
rect 12158 6644 12164 6656
rect 11839 6616 12164 6644
rect 11839 6613 11851 6616
rect 11793 6607 11851 6613
rect 12158 6604 12164 6616
rect 12216 6604 12222 6656
rect 14090 6604 14096 6656
rect 14148 6604 14154 6656
rect 16853 6647 16911 6653
rect 16853 6613 16865 6647
rect 16899 6644 16911 6647
rect 17126 6644 17132 6656
rect 16899 6616 17132 6644
rect 16899 6613 16911 6616
rect 16853 6607 16911 6613
rect 17126 6604 17132 6616
rect 17184 6604 17190 6656
rect 17221 6647 17279 6653
rect 17221 6613 17233 6647
rect 17267 6644 17279 6647
rect 17696 6644 17724 6684
rect 18064 6656 18092 6684
rect 20806 6672 20812 6724
rect 20864 6712 20870 6724
rect 20864 6684 21298 6712
rect 23124 6684 23230 6712
rect 20864 6672 20870 6684
rect 17267 6616 17724 6644
rect 17267 6613 17279 6616
rect 17221 6607 17279 6613
rect 17770 6604 17776 6656
rect 17828 6604 17834 6656
rect 17954 6604 17960 6656
rect 18012 6604 18018 6656
rect 18046 6604 18052 6656
rect 18104 6604 18110 6656
rect 21192 6644 21220 6684
rect 23124 6644 23152 6684
rect 26510 6644 26516 6656
rect 21192 6616 26516 6644
rect 26510 6604 26516 6616
rect 26568 6604 26574 6656
rect 1104 6554 29595 6576
rect 1104 6502 8032 6554
rect 8084 6502 8096 6554
rect 8148 6502 8160 6554
rect 8212 6502 8224 6554
rect 8276 6502 8288 6554
rect 8340 6502 15115 6554
rect 15167 6502 15179 6554
rect 15231 6502 15243 6554
rect 15295 6502 15307 6554
rect 15359 6502 15371 6554
rect 15423 6502 22198 6554
rect 22250 6502 22262 6554
rect 22314 6502 22326 6554
rect 22378 6502 22390 6554
rect 22442 6502 22454 6554
rect 22506 6502 29281 6554
rect 29333 6502 29345 6554
rect 29397 6502 29409 6554
rect 29461 6502 29473 6554
rect 29525 6502 29537 6554
rect 29589 6502 29595 6554
rect 1104 6480 29595 6502
rect 5074 6440 5080 6452
rect 4172 6412 5080 6440
rect 4172 6381 4200 6412
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 5629 6443 5687 6449
rect 5629 6409 5641 6443
rect 5675 6440 5687 6443
rect 5902 6440 5908 6452
rect 5675 6412 5908 6440
rect 5675 6409 5687 6412
rect 5629 6403 5687 6409
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 7009 6443 7067 6449
rect 7009 6440 7021 6443
rect 6328 6412 7021 6440
rect 6328 6400 6334 6412
rect 7009 6409 7021 6412
rect 7055 6409 7067 6443
rect 7009 6403 7067 6409
rect 7466 6400 7472 6452
rect 7524 6440 7530 6452
rect 8757 6443 8815 6449
rect 8757 6440 8769 6443
rect 7524 6412 8769 6440
rect 7524 6400 7530 6412
rect 8757 6409 8769 6412
rect 8803 6409 8815 6443
rect 8757 6403 8815 6409
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 10873 6443 10931 6449
rect 10873 6440 10885 6443
rect 10284 6412 10885 6440
rect 10284 6400 10290 6412
rect 10873 6409 10885 6412
rect 10919 6409 10931 6443
rect 10873 6403 10931 6409
rect 11057 6443 11115 6449
rect 11057 6409 11069 6443
rect 11103 6440 11115 6443
rect 11422 6440 11428 6452
rect 11103 6412 11428 6440
rect 11103 6409 11115 6412
rect 11057 6403 11115 6409
rect 11422 6400 11428 6412
rect 11480 6400 11486 6452
rect 11698 6400 11704 6452
rect 11756 6400 11762 6452
rect 11790 6400 11796 6452
rect 11848 6400 11854 6452
rect 14090 6440 14096 6452
rect 13740 6412 14096 6440
rect 4157 6375 4215 6381
rect 4157 6341 4169 6375
rect 4203 6341 4215 6375
rect 4157 6335 4215 6341
rect 6822 6332 6828 6384
rect 6880 6372 6886 6384
rect 8021 6375 8079 6381
rect 8021 6372 8033 6375
rect 6880 6344 8033 6372
rect 6880 6332 6886 6344
rect 8021 6341 8033 6344
rect 8067 6341 8079 6375
rect 8021 6335 8079 6341
rect 10045 6375 10103 6381
rect 10045 6341 10057 6375
rect 10091 6372 10103 6375
rect 10502 6372 10508 6384
rect 10091 6344 10508 6372
rect 10091 6341 10103 6344
rect 10045 6335 10103 6341
rect 10502 6332 10508 6344
rect 10560 6372 10566 6384
rect 11716 6372 11744 6400
rect 10560 6344 11744 6372
rect 10560 6332 10566 6344
rect 2682 6264 2688 6316
rect 2740 6304 2746 6316
rect 3881 6307 3939 6313
rect 3881 6304 3893 6307
rect 2740 6276 3893 6304
rect 2740 6264 2746 6276
rect 3881 6273 3893 6276
rect 3927 6273 3939 6307
rect 3881 6267 3939 6273
rect 3786 6196 3792 6248
rect 3844 6236 3850 6248
rect 5276 6236 5304 6290
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 6236 6276 6500 6304
rect 6236 6264 6242 6276
rect 5350 6236 5356 6248
rect 3844 6208 5356 6236
rect 3844 6196 3850 6208
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 5718 6196 5724 6248
rect 5776 6236 5782 6248
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 5776 6208 6377 6236
rect 5776 6196 5782 6208
rect 6365 6205 6377 6208
rect 6411 6205 6423 6239
rect 6472 6236 6500 6276
rect 7190 6264 7196 6316
rect 7248 6304 7254 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7248 6276 7389 6304
rect 7248 6264 7254 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 7926 6264 7932 6316
rect 7984 6304 7990 6316
rect 8113 6307 8171 6313
rect 8113 6304 8125 6307
rect 7984 6276 8125 6304
rect 7984 6264 7990 6276
rect 8113 6273 8125 6276
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 9950 6264 9956 6316
rect 10008 6264 10014 6316
rect 10134 6264 10140 6316
rect 10192 6304 10198 6316
rect 10229 6307 10287 6313
rect 10229 6304 10241 6307
rect 10192 6276 10241 6304
rect 10192 6264 10198 6276
rect 10229 6273 10241 6276
rect 10275 6304 10287 6307
rect 10275 6276 10548 6304
rect 10275 6273 10287 6276
rect 10229 6267 10287 6273
rect 10410 6236 10416 6248
rect 6472 6208 10416 6236
rect 6365 6199 6423 6205
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 7374 6128 7380 6180
rect 7432 6168 7438 6180
rect 7834 6168 7840 6180
rect 7432 6140 7840 6168
rect 7432 6128 7438 6140
rect 7834 6128 7840 6140
rect 7892 6168 7898 6180
rect 10520 6168 10548 6276
rect 10594 6264 10600 6316
rect 10652 6264 10658 6316
rect 10962 6264 10968 6316
rect 11020 6264 11026 6316
rect 11146 6264 11152 6316
rect 11204 6264 11210 6316
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6304 11575 6307
rect 11808 6304 11836 6400
rect 13740 6381 13768 6412
rect 14090 6400 14096 6412
rect 14148 6400 14154 6452
rect 16574 6400 16580 6452
rect 16632 6440 16638 6452
rect 17129 6443 17187 6449
rect 17129 6440 17141 6443
rect 16632 6412 17141 6440
rect 16632 6400 16638 6412
rect 17129 6409 17141 6412
rect 17175 6440 17187 6443
rect 17770 6440 17776 6452
rect 17175 6412 17776 6440
rect 17175 6409 17187 6412
rect 17129 6403 17187 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 17954 6400 17960 6452
rect 18012 6400 18018 6452
rect 20070 6400 20076 6452
rect 20128 6400 20134 6452
rect 20441 6443 20499 6449
rect 20441 6409 20453 6443
rect 20487 6440 20499 6443
rect 20530 6440 20536 6452
rect 20487 6412 20536 6440
rect 20487 6409 20499 6412
rect 20441 6403 20499 6409
rect 20530 6400 20536 6412
rect 20588 6400 20594 6452
rect 20625 6443 20683 6449
rect 20625 6409 20637 6443
rect 20671 6440 20683 6443
rect 28718 6440 28724 6452
rect 20671 6412 28724 6440
rect 20671 6409 20683 6412
rect 20625 6403 20683 6409
rect 28718 6400 28724 6412
rect 28776 6400 28782 6452
rect 13725 6375 13783 6381
rect 13725 6341 13737 6375
rect 13771 6341 13783 6375
rect 13725 6335 13783 6341
rect 14182 6332 14188 6384
rect 14240 6332 14246 6384
rect 15470 6332 15476 6384
rect 15528 6332 15534 6384
rect 16850 6332 16856 6384
rect 16908 6372 16914 6384
rect 16945 6375 17003 6381
rect 16945 6372 16957 6375
rect 16908 6344 16957 6372
rect 16908 6332 16914 6344
rect 16945 6341 16957 6344
rect 16991 6372 17003 6375
rect 17862 6372 17868 6384
rect 16991 6344 17868 6372
rect 16991 6341 17003 6344
rect 16945 6335 17003 6341
rect 17862 6332 17868 6344
rect 17920 6332 17926 6384
rect 11563 6276 11836 6304
rect 17221 6307 17279 6313
rect 11563 6273 11575 6276
rect 11517 6267 11575 6273
rect 17221 6273 17233 6307
rect 17267 6304 17279 6307
rect 17972 6304 18000 6400
rect 20993 6375 21051 6381
rect 20272 6344 20852 6372
rect 20272 6316 20300 6344
rect 17267 6276 18000 6304
rect 17267 6273 17279 6276
rect 17221 6267 17279 6273
rect 20254 6264 20260 6316
rect 20312 6264 20318 6316
rect 20824 6313 20852 6344
rect 20993 6341 21005 6375
rect 21039 6372 21051 6375
rect 21039 6344 21220 6372
rect 21039 6341 21051 6344
rect 20993 6335 21051 6341
rect 20533 6307 20591 6313
rect 20533 6273 20545 6307
rect 20579 6273 20591 6307
rect 20533 6267 20591 6273
rect 20809 6307 20867 6313
rect 20809 6273 20821 6307
rect 20855 6273 20867 6307
rect 20809 6267 20867 6273
rect 21085 6307 21143 6313
rect 21085 6273 21097 6307
rect 21131 6273 21143 6307
rect 21085 6267 21143 6273
rect 10714 6239 10772 6245
rect 10714 6205 10726 6239
rect 10760 6236 10772 6239
rect 11164 6236 11192 6264
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 10760 6208 11192 6236
rect 11256 6208 11713 6236
rect 10760 6205 10772 6208
rect 10714 6199 10772 6205
rect 11146 6168 11152 6180
rect 7892 6140 10364 6168
rect 10520 6140 11152 6168
rect 7892 6128 7898 6140
rect 4614 6060 4620 6112
rect 4672 6100 4678 6112
rect 7558 6100 7564 6112
rect 4672 6072 7564 6100
rect 4672 6060 4678 6072
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 10336 6100 10364 6140
rect 11146 6128 11152 6140
rect 11204 6128 11210 6180
rect 11256 6100 11284 6208
rect 11701 6205 11713 6208
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 12434 6196 12440 6248
rect 12492 6236 12498 6248
rect 13446 6236 13452 6248
rect 12492 6208 13452 6236
rect 12492 6196 12498 6208
rect 13446 6196 13452 6208
rect 13504 6196 13510 6248
rect 20548 6236 20576 6267
rect 21100 6236 21128 6267
rect 20456 6208 21128 6236
rect 20456 6112 20484 6208
rect 20530 6128 20536 6180
rect 20588 6168 20594 6180
rect 21192 6168 21220 6344
rect 20588 6140 21220 6168
rect 20588 6128 20594 6140
rect 10336 6072 11284 6100
rect 16945 6103 17003 6109
rect 16945 6069 16957 6103
rect 16991 6100 17003 6103
rect 17586 6100 17592 6112
rect 16991 6072 17592 6100
rect 16991 6069 17003 6072
rect 16945 6063 17003 6069
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 20438 6060 20444 6112
rect 20496 6060 20502 6112
rect 1104 6010 29440 6032
rect 1104 5958 4491 6010
rect 4543 5958 4555 6010
rect 4607 5958 4619 6010
rect 4671 5958 4683 6010
rect 4735 5958 4747 6010
rect 4799 5958 11574 6010
rect 11626 5958 11638 6010
rect 11690 5958 11702 6010
rect 11754 5958 11766 6010
rect 11818 5958 11830 6010
rect 11882 5958 18657 6010
rect 18709 5958 18721 6010
rect 18773 5958 18785 6010
rect 18837 5958 18849 6010
rect 18901 5958 18913 6010
rect 18965 5958 25740 6010
rect 25792 5958 25804 6010
rect 25856 5958 25868 6010
rect 25920 5958 25932 6010
rect 25984 5958 25996 6010
rect 26048 5958 29440 6010
rect 1104 5936 29440 5958
rect 4236 5899 4294 5905
rect 4236 5865 4248 5899
rect 4282 5896 4294 5899
rect 6546 5896 6552 5908
rect 4282 5868 6552 5896
rect 4282 5865 4294 5868
rect 4236 5859 4294 5865
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 8021 5899 8079 5905
rect 8021 5896 8033 5899
rect 7248 5868 8033 5896
rect 7248 5856 7254 5868
rect 8021 5865 8033 5868
rect 8067 5865 8079 5899
rect 8021 5859 8079 5865
rect 9628 5856 9634 5908
rect 9686 5896 9692 5908
rect 10042 5896 10048 5908
rect 9686 5868 10048 5896
rect 9686 5856 9692 5868
rect 10042 5856 10048 5868
rect 10100 5896 10106 5908
rect 10781 5899 10839 5905
rect 10781 5896 10793 5899
rect 10100 5868 10793 5896
rect 10100 5856 10106 5868
rect 10781 5865 10793 5868
rect 10827 5865 10839 5899
rect 10781 5859 10839 5865
rect 11054 5856 11060 5908
rect 11112 5856 11118 5908
rect 11146 5856 11152 5908
rect 11204 5896 11210 5908
rect 11330 5896 11336 5908
rect 11204 5868 11336 5896
rect 11204 5856 11210 5868
rect 11330 5856 11336 5868
rect 11388 5856 11394 5908
rect 16942 5856 16948 5908
rect 17000 5896 17006 5908
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 17000 5868 17693 5896
rect 17000 5856 17006 5868
rect 17681 5865 17693 5868
rect 17727 5865 17739 5899
rect 17681 5859 17739 5865
rect 5718 5788 5724 5840
rect 5776 5788 5782 5840
rect 7558 5788 7564 5840
rect 7616 5828 7622 5840
rect 13998 5828 14004 5840
rect 7616 5800 14004 5828
rect 7616 5788 7622 5800
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 17218 5788 17224 5840
rect 17276 5828 17282 5840
rect 17865 5831 17923 5837
rect 17865 5828 17877 5831
rect 17276 5800 17877 5828
rect 17276 5788 17282 5800
rect 17865 5797 17877 5800
rect 17911 5797 17923 5831
rect 17865 5791 17923 5797
rect 2682 5720 2688 5772
rect 2740 5720 2746 5772
rect 6270 5760 6276 5772
rect 3988 5732 6276 5760
rect 2700 5692 2728 5720
rect 3988 5701 4016 5732
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 6549 5763 6607 5769
rect 6549 5729 6561 5763
rect 6595 5760 6607 5763
rect 6914 5760 6920 5772
rect 6595 5732 6920 5760
rect 6595 5729 6607 5732
rect 6549 5723 6607 5729
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 10873 5763 10931 5769
rect 10873 5760 10885 5763
rect 9692 5732 10885 5760
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 2700 5664 3985 5692
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 5350 5652 5356 5704
rect 5408 5652 5414 5704
rect 9401 5695 9459 5701
rect 9401 5661 9413 5695
rect 9447 5692 9459 5695
rect 9490 5692 9496 5704
rect 9447 5664 9496 5692
rect 9447 5661 9459 5664
rect 9401 5655 9459 5661
rect 9490 5652 9496 5664
rect 9548 5652 9554 5704
rect 9692 5701 9720 5732
rect 10873 5729 10885 5732
rect 10919 5760 10931 5763
rect 11422 5760 11428 5772
rect 10919 5732 11428 5760
rect 10919 5729 10931 5732
rect 10873 5723 10931 5729
rect 11422 5720 11428 5732
rect 11480 5760 11486 5772
rect 11480 5732 11652 5760
rect 11480 5720 11486 5732
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5661 9735 5695
rect 9677 5655 9735 5661
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 10045 5695 10103 5701
rect 10045 5661 10057 5695
rect 10091 5661 10103 5695
rect 10045 5655 10103 5661
rect 5368 5556 5396 5652
rect 7006 5624 7012 5636
rect 5552 5596 7012 5624
rect 5552 5556 5580 5596
rect 7006 5584 7012 5596
rect 7064 5584 7070 5636
rect 9585 5627 9643 5633
rect 9585 5593 9597 5627
rect 9631 5624 9643 5627
rect 9631 5596 9904 5624
rect 9631 5593 9643 5596
rect 9585 5587 9643 5593
rect 9876 5568 9904 5596
rect 5368 5528 5580 5556
rect 9217 5559 9275 5565
rect 9217 5525 9229 5559
rect 9263 5556 9275 5559
rect 9306 5556 9312 5568
rect 9263 5528 9312 5556
rect 9263 5525 9275 5528
rect 9217 5519 9275 5525
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 9766 5516 9772 5568
rect 9824 5516 9830 5568
rect 9858 5516 9864 5568
rect 9916 5516 9922 5568
rect 9968 5556 9996 5655
rect 10060 5624 10088 5655
rect 10134 5652 10140 5704
rect 10192 5652 10198 5704
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5692 10287 5695
rect 10413 5695 10471 5701
rect 10413 5692 10425 5695
rect 10275 5664 10425 5692
rect 10275 5661 10287 5664
rect 10229 5655 10287 5661
rect 10413 5661 10425 5664
rect 10459 5661 10471 5695
rect 10413 5655 10471 5661
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5692 10655 5695
rect 10965 5695 11023 5701
rect 10965 5692 10977 5695
rect 10643 5664 10977 5692
rect 10643 5661 10655 5664
rect 10597 5655 10655 5661
rect 10888 5636 10916 5664
rect 10965 5661 10977 5664
rect 11011 5661 11023 5695
rect 10965 5655 11023 5661
rect 11146 5652 11152 5704
rect 11204 5652 11210 5704
rect 11238 5652 11244 5704
rect 11296 5652 11302 5704
rect 11624 5701 11652 5732
rect 17034 5720 17040 5772
rect 17092 5760 17098 5772
rect 17402 5760 17408 5772
rect 17092 5732 17408 5760
rect 17092 5720 17098 5732
rect 17402 5720 17408 5732
rect 17460 5760 17466 5772
rect 17460 5732 18276 5760
rect 17460 5720 17466 5732
rect 17604 5701 17632 5732
rect 18248 5701 18276 5732
rect 11517 5695 11575 5701
rect 11517 5692 11529 5695
rect 11348 5664 11529 5692
rect 10318 5624 10324 5636
rect 10060 5596 10324 5624
rect 10318 5584 10324 5596
rect 10376 5584 10382 5636
rect 10870 5584 10876 5636
rect 10928 5584 10934 5636
rect 11256 5556 11284 5652
rect 11348 5636 11376 5664
rect 11517 5661 11529 5664
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 11609 5695 11667 5701
rect 11609 5661 11621 5695
rect 11655 5661 11667 5695
rect 11609 5655 11667 5661
rect 17589 5695 17647 5701
rect 17589 5661 17601 5695
rect 17635 5661 17647 5695
rect 18141 5695 18199 5701
rect 18141 5692 18153 5695
rect 17589 5655 17647 5661
rect 17972 5664 18153 5692
rect 11330 5584 11336 5636
rect 11388 5584 11394 5636
rect 11422 5584 11428 5636
rect 11480 5584 11486 5636
rect 17405 5627 17463 5633
rect 17405 5593 17417 5627
rect 17451 5624 17463 5627
rect 17494 5624 17500 5636
rect 17451 5596 17500 5624
rect 17451 5593 17463 5596
rect 17405 5587 17463 5593
rect 17494 5584 17500 5596
rect 17552 5584 17558 5636
rect 17865 5627 17923 5633
rect 17865 5593 17877 5627
rect 17911 5593 17923 5627
rect 17865 5587 17923 5593
rect 9968 5528 11284 5556
rect 11790 5516 11796 5568
rect 11848 5516 11854 5568
rect 16298 5516 16304 5568
rect 16356 5556 16362 5568
rect 17512 5556 17540 5584
rect 17770 5556 17776 5568
rect 16356 5528 17776 5556
rect 16356 5516 16362 5528
rect 17770 5516 17776 5528
rect 17828 5556 17834 5568
rect 17880 5556 17908 5587
rect 17972 5568 18000 5664
rect 18141 5661 18153 5664
rect 18187 5661 18199 5695
rect 18141 5655 18199 5661
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5661 18291 5695
rect 18233 5655 18291 5661
rect 18248 5624 18276 5655
rect 18322 5652 18328 5704
rect 18380 5692 18386 5704
rect 18417 5695 18475 5701
rect 18417 5692 18429 5695
rect 18380 5664 18429 5692
rect 18380 5652 18386 5664
rect 18417 5661 18429 5664
rect 18463 5661 18475 5695
rect 18417 5655 18475 5661
rect 18248 5596 18552 5624
rect 18524 5568 18552 5596
rect 17828 5528 17908 5556
rect 17828 5516 17834 5528
rect 17954 5516 17960 5568
rect 18012 5516 18018 5568
rect 18049 5559 18107 5565
rect 18049 5525 18061 5559
rect 18095 5556 18107 5559
rect 18230 5556 18236 5568
rect 18095 5528 18236 5556
rect 18095 5525 18107 5528
rect 18049 5519 18107 5525
rect 18230 5516 18236 5528
rect 18288 5556 18294 5568
rect 18325 5559 18383 5565
rect 18325 5556 18337 5559
rect 18288 5528 18337 5556
rect 18288 5516 18294 5528
rect 18325 5525 18337 5528
rect 18371 5525 18383 5559
rect 18325 5519 18383 5525
rect 18506 5516 18512 5568
rect 18564 5516 18570 5568
rect 1104 5466 29595 5488
rect 1104 5414 8032 5466
rect 8084 5414 8096 5466
rect 8148 5414 8160 5466
rect 8212 5414 8224 5466
rect 8276 5414 8288 5466
rect 8340 5414 15115 5466
rect 15167 5414 15179 5466
rect 15231 5414 15243 5466
rect 15295 5414 15307 5466
rect 15359 5414 15371 5466
rect 15423 5414 22198 5466
rect 22250 5414 22262 5466
rect 22314 5414 22326 5466
rect 22378 5414 22390 5466
rect 22442 5414 22454 5466
rect 22506 5414 29281 5466
rect 29333 5414 29345 5466
rect 29397 5414 29409 5466
rect 29461 5414 29473 5466
rect 29525 5414 29537 5466
rect 29589 5414 29595 5466
rect 1104 5392 29595 5414
rect 7282 5352 7288 5364
rect 6656 5324 7288 5352
rect 6656 5293 6684 5324
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 7926 5312 7932 5364
rect 7984 5352 7990 5364
rect 8113 5355 8171 5361
rect 8113 5352 8125 5355
rect 7984 5324 8125 5352
rect 7984 5312 7990 5324
rect 8113 5321 8125 5324
rect 8159 5321 8171 5355
rect 8938 5352 8944 5364
rect 8113 5315 8171 5321
rect 8496 5324 8944 5352
rect 6641 5287 6699 5293
rect 6641 5253 6653 5287
rect 6687 5253 6699 5287
rect 6641 5247 6699 5253
rect 7098 5244 7104 5296
rect 7156 5244 7162 5296
rect 6270 5176 6276 5228
rect 6328 5216 6334 5228
rect 8496 5225 8524 5324
rect 8938 5312 8944 5324
rect 8996 5352 9002 5364
rect 12342 5352 12348 5364
rect 8996 5324 12348 5352
rect 8996 5312 9002 5324
rect 11057 5287 11115 5293
rect 11057 5284 11069 5287
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 6328 5188 6377 5216
rect 6328 5176 6334 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 8481 5219 8539 5225
rect 8481 5185 8493 5219
rect 8527 5185 8539 5219
rect 8481 5179 8539 5185
rect 9766 5176 9772 5228
rect 9824 5176 9830 5228
rect 8849 5151 8907 5157
rect 8849 5117 8861 5151
rect 8895 5148 8907 5151
rect 9784 5148 9812 5176
rect 8895 5120 9812 5148
rect 9876 5148 9904 5270
rect 9968 5256 11069 5284
rect 9968 5228 9996 5256
rect 11057 5253 11069 5256
rect 11103 5253 11115 5287
rect 11057 5247 11115 5253
rect 9950 5176 9956 5228
rect 10008 5176 10014 5228
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 10505 5219 10563 5225
rect 10505 5216 10517 5219
rect 10192 5188 10517 5216
rect 10192 5176 10198 5188
rect 10505 5185 10517 5188
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 10870 5176 10876 5228
rect 10928 5176 10934 5228
rect 11532 5225 11560 5324
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 12492 5324 13032 5352
rect 12492 5312 12498 5324
rect 13004 5284 13032 5324
rect 14550 5312 14556 5364
rect 14608 5312 14614 5364
rect 16879 5355 16937 5361
rect 16879 5321 16891 5355
rect 16925 5352 16937 5355
rect 17218 5352 17224 5364
rect 16925 5324 17224 5352
rect 16925 5321 16937 5324
rect 16879 5315 16937 5321
rect 17218 5312 17224 5324
rect 17276 5312 17282 5364
rect 17310 5312 17316 5364
rect 17368 5352 17374 5364
rect 17368 5324 19656 5352
rect 17368 5312 17374 5324
rect 13311 5287 13369 5293
rect 13311 5284 13323 5287
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 11848 5188 11897 5216
rect 11848 5176 11854 5188
rect 11885 5185 11897 5188
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 12728 5216 12756 5270
rect 13004 5256 13323 5284
rect 13311 5253 13323 5256
rect 13357 5253 13369 5287
rect 13311 5247 13369 5253
rect 14182 5216 14188 5228
rect 12728 5188 14188 5216
rect 9876 5120 9996 5148
rect 8895 5117 8907 5120
rect 8849 5111 8907 5117
rect 9968 5012 9996 5120
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10321 5151 10379 5157
rect 10321 5148 10333 5151
rect 10100 5120 10333 5148
rect 10100 5108 10106 5120
rect 10321 5117 10333 5120
rect 10367 5148 10379 5151
rect 10888 5148 10916 5176
rect 10367 5120 10916 5148
rect 10367 5117 10379 5120
rect 10321 5111 10379 5117
rect 11330 5108 11336 5160
rect 11388 5148 11394 5160
rect 12066 5148 12072 5160
rect 11388 5120 12072 5148
rect 11388 5108 11394 5120
rect 12066 5108 12072 5120
rect 12124 5148 12130 5160
rect 12434 5148 12440 5160
rect 12124 5120 12440 5148
rect 12124 5108 12130 5120
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 10318 5012 10324 5024
rect 9968 4984 10324 5012
rect 10318 4972 10324 4984
rect 10376 5012 10382 5024
rect 12728 5012 12756 5188
rect 14182 5176 14188 5188
rect 14240 5176 14246 5228
rect 14568 5216 14596 5312
rect 16669 5287 16727 5293
rect 16669 5253 16681 5287
rect 16715 5284 16727 5287
rect 16758 5284 16764 5296
rect 16715 5256 16764 5284
rect 16715 5253 16727 5256
rect 16669 5247 16727 5253
rect 16758 5244 16764 5256
rect 16816 5284 16822 5296
rect 17678 5284 17684 5296
rect 16816 5256 17684 5284
rect 16816 5244 16822 5256
rect 17034 5216 17040 5228
rect 14568 5188 17040 5216
rect 17034 5176 17040 5188
rect 17092 5176 17098 5228
rect 17129 5219 17187 5225
rect 17129 5185 17141 5219
rect 17175 5216 17187 5219
rect 17402 5216 17408 5228
rect 17175 5188 17408 5216
rect 17175 5185 17187 5188
rect 17129 5179 17187 5185
rect 16390 5108 16396 5160
rect 16448 5148 16454 5160
rect 17144 5148 17172 5179
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 17512 5225 17540 5256
rect 17678 5244 17684 5256
rect 17736 5284 17742 5296
rect 17736 5256 17816 5284
rect 17736 5244 17742 5256
rect 17788 5225 17816 5256
rect 17880 5256 19012 5284
rect 17880 5228 17908 5256
rect 17497 5219 17555 5225
rect 17497 5185 17509 5219
rect 17543 5185 17555 5219
rect 17497 5179 17555 5185
rect 17773 5219 17831 5225
rect 17773 5185 17785 5219
rect 17819 5185 17831 5219
rect 17773 5179 17831 5185
rect 17862 5176 17868 5228
rect 17920 5176 17926 5228
rect 17957 5219 18015 5225
rect 17957 5185 17969 5219
rect 18003 5185 18015 5219
rect 17957 5179 18015 5185
rect 16448 5120 17172 5148
rect 16448 5108 16454 5120
rect 17972 5080 18000 5179
rect 18230 5176 18236 5228
rect 18288 5176 18294 5228
rect 18322 5176 18328 5228
rect 18380 5176 18386 5228
rect 18506 5176 18512 5228
rect 18564 5176 18570 5228
rect 18984 5225 19012 5256
rect 19628 5225 19656 5324
rect 20254 5312 20260 5364
rect 20312 5352 20318 5364
rect 20349 5355 20407 5361
rect 20349 5352 20361 5355
rect 20312 5324 20361 5352
rect 20312 5312 20318 5324
rect 20349 5321 20361 5324
rect 20395 5321 20407 5355
rect 20349 5315 20407 5321
rect 28258 5312 28264 5364
rect 28316 5312 28322 5364
rect 18693 5219 18751 5225
rect 18693 5185 18705 5219
rect 18739 5185 18751 5219
rect 18693 5179 18751 5185
rect 18969 5219 19027 5225
rect 18969 5185 18981 5219
rect 19015 5185 19027 5219
rect 18969 5179 19027 5185
rect 19153 5219 19211 5225
rect 19153 5185 19165 5219
rect 19199 5185 19211 5219
rect 19153 5179 19211 5185
rect 19613 5219 19671 5225
rect 19613 5185 19625 5219
rect 19659 5185 19671 5219
rect 20257 5219 20315 5225
rect 20257 5216 20269 5219
rect 19613 5179 19671 5185
rect 20088 5188 20269 5216
rect 18340 5148 18368 5176
rect 18708 5148 18736 5179
rect 19168 5148 19196 5179
rect 18340 5120 19196 5148
rect 18046 5080 18052 5092
rect 17788 5052 18052 5080
rect 10376 4984 12756 5012
rect 10376 4972 10382 4984
rect 16850 4972 16856 5024
rect 16908 4972 16914 5024
rect 17034 4972 17040 5024
rect 17092 4972 17098 5024
rect 17126 4972 17132 5024
rect 17184 5012 17190 5024
rect 17497 5015 17555 5021
rect 17497 5012 17509 5015
rect 17184 4984 17509 5012
rect 17184 4972 17190 4984
rect 17497 4981 17509 4984
rect 17543 5012 17555 5015
rect 17788 5012 17816 5052
rect 18046 5040 18052 5052
rect 18104 5040 18110 5092
rect 18138 5040 18144 5092
rect 18196 5080 18202 5092
rect 18969 5083 19027 5089
rect 18969 5080 18981 5083
rect 18196 5052 18981 5080
rect 18196 5040 18202 5052
rect 18969 5049 18981 5052
rect 19015 5049 19027 5083
rect 19628 5080 19656 5179
rect 20088 5157 20116 5188
rect 20257 5185 20269 5188
rect 20303 5185 20315 5219
rect 20257 5179 20315 5185
rect 28074 5176 28080 5228
rect 28132 5176 28138 5228
rect 20073 5151 20131 5157
rect 20073 5117 20085 5151
rect 20119 5117 20131 5151
rect 20073 5111 20131 5117
rect 19628 5052 20760 5080
rect 18969 5043 19027 5049
rect 20732 5024 20760 5052
rect 17543 4984 17816 5012
rect 17543 4981 17555 4984
rect 17497 4975 17555 4981
rect 17862 4972 17868 5024
rect 17920 4972 17926 5024
rect 17954 4972 17960 5024
rect 18012 5012 18018 5024
rect 18877 5015 18935 5021
rect 18877 5012 18889 5015
rect 18012 4984 18889 5012
rect 18012 4972 18018 4984
rect 18877 4981 18889 4984
rect 18923 4981 18935 5015
rect 18877 4975 18935 4981
rect 19518 4972 19524 5024
rect 19576 5012 19582 5024
rect 19705 5015 19763 5021
rect 19705 5012 19717 5015
rect 19576 4984 19717 5012
rect 19576 4972 19582 4984
rect 19705 4981 19717 4984
rect 19751 4981 19763 5015
rect 19705 4975 19763 4981
rect 20714 4972 20720 5024
rect 20772 4972 20778 5024
rect 1104 4922 29440 4944
rect 1104 4870 4491 4922
rect 4543 4870 4555 4922
rect 4607 4870 4619 4922
rect 4671 4870 4683 4922
rect 4735 4870 4747 4922
rect 4799 4870 11574 4922
rect 11626 4870 11638 4922
rect 11690 4870 11702 4922
rect 11754 4870 11766 4922
rect 11818 4870 11830 4922
rect 11882 4870 18657 4922
rect 18709 4870 18721 4922
rect 18773 4870 18785 4922
rect 18837 4870 18849 4922
rect 18901 4870 18913 4922
rect 18965 4870 25740 4922
rect 25792 4870 25804 4922
rect 25856 4870 25868 4922
rect 25920 4870 25932 4922
rect 25984 4870 25996 4922
rect 26048 4870 29440 4922
rect 1104 4848 29440 4870
rect 10134 4768 10140 4820
rect 10192 4808 10198 4820
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 10192 4780 10701 4808
rect 10192 4768 10198 4780
rect 10689 4777 10701 4780
rect 10735 4777 10747 4811
rect 10689 4771 10747 4777
rect 11054 4768 11060 4820
rect 11112 4768 11118 4820
rect 11333 4811 11391 4817
rect 11333 4777 11345 4811
rect 11379 4808 11391 4811
rect 11422 4808 11428 4820
rect 11379 4780 11428 4808
rect 11379 4777 11391 4780
rect 11333 4771 11391 4777
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 16298 4808 16304 4820
rect 15948 4780 16304 4808
rect 8938 4632 8944 4684
rect 8996 4632 9002 4684
rect 9306 4632 9312 4684
rect 9364 4632 9370 4684
rect 10318 4632 10324 4684
rect 10376 4632 10382 4684
rect 11072 4672 11100 4768
rect 11149 4675 11207 4681
rect 11149 4672 11161 4675
rect 11072 4644 11161 4672
rect 11149 4641 11161 4644
rect 11195 4641 11207 4675
rect 13357 4675 13415 4681
rect 13357 4672 13369 4675
rect 11149 4635 11207 4641
rect 13004 4644 13369 4672
rect 10336 4522 10364 4632
rect 13004 4616 13032 4644
rect 13357 4641 13369 4644
rect 13403 4641 13415 4675
rect 13357 4635 13415 4641
rect 11057 4607 11115 4613
rect 11057 4573 11069 4607
rect 11103 4604 11115 4607
rect 11330 4604 11336 4616
rect 11103 4576 11336 4604
rect 11103 4573 11115 4576
rect 11057 4567 11115 4573
rect 11330 4564 11336 4576
rect 11388 4564 11394 4616
rect 12986 4564 12992 4616
rect 13044 4564 13050 4616
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4573 13139 4607
rect 13081 4567 13139 4573
rect 13096 4536 13124 4567
rect 13262 4564 13268 4616
rect 13320 4564 13326 4616
rect 15948 4613 15976 4780
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 16482 4768 16488 4820
rect 16540 4808 16546 4820
rect 16942 4808 16948 4820
rect 16540 4780 16948 4808
rect 16540 4768 16546 4780
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 17586 4768 17592 4820
rect 17644 4768 17650 4820
rect 17862 4768 17868 4820
rect 17920 4808 17926 4820
rect 17920 4780 18920 4808
rect 17920 4768 17926 4780
rect 16209 4743 16267 4749
rect 16209 4709 16221 4743
rect 16255 4740 16267 4743
rect 18785 4743 18843 4749
rect 18785 4740 18797 4743
rect 16255 4712 18797 4740
rect 16255 4709 16267 4712
rect 16209 4703 16267 4709
rect 18785 4709 18797 4712
rect 18831 4709 18843 4743
rect 18785 4703 18843 4709
rect 18892 4740 18920 4780
rect 19794 4768 19800 4820
rect 19852 4808 19858 4820
rect 19981 4811 20039 4817
rect 19981 4808 19993 4811
rect 19852 4780 19993 4808
rect 19852 4768 19858 4780
rect 19981 4777 19993 4780
rect 20027 4777 20039 4811
rect 19981 4771 20039 4777
rect 20441 4811 20499 4817
rect 20441 4777 20453 4811
rect 20487 4808 20499 4811
rect 28074 4808 28080 4820
rect 20487 4780 28080 4808
rect 20487 4777 20499 4780
rect 20441 4771 20499 4777
rect 28074 4768 28080 4780
rect 28132 4768 28138 4820
rect 19334 4740 19340 4752
rect 18892 4712 19340 4740
rect 16022 4632 16028 4684
rect 16080 4672 16086 4684
rect 16080 4644 16712 4672
rect 16080 4632 16086 4644
rect 15933 4607 15991 4613
rect 15933 4573 15945 4607
rect 15979 4573 15991 4607
rect 15933 4567 15991 4573
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4604 16175 4607
rect 16390 4604 16396 4616
rect 16163 4576 16396 4604
rect 16163 4573 16175 4576
rect 16117 4567 16175 4573
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 16482 4564 16488 4616
rect 16540 4564 16546 4616
rect 16574 4564 16580 4616
rect 16632 4564 16638 4616
rect 16684 4604 16712 4644
rect 17034 4632 17040 4684
rect 17092 4672 17098 4684
rect 18892 4681 18920 4712
rect 19334 4700 19340 4712
rect 19392 4740 19398 4752
rect 20530 4740 20536 4752
rect 19392 4712 20536 4740
rect 19392 4700 19398 4712
rect 20530 4700 20536 4712
rect 20588 4700 20594 4752
rect 17681 4675 17739 4681
rect 17681 4672 17693 4675
rect 17092 4644 17693 4672
rect 17092 4632 17098 4644
rect 17681 4641 17693 4644
rect 17727 4641 17739 4675
rect 18141 4675 18199 4681
rect 18141 4672 18153 4675
rect 17681 4635 17739 4641
rect 17788 4644 18153 4672
rect 16684 4576 17264 4604
rect 13998 4536 14004 4548
rect 13096 4508 14004 4536
rect 13998 4496 14004 4508
rect 14056 4496 14062 4548
rect 16206 4496 16212 4548
rect 16264 4496 16270 4548
rect 16298 4496 16304 4548
rect 16356 4536 16362 4548
rect 17236 4536 17264 4576
rect 17402 4564 17408 4616
rect 17460 4564 17466 4616
rect 17788 4604 17816 4644
rect 18141 4641 18153 4644
rect 18187 4641 18199 4675
rect 18141 4635 18199 4641
rect 18417 4675 18475 4681
rect 18417 4641 18429 4675
rect 18463 4672 18475 4675
rect 18877 4675 18935 4681
rect 18463 4644 18828 4672
rect 18463 4641 18475 4644
rect 18417 4635 18475 4641
rect 17512 4576 17816 4604
rect 17512 4536 17540 4576
rect 17862 4564 17868 4616
rect 17920 4604 17926 4616
rect 17957 4607 18015 4613
rect 17957 4604 17969 4607
rect 17920 4576 17969 4604
rect 17920 4564 17926 4576
rect 17957 4573 17969 4576
rect 18003 4573 18015 4607
rect 17957 4567 18015 4573
rect 18046 4564 18052 4616
rect 18104 4604 18110 4616
rect 18233 4607 18291 4613
rect 18233 4604 18245 4607
rect 18104 4576 18245 4604
rect 18104 4564 18110 4576
rect 18233 4573 18245 4576
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 18601 4607 18659 4613
rect 18601 4573 18613 4607
rect 18647 4573 18659 4607
rect 18601 4567 18659 4573
rect 16356 4508 17172 4536
rect 17236 4508 17540 4536
rect 16356 4496 16362 4508
rect 6454 4428 6460 4480
rect 6512 4468 6518 4480
rect 12897 4471 12955 4477
rect 12897 4468 12909 4471
rect 6512 4440 12909 4468
rect 6512 4428 6518 4440
rect 12897 4437 12909 4440
rect 12943 4437 12955 4471
rect 12897 4431 12955 4437
rect 16393 4471 16451 4477
rect 16393 4437 16405 4471
rect 16439 4468 16451 4471
rect 16850 4468 16856 4480
rect 16439 4440 16856 4468
rect 16439 4437 16451 4440
rect 16393 4431 16451 4437
rect 16850 4428 16856 4440
rect 16908 4468 16914 4480
rect 17144 4477 17172 4508
rect 17586 4496 17592 4548
rect 17644 4536 17650 4548
rect 17773 4539 17831 4545
rect 17773 4536 17785 4539
rect 17644 4508 17785 4536
rect 17644 4496 17650 4508
rect 17773 4505 17785 4508
rect 17819 4536 17831 4539
rect 18616 4536 18644 4567
rect 17819 4508 18644 4536
rect 18800 4536 18828 4644
rect 18877 4641 18889 4675
rect 18923 4641 18935 4675
rect 19518 4672 19524 4684
rect 18877 4635 18935 4641
rect 19168 4644 19524 4672
rect 19168 4536 19196 4644
rect 19518 4632 19524 4644
rect 19576 4632 19582 4684
rect 19613 4675 19671 4681
rect 19613 4641 19625 4675
rect 19659 4672 19671 4675
rect 19659 4644 20208 4672
rect 19659 4641 19671 4644
rect 19613 4635 19671 4641
rect 20180 4616 20208 4644
rect 19242 4564 19248 4616
rect 19300 4564 19306 4616
rect 19426 4564 19432 4616
rect 19484 4564 19490 4616
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4604 19763 4607
rect 19794 4604 19800 4616
rect 19751 4576 19800 4604
rect 19751 4573 19763 4576
rect 19705 4567 19763 4573
rect 19794 4564 19800 4576
rect 19852 4564 19858 4616
rect 19889 4607 19947 4613
rect 19889 4573 19901 4607
rect 19935 4573 19947 4607
rect 19889 4567 19947 4573
rect 18800 4508 19196 4536
rect 19260 4536 19288 4564
rect 19904 4536 19932 4567
rect 20162 4564 20168 4616
rect 20220 4564 20226 4616
rect 20438 4564 20444 4616
rect 20496 4604 20502 4616
rect 20533 4607 20591 4613
rect 20533 4604 20545 4607
rect 20496 4576 20545 4604
rect 20496 4564 20502 4576
rect 20533 4573 20545 4576
rect 20579 4573 20591 4607
rect 20533 4567 20591 4573
rect 20714 4564 20720 4616
rect 20772 4564 20778 4616
rect 20625 4539 20683 4545
rect 20625 4536 20637 4539
rect 19260 4508 20637 4536
rect 17819 4505 17831 4508
rect 17773 4499 17831 4505
rect 20625 4505 20637 4508
rect 20671 4505 20683 4539
rect 20625 4499 20683 4505
rect 16945 4471 17003 4477
rect 16945 4468 16957 4471
rect 16908 4440 16957 4468
rect 16908 4428 16914 4440
rect 16945 4437 16957 4440
rect 16991 4437 17003 4471
rect 16945 4431 17003 4437
rect 17129 4471 17187 4477
rect 17129 4437 17141 4471
rect 17175 4437 17187 4471
rect 17129 4431 17187 4437
rect 17218 4428 17224 4480
rect 17276 4428 17282 4480
rect 17678 4428 17684 4480
rect 17736 4468 17742 4480
rect 17862 4468 17868 4480
rect 17736 4440 17868 4468
rect 17736 4428 17742 4440
rect 17862 4428 17868 4440
rect 17920 4468 17926 4480
rect 18230 4468 18236 4480
rect 17920 4440 18236 4468
rect 17920 4428 17926 4440
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 18322 4428 18328 4480
rect 18380 4468 18386 4480
rect 19245 4471 19303 4477
rect 19245 4468 19257 4471
rect 18380 4440 19257 4468
rect 18380 4428 18386 4440
rect 19245 4437 19257 4440
rect 19291 4437 19303 4471
rect 19245 4431 19303 4437
rect 1104 4378 29595 4400
rect 1104 4326 8032 4378
rect 8084 4326 8096 4378
rect 8148 4326 8160 4378
rect 8212 4326 8224 4378
rect 8276 4326 8288 4378
rect 8340 4326 15115 4378
rect 15167 4326 15179 4378
rect 15231 4326 15243 4378
rect 15295 4326 15307 4378
rect 15359 4326 15371 4378
rect 15423 4326 22198 4378
rect 22250 4326 22262 4378
rect 22314 4326 22326 4378
rect 22378 4326 22390 4378
rect 22442 4326 22454 4378
rect 22506 4326 29281 4378
rect 29333 4326 29345 4378
rect 29397 4326 29409 4378
rect 29461 4326 29473 4378
rect 29525 4326 29537 4378
rect 29589 4326 29595 4378
rect 1104 4304 29595 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 2464 4236 2774 4264
rect 2464 4224 2470 4236
rect 2746 4196 2774 4236
rect 13170 4224 13176 4276
rect 13228 4224 13234 4276
rect 13909 4267 13967 4273
rect 13909 4233 13921 4267
rect 13955 4233 13967 4267
rect 13909 4227 13967 4233
rect 13924 4196 13952 4227
rect 14182 4224 14188 4276
rect 14240 4264 14246 4276
rect 14461 4267 14519 4273
rect 14461 4264 14473 4267
rect 14240 4236 14473 4264
rect 14240 4224 14246 4236
rect 14461 4233 14473 4236
rect 14507 4233 14519 4267
rect 14461 4227 14519 4233
rect 15562 4224 15568 4276
rect 15620 4224 15626 4276
rect 15749 4267 15807 4273
rect 15749 4233 15761 4267
rect 15795 4264 15807 4267
rect 15838 4264 15844 4276
rect 15795 4236 15844 4264
rect 15795 4233 15807 4236
rect 15749 4227 15807 4233
rect 15838 4224 15844 4236
rect 15896 4224 15902 4276
rect 16022 4224 16028 4276
rect 16080 4224 16086 4276
rect 16850 4224 16856 4276
rect 16908 4264 16914 4276
rect 16908 4236 17632 4264
rect 16908 4224 16914 4236
rect 14274 4196 14280 4208
rect 2746 4168 13952 4196
rect 14200 4168 14280 4196
rect 2406 4088 2412 4140
rect 2464 4088 2470 4140
rect 12986 4088 12992 4140
rect 13044 4128 13050 4140
rect 13111 4131 13169 4137
rect 13111 4128 13123 4131
rect 13044 4100 13123 4128
rect 13044 4088 13050 4100
rect 13111 4097 13123 4100
rect 13157 4097 13169 4131
rect 13633 4131 13691 4137
rect 13633 4128 13645 4131
rect 13111 4091 13169 4097
rect 13556 4100 13645 4128
rect 13556 4060 13584 4100
rect 13633 4097 13645 4100
rect 13679 4097 13691 4131
rect 13633 4091 13691 4097
rect 13725 4131 13783 4137
rect 13725 4097 13737 4131
rect 13771 4128 13783 4131
rect 14200 4128 14228 4168
rect 14274 4156 14280 4168
rect 14332 4156 14338 4208
rect 15580 4196 15608 4224
rect 16040 4196 16068 4224
rect 14384 4168 15608 4196
rect 15764 4168 16068 4196
rect 16224 4168 17356 4196
rect 14384 4137 14412 4168
rect 15764 4137 15792 4168
rect 13771 4100 14228 4128
rect 14369 4131 14427 4137
rect 13771 4097 13783 4100
rect 13725 4091 13783 4097
rect 14369 4097 14381 4131
rect 14415 4097 14427 4131
rect 14369 4091 14427 4097
rect 14553 4131 14611 4137
rect 14553 4097 14565 4131
rect 14599 4097 14611 4131
rect 14553 4091 14611 4097
rect 15565 4131 15623 4137
rect 15565 4097 15577 4131
rect 15611 4097 15623 4131
rect 15565 4091 15623 4097
rect 15749 4131 15807 4137
rect 15749 4097 15761 4131
rect 15795 4097 15807 4131
rect 15749 4091 15807 4097
rect 13096 4032 13584 4060
rect 3602 3952 3608 4004
rect 3660 3992 3666 4004
rect 12989 3995 13047 4001
rect 12989 3992 13001 3995
rect 3660 3964 13001 3992
rect 3660 3952 3666 3964
rect 12989 3961 13001 3964
rect 13035 3961 13047 3995
rect 12989 3955 13047 3961
rect 13096 3936 13124 4032
rect 13354 3952 13360 4004
rect 13412 3992 13418 4004
rect 13740 3992 13768 4091
rect 14090 4069 14096 4072
rect 14047 4063 14096 4069
rect 14047 4029 14059 4063
rect 14093 4029 14096 4063
rect 14047 4023 14096 4029
rect 14090 4020 14096 4023
rect 14148 4020 14154 4072
rect 13412 3964 13768 3992
rect 13412 3952 13418 3964
rect 2222 3884 2228 3936
rect 2280 3884 2286 3936
rect 13078 3884 13084 3936
rect 13136 3884 13142 3936
rect 13446 3884 13452 3936
rect 13504 3924 13510 3936
rect 13541 3927 13599 3933
rect 13541 3924 13553 3927
rect 13504 3896 13553 3924
rect 13504 3884 13510 3896
rect 13541 3893 13553 3896
rect 13587 3893 13599 3927
rect 13541 3887 13599 3893
rect 13906 3884 13912 3936
rect 13964 3924 13970 3936
rect 14277 3927 14335 3933
rect 14277 3924 14289 3927
rect 13964 3896 14289 3924
rect 13964 3884 13970 3896
rect 14277 3893 14289 3896
rect 14323 3924 14335 3927
rect 14384 3924 14412 4091
rect 14458 4020 14464 4072
rect 14516 4060 14522 4072
rect 14568 4060 14596 4091
rect 14516 4032 14596 4060
rect 15580 4060 15608 4091
rect 16022 4088 16028 4140
rect 16080 4088 16086 4140
rect 16224 4128 16252 4168
rect 16960 4140 16988 4168
rect 16132 4100 16252 4128
rect 16132 4060 16160 4100
rect 16298 4088 16304 4140
rect 16356 4088 16362 4140
rect 16574 4088 16580 4140
rect 16632 4128 16638 4140
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16632 4100 16681 4128
rect 16632 4088 16638 4100
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 16942 4088 16948 4140
rect 17000 4088 17006 4140
rect 17218 4088 17224 4140
rect 17276 4088 17282 4140
rect 17328 4137 17356 4168
rect 17604 4137 17632 4236
rect 17770 4224 17776 4276
rect 17828 4224 17834 4276
rect 19518 4224 19524 4276
rect 19576 4224 19582 4276
rect 19981 4267 20039 4273
rect 19981 4233 19993 4267
rect 20027 4264 20039 4267
rect 20438 4264 20444 4276
rect 20027 4236 20444 4264
rect 20027 4233 20039 4236
rect 19981 4227 20039 4233
rect 20438 4224 20444 4236
rect 20496 4224 20502 4276
rect 20530 4224 20536 4276
rect 20588 4224 20594 4276
rect 17788 4196 17816 4224
rect 17788 4168 17908 4196
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4097 17371 4131
rect 17313 4091 17371 4097
rect 17589 4131 17647 4137
rect 17589 4097 17601 4131
rect 17635 4097 17647 4131
rect 17880 4128 17908 4168
rect 18785 4131 18843 4137
rect 18785 4128 18797 4131
rect 17880 4100 18797 4128
rect 17589 4091 17647 4097
rect 18785 4097 18797 4100
rect 18831 4097 18843 4131
rect 18785 4091 18843 4097
rect 19242 4088 19248 4140
rect 19300 4088 19306 4140
rect 19426 4088 19432 4140
rect 19484 4088 19490 4140
rect 19536 4128 19564 4224
rect 19705 4131 19763 4137
rect 19705 4128 19717 4131
rect 19536 4100 19717 4128
rect 19705 4097 19717 4100
rect 19751 4097 19763 4131
rect 19705 4091 19763 4097
rect 19794 4088 19800 4140
rect 19852 4088 19858 4140
rect 20073 4131 20131 4137
rect 20073 4097 20085 4131
rect 20119 4128 20131 4131
rect 20548 4128 20576 4224
rect 24029 4199 24087 4205
rect 24029 4165 24041 4199
rect 24075 4196 24087 4199
rect 24213 4199 24271 4205
rect 24075 4168 24164 4196
rect 24075 4165 24087 4168
rect 24029 4159 24087 4165
rect 20119 4100 20576 4128
rect 24136 4128 24164 4168
rect 24213 4165 24225 4199
rect 24259 4196 24271 4199
rect 24302 4196 24308 4208
rect 24259 4168 24308 4196
rect 24259 4165 24271 4168
rect 24213 4159 24271 4165
rect 24302 4156 24308 4168
rect 24360 4196 24366 4208
rect 24765 4199 24823 4205
rect 24765 4196 24777 4199
rect 24360 4168 24777 4196
rect 24360 4156 24366 4168
rect 24765 4165 24777 4168
rect 24811 4165 24823 4199
rect 24765 4159 24823 4165
rect 24486 4128 24492 4140
rect 24136 4100 24492 4128
rect 20119 4097 20131 4100
rect 20073 4091 20131 4097
rect 24486 4088 24492 4100
rect 24544 4128 24550 4140
rect 24581 4131 24639 4137
rect 24581 4128 24593 4131
rect 24544 4100 24593 4128
rect 24544 4088 24550 4100
rect 24581 4097 24593 4100
rect 24627 4097 24639 4131
rect 24581 4091 24639 4097
rect 15580 4032 16160 4060
rect 16209 4063 16267 4069
rect 14516 4020 14522 4032
rect 16209 4029 16221 4063
rect 16255 4060 16267 4063
rect 17236 4060 17264 4088
rect 16255 4032 17264 4060
rect 16255 4029 16267 4032
rect 16209 4023 16267 4029
rect 17402 4020 17408 4072
rect 17460 4060 17466 4072
rect 19444 4060 19472 4088
rect 17460 4032 19472 4060
rect 17460 4020 17466 4032
rect 19518 4020 19524 4072
rect 19576 4020 19582 4072
rect 19610 4020 19616 4072
rect 19668 4060 19674 4072
rect 19981 4063 20039 4069
rect 19981 4060 19993 4063
rect 19668 4032 19993 4060
rect 19668 4020 19674 4032
rect 19981 4029 19993 4032
rect 20027 4029 20039 4063
rect 19981 4023 20039 4029
rect 15562 3952 15568 4004
rect 15620 3992 15626 4004
rect 22094 3992 22100 4004
rect 15620 3964 22100 3992
rect 15620 3952 15626 3964
rect 22094 3952 22100 3964
rect 22152 3952 22158 4004
rect 14323 3896 14412 3924
rect 14323 3893 14335 3896
rect 14277 3887 14335 3893
rect 14550 3884 14556 3936
rect 14608 3924 14614 3936
rect 15841 3927 15899 3933
rect 15841 3924 15853 3927
rect 14608 3896 15853 3924
rect 14608 3884 14614 3896
rect 15841 3893 15853 3896
rect 15887 3893 15899 3927
rect 15841 3887 15899 3893
rect 16022 3884 16028 3936
rect 16080 3924 16086 3936
rect 17034 3924 17040 3936
rect 16080 3896 17040 3924
rect 16080 3884 16086 3896
rect 17034 3884 17040 3896
rect 17092 3884 17098 3936
rect 17126 3884 17132 3936
rect 17184 3924 17190 3936
rect 18506 3924 18512 3936
rect 17184 3896 18512 3924
rect 17184 3884 17190 3896
rect 18506 3884 18512 3896
rect 18564 3884 18570 3936
rect 20162 3884 20168 3936
rect 20220 3884 20226 3936
rect 24394 3884 24400 3936
rect 24452 3884 24458 3936
rect 24946 3884 24952 3936
rect 25004 3884 25010 3936
rect 1104 3834 29440 3856
rect 1104 3782 4491 3834
rect 4543 3782 4555 3834
rect 4607 3782 4619 3834
rect 4671 3782 4683 3834
rect 4735 3782 4747 3834
rect 4799 3782 11574 3834
rect 11626 3782 11638 3834
rect 11690 3782 11702 3834
rect 11754 3782 11766 3834
rect 11818 3782 11830 3834
rect 11882 3782 18657 3834
rect 18709 3782 18721 3834
rect 18773 3782 18785 3834
rect 18837 3782 18849 3834
rect 18901 3782 18913 3834
rect 18965 3782 25740 3834
rect 25792 3782 25804 3834
rect 25856 3782 25868 3834
rect 25920 3782 25932 3834
rect 25984 3782 25996 3834
rect 26048 3782 29440 3834
rect 1104 3760 29440 3782
rect 2222 3680 2228 3732
rect 2280 3680 2286 3732
rect 12621 3723 12679 3729
rect 12621 3689 12633 3723
rect 12667 3720 12679 3723
rect 13170 3720 13176 3732
rect 12667 3692 13176 3720
rect 12667 3689 12679 3692
rect 12621 3683 12679 3689
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 14274 3680 14280 3732
rect 14332 3680 14338 3732
rect 14737 3723 14795 3729
rect 14737 3720 14749 3723
rect 14384 3692 14749 3720
rect 1489 3519 1547 3525
rect 1489 3485 1501 3519
rect 1535 3516 1547 3519
rect 2240 3516 2268 3680
rect 13538 3652 13544 3664
rect 13004 3624 13544 3652
rect 1535 3488 2268 3516
rect 2409 3519 2467 3525
rect 1535 3485 1547 3488
rect 1489 3479 1547 3485
rect 2409 3485 2421 3519
rect 2455 3516 2467 3519
rect 12529 3519 12587 3525
rect 2455 3488 2774 3516
rect 2455 3485 2467 3488
rect 2409 3479 2467 3485
rect 2746 3448 2774 3488
rect 12529 3485 12541 3519
rect 12575 3516 12587 3519
rect 12894 3516 12900 3528
rect 12575 3488 12900 3516
rect 12575 3485 12587 3488
rect 12529 3479 12587 3485
rect 12894 3476 12900 3488
rect 12952 3476 12958 3528
rect 13004 3525 13032 3624
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 13998 3612 14004 3664
rect 14056 3652 14062 3664
rect 14384 3652 14412 3692
rect 14737 3689 14749 3692
rect 14783 3689 14795 3723
rect 14737 3683 14795 3689
rect 15473 3723 15531 3729
rect 15473 3689 15485 3723
rect 15519 3720 15531 3723
rect 15562 3720 15568 3732
rect 15519 3692 15568 3720
rect 15519 3689 15531 3692
rect 15473 3683 15531 3689
rect 15562 3680 15568 3692
rect 15620 3680 15626 3732
rect 15654 3680 15660 3732
rect 15712 3720 15718 3732
rect 19518 3720 19524 3732
rect 15712 3692 19524 3720
rect 15712 3680 15718 3692
rect 19518 3680 19524 3692
rect 19576 3680 19582 3732
rect 24394 3720 24400 3732
rect 22066 3692 24400 3720
rect 14056 3624 14412 3652
rect 14056 3612 14062 3624
rect 14550 3612 14556 3664
rect 14608 3652 14614 3664
rect 15105 3655 15163 3661
rect 15105 3652 15117 3655
rect 14608 3624 15117 3652
rect 14608 3612 14614 3624
rect 15105 3621 15117 3624
rect 15151 3621 15163 3655
rect 15105 3615 15163 3621
rect 15194 3612 15200 3664
rect 15252 3652 15258 3664
rect 22066 3652 22094 3692
rect 24394 3680 24400 3692
rect 24452 3680 24458 3732
rect 24946 3680 24952 3732
rect 25004 3680 25010 3732
rect 15252 3624 22094 3652
rect 15252 3612 15258 3624
rect 14090 3584 14096 3596
rect 13740 3556 14096 3584
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3485 13047 3519
rect 12989 3479 13047 3485
rect 13265 3519 13323 3525
rect 13265 3485 13277 3519
rect 13311 3516 13323 3519
rect 13354 3516 13360 3528
rect 13311 3488 13360 3516
rect 13311 3485 13323 3488
rect 13265 3479 13323 3485
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 13446 3476 13452 3528
rect 13504 3476 13510 3528
rect 13740 3525 13768 3556
rect 14090 3544 14096 3556
rect 14148 3584 14154 3596
rect 14148 3556 15608 3584
rect 14148 3544 14154 3556
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3485 13783 3519
rect 13725 3479 13783 3485
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 14182 3516 14188 3528
rect 13872 3488 14188 3516
rect 13872 3476 13878 3488
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 14458 3476 14464 3528
rect 14516 3476 14522 3528
rect 14568 3525 14596 3556
rect 15580 3525 15608 3556
rect 15838 3544 15844 3596
rect 15896 3584 15902 3596
rect 15896 3556 17172 3584
rect 15896 3544 15902 3556
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 15381 3519 15439 3525
rect 15381 3485 15393 3519
rect 15427 3485 15439 3519
rect 15381 3479 15439 3485
rect 15565 3519 15623 3525
rect 15565 3485 15577 3519
rect 15611 3516 15623 3519
rect 15611 3488 16436 3516
rect 15611 3485 15623 3488
rect 15565 3479 15623 3485
rect 13170 3448 13176 3460
rect 2746 3420 13176 3448
rect 13170 3408 13176 3420
rect 13228 3408 13234 3460
rect 13464 3448 13492 3476
rect 13464 3420 13860 3448
rect 934 3340 940 3392
rect 992 3380 998 3392
rect 1581 3383 1639 3389
rect 1581 3380 1593 3383
rect 992 3352 1593 3380
rect 992 3340 998 3352
rect 1581 3349 1593 3352
rect 1627 3349 1639 3383
rect 1581 3343 1639 3349
rect 2222 3340 2228 3392
rect 2280 3340 2286 3392
rect 12802 3340 12808 3392
rect 12860 3340 12866 3392
rect 12894 3340 12900 3392
rect 12952 3380 12958 3392
rect 13722 3380 13728 3392
rect 12952 3352 13728 3380
rect 12952 3340 12958 3352
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 13832 3389 13860 3420
rect 13906 3408 13912 3460
rect 13964 3448 13970 3460
rect 14093 3451 14151 3457
rect 14093 3448 14105 3451
rect 13964 3420 14105 3448
rect 13964 3408 13970 3420
rect 14093 3417 14105 3420
rect 14139 3417 14151 3451
rect 14200 3448 14228 3476
rect 14829 3451 14887 3457
rect 14829 3448 14841 3451
rect 14200 3420 14841 3448
rect 14093 3411 14151 3417
rect 14829 3417 14841 3420
rect 14875 3417 14887 3451
rect 14829 3411 14887 3417
rect 13817 3383 13875 3389
rect 13817 3349 13829 3383
rect 13863 3380 13875 3383
rect 14274 3380 14280 3392
rect 13863 3352 14280 3380
rect 13863 3349 13875 3352
rect 13817 3343 13875 3349
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 14366 3340 14372 3392
rect 14424 3380 14430 3392
rect 14642 3380 14648 3392
rect 14424 3352 14648 3380
rect 14424 3340 14430 3352
rect 14642 3340 14648 3352
rect 14700 3340 14706 3392
rect 14918 3340 14924 3392
rect 14976 3380 14982 3392
rect 15289 3383 15347 3389
rect 15289 3380 15301 3383
rect 14976 3352 15301 3380
rect 14976 3340 14982 3352
rect 15289 3349 15301 3352
rect 15335 3380 15347 3383
rect 15396 3380 15424 3479
rect 16408 3457 16436 3488
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 16776 3525 16804 3556
rect 16669 3519 16727 3525
rect 16669 3516 16681 3519
rect 16632 3488 16681 3516
rect 16632 3476 16638 3488
rect 16669 3485 16681 3488
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 16761 3519 16819 3525
rect 16761 3485 16773 3519
rect 16807 3485 16819 3519
rect 16761 3479 16819 3485
rect 16853 3519 16911 3525
rect 16853 3485 16865 3519
rect 16899 3485 16911 3519
rect 16853 3479 16911 3485
rect 16393 3451 16451 3457
rect 16393 3417 16405 3451
rect 16439 3417 16451 3451
rect 16868 3448 16896 3479
rect 17034 3476 17040 3528
rect 17092 3476 17098 3528
rect 17144 3516 17172 3556
rect 17586 3544 17592 3596
rect 17644 3584 17650 3596
rect 18049 3587 18107 3593
rect 18049 3584 18061 3587
rect 17644 3556 18061 3584
rect 17644 3544 17650 3556
rect 18049 3553 18061 3556
rect 18095 3553 18107 3587
rect 18049 3547 18107 3553
rect 18969 3587 19027 3593
rect 18969 3553 18981 3587
rect 19015 3584 19027 3587
rect 20162 3584 20168 3596
rect 19015 3556 20168 3584
rect 19015 3553 19027 3556
rect 18969 3547 19027 3553
rect 20162 3544 20168 3556
rect 20220 3544 20226 3596
rect 17144 3488 17908 3516
rect 16868 3420 17632 3448
rect 16393 3411 16451 3417
rect 17604 3392 17632 3420
rect 17770 3408 17776 3460
rect 17828 3448 17834 3460
rect 17880 3457 17908 3488
rect 18506 3476 18512 3528
rect 18564 3516 18570 3528
rect 18693 3519 18751 3525
rect 18693 3516 18705 3519
rect 18564 3488 18705 3516
rect 18564 3476 18570 3488
rect 18693 3485 18705 3488
rect 18739 3485 18751 3519
rect 24964 3516 24992 3680
rect 25409 3519 25467 3525
rect 25409 3516 25421 3519
rect 24964 3488 25421 3516
rect 18693 3479 18751 3485
rect 25409 3485 25421 3488
rect 25455 3485 25467 3519
rect 25409 3479 25467 3485
rect 17865 3451 17923 3457
rect 17865 3448 17877 3451
rect 17828 3420 17877 3448
rect 17828 3408 17834 3420
rect 17865 3417 17877 3420
rect 17911 3417 17923 3451
rect 17865 3411 17923 3417
rect 15335 3352 15424 3380
rect 15335 3349 15347 3352
rect 15289 3343 15347 3349
rect 17494 3340 17500 3392
rect 17552 3340 17558 3392
rect 17586 3340 17592 3392
rect 17644 3340 17650 3392
rect 17957 3383 18015 3389
rect 17957 3349 17969 3383
rect 18003 3380 18015 3383
rect 18325 3383 18383 3389
rect 18325 3380 18337 3383
rect 18003 3352 18337 3380
rect 18003 3349 18015 3352
rect 17957 3343 18015 3349
rect 18325 3349 18337 3352
rect 18371 3349 18383 3383
rect 18325 3343 18383 3349
rect 18782 3340 18788 3392
rect 18840 3340 18846 3392
rect 25222 3340 25228 3392
rect 25280 3340 25286 3392
rect 1104 3290 29595 3312
rect 1104 3238 8032 3290
rect 8084 3238 8096 3290
rect 8148 3238 8160 3290
rect 8212 3238 8224 3290
rect 8276 3238 8288 3290
rect 8340 3238 15115 3290
rect 15167 3238 15179 3290
rect 15231 3238 15243 3290
rect 15295 3238 15307 3290
rect 15359 3238 15371 3290
rect 15423 3238 22198 3290
rect 22250 3238 22262 3290
rect 22314 3238 22326 3290
rect 22378 3238 22390 3290
rect 22442 3238 22454 3290
rect 22506 3238 29281 3290
rect 29333 3238 29345 3290
rect 29397 3238 29409 3290
rect 29461 3238 29473 3290
rect 29525 3238 29537 3290
rect 29589 3238 29595 3290
rect 1104 3216 29595 3238
rect 12986 3136 12992 3188
rect 13044 3136 13050 3188
rect 13078 3136 13084 3188
rect 13136 3176 13142 3188
rect 14550 3176 14556 3188
rect 13136 3148 14556 3176
rect 13136 3136 13142 3148
rect 13372 3049 13400 3148
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 15654 3136 15660 3188
rect 15712 3136 15718 3188
rect 17494 3136 17500 3188
rect 17552 3136 17558 3188
rect 17586 3136 17592 3188
rect 17644 3136 17650 3188
rect 17770 3136 17776 3188
rect 17828 3136 17834 3188
rect 17957 3179 18015 3185
rect 17957 3145 17969 3179
rect 18003 3176 18015 3179
rect 18782 3176 18788 3188
rect 18003 3148 18788 3176
rect 18003 3145 18015 3148
rect 17957 3139 18015 3145
rect 18782 3136 18788 3148
rect 18840 3136 18846 3188
rect 14090 3108 14096 3120
rect 13464 3080 14096 3108
rect 13464 3049 13492 3080
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 14918 3108 14924 3120
rect 14200 3080 14924 3108
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3009 13139 3043
rect 13081 3003 13139 3009
rect 13357 3043 13415 3049
rect 13357 3009 13369 3043
rect 13403 3009 13415 3043
rect 13357 3003 13415 3009
rect 13449 3043 13507 3049
rect 13449 3009 13461 3043
rect 13495 3009 13507 3043
rect 13449 3003 13507 3009
rect 12912 2904 12940 3003
rect 13096 2972 13124 3003
rect 13464 2972 13492 3003
rect 13538 3000 13544 3052
rect 13596 3040 13602 3052
rect 13633 3043 13691 3049
rect 13633 3040 13645 3043
rect 13596 3012 13645 3040
rect 13596 3000 13602 3012
rect 13633 3009 13645 3012
rect 13679 3009 13691 3043
rect 13633 3003 13691 3009
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 13096 2944 13492 2972
rect 13354 2904 13360 2916
rect 12912 2876 13360 2904
rect 13354 2864 13360 2876
rect 13412 2864 13418 2916
rect 13740 2848 13768 3003
rect 13906 3000 13912 3052
rect 13964 3000 13970 3052
rect 13998 3000 14004 3052
rect 14056 3000 14062 3052
rect 14200 3049 14228 3080
rect 14918 3068 14924 3080
rect 14976 3068 14982 3120
rect 14185 3043 14243 3049
rect 14185 3009 14197 3043
rect 14231 3009 14243 3043
rect 14185 3003 14243 3009
rect 14274 3000 14280 3052
rect 14332 3000 14338 3052
rect 14369 3043 14427 3049
rect 14369 3009 14381 3043
rect 14415 3009 14427 3043
rect 14369 3003 14427 3009
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3040 14611 3043
rect 14642 3040 14648 3052
rect 14599 3012 14648 3040
rect 14599 3009 14611 3012
rect 14553 3003 14611 3009
rect 13924 2972 13952 3000
rect 14384 2972 14412 3003
rect 14642 3000 14648 3012
rect 14700 3040 14706 3052
rect 15672 3040 15700 3136
rect 16868 3080 17172 3108
rect 16868 3049 16896 3080
rect 17144 3052 17172 3080
rect 14700 3012 15700 3040
rect 16853 3043 16911 3049
rect 14700 3000 14706 3012
rect 16853 3009 16865 3043
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 17034 3000 17040 3052
rect 17092 3000 17098 3052
rect 17126 3000 17132 3052
rect 17184 3000 17190 3052
rect 17221 3043 17279 3049
rect 17221 3009 17233 3043
rect 17267 3040 17279 3043
rect 17512 3040 17540 3136
rect 17788 3049 17816 3136
rect 17267 3012 17540 3040
rect 17681 3043 17739 3049
rect 17267 3009 17279 3012
rect 17221 3003 17279 3009
rect 17681 3009 17693 3043
rect 17727 3009 17739 3043
rect 17681 3003 17739 3009
rect 17773 3043 17831 3049
rect 17773 3009 17785 3043
rect 17819 3009 17831 3043
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 17773 3003 17831 3009
rect 17880 3012 18061 3040
rect 13924 2944 14412 2972
rect 16945 2975 17003 2981
rect 16945 2941 16957 2975
rect 16991 2972 17003 2975
rect 17405 2975 17463 2981
rect 17405 2972 17417 2975
rect 16991 2944 17417 2972
rect 16991 2941 17003 2944
rect 16945 2935 17003 2941
rect 17405 2941 17417 2944
rect 17451 2941 17463 2975
rect 17405 2935 17463 2941
rect 17494 2932 17500 2984
rect 17552 2932 17558 2984
rect 17696 2972 17724 3003
rect 17880 2972 17908 3012
rect 18049 3009 18061 3012
rect 18095 3040 18107 3043
rect 18138 3040 18144 3052
rect 18095 3012 18144 3040
rect 18095 3009 18107 3012
rect 18049 3003 18107 3009
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 18230 3000 18236 3052
rect 18288 3000 18294 3052
rect 28813 3043 28871 3049
rect 28813 3040 28825 3043
rect 22066 3012 28825 3040
rect 17696 2944 17908 2972
rect 17954 2932 17960 2984
rect 18012 2932 18018 2984
rect 13817 2907 13875 2913
rect 13817 2873 13829 2907
rect 13863 2904 13875 2907
rect 22066 2904 22094 3012
rect 28813 3009 28825 3012
rect 28859 3009 28871 3043
rect 28813 3003 28871 3009
rect 13863 2876 22094 2904
rect 13863 2873 13875 2876
rect 13817 2867 13875 2873
rect 13170 2796 13176 2848
rect 13228 2796 13234 2848
rect 13722 2796 13728 2848
rect 13780 2836 13786 2848
rect 14458 2836 14464 2848
rect 13780 2808 14464 2836
rect 13780 2796 13786 2808
rect 14458 2796 14464 2808
rect 14516 2796 14522 2848
rect 17126 2796 17132 2848
rect 17184 2836 17190 2848
rect 18049 2839 18107 2845
rect 18049 2836 18061 2839
rect 17184 2808 18061 2836
rect 17184 2796 17190 2808
rect 18049 2805 18061 2808
rect 18095 2836 18107 2839
rect 19794 2836 19800 2848
rect 18095 2808 19800 2836
rect 18095 2805 18107 2808
rect 18049 2799 18107 2805
rect 19794 2796 19800 2808
rect 19852 2796 19858 2848
rect 28994 2796 29000 2848
rect 29052 2796 29058 2848
rect 1104 2746 29440 2768
rect 1104 2694 4491 2746
rect 4543 2694 4555 2746
rect 4607 2694 4619 2746
rect 4671 2694 4683 2746
rect 4735 2694 4747 2746
rect 4799 2694 11574 2746
rect 11626 2694 11638 2746
rect 11690 2694 11702 2746
rect 11754 2694 11766 2746
rect 11818 2694 11830 2746
rect 11882 2694 18657 2746
rect 18709 2694 18721 2746
rect 18773 2694 18785 2746
rect 18837 2694 18849 2746
rect 18901 2694 18913 2746
rect 18965 2694 25740 2746
rect 25792 2694 25804 2746
rect 25856 2694 25868 2746
rect 25920 2694 25932 2746
rect 25984 2694 25996 2746
rect 26048 2694 29440 2746
rect 1104 2672 29440 2694
rect 12802 2632 12808 2644
rect 6886 2604 12808 2632
rect 1489 2431 1547 2437
rect 1489 2397 1501 2431
rect 1535 2428 1547 2431
rect 2222 2428 2228 2440
rect 1535 2400 2228 2428
rect 1535 2397 1547 2400
rect 1489 2391 1547 2397
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 3881 2431 3939 2437
rect 3881 2397 3893 2431
rect 3927 2428 3939 2431
rect 6886 2428 6914 2604
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 13262 2592 13268 2644
rect 13320 2632 13326 2644
rect 13449 2635 13507 2641
rect 13449 2632 13461 2635
rect 13320 2604 13461 2632
rect 13320 2592 13326 2604
rect 13449 2601 13461 2604
rect 13495 2601 13507 2635
rect 13449 2595 13507 2601
rect 27062 2564 27068 2576
rect 16546 2536 27068 2564
rect 3927 2400 6914 2428
rect 7300 2468 13216 2496
rect 3927 2397 3939 2400
rect 3881 2391 3939 2397
rect 7300 2369 7328 2468
rect 13188 2440 13216 2468
rect 13170 2388 13176 2440
rect 13228 2388 13234 2440
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2428 13507 2431
rect 13538 2428 13544 2440
rect 13495 2400 13544 2428
rect 13495 2397 13507 2400
rect 13449 2391 13507 2397
rect 13538 2388 13544 2400
rect 13596 2388 13602 2440
rect 13633 2431 13691 2437
rect 13633 2397 13645 2431
rect 13679 2428 13691 2431
rect 13722 2428 13728 2440
rect 13679 2400 13728 2428
rect 13679 2397 13691 2400
rect 13633 2391 13691 2397
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 15013 2431 15071 2437
rect 15013 2397 15025 2431
rect 15059 2428 15071 2431
rect 16546 2428 16574 2536
rect 27062 2524 27068 2536
rect 27120 2524 27126 2576
rect 15059 2400 16574 2428
rect 15059 2397 15071 2400
rect 15013 2391 15071 2397
rect 19334 2388 19340 2440
rect 19392 2388 19398 2440
rect 22094 2388 22100 2440
rect 22152 2388 22158 2440
rect 25222 2388 25228 2440
rect 25280 2428 25286 2440
rect 25961 2431 26019 2437
rect 25961 2428 25973 2431
rect 25280 2400 25973 2428
rect 25280 2388 25286 2400
rect 25961 2397 25973 2400
rect 26007 2397 26019 2431
rect 25961 2391 26019 2397
rect 28534 2388 28540 2440
rect 28592 2428 28598 2440
rect 28721 2431 28779 2437
rect 28721 2428 28733 2431
rect 28592 2400 28733 2428
rect 28592 2388 28598 2400
rect 28721 2397 28733 2400
rect 28767 2397 28779 2431
rect 28721 2391 28779 2397
rect 7285 2363 7343 2369
rect 7285 2329 7297 2363
rect 7331 2329 7343 2363
rect 7285 2323 7343 2329
rect 11609 2363 11667 2369
rect 11609 2329 11621 2363
rect 11655 2360 11667 2363
rect 17494 2360 17500 2372
rect 11655 2332 17500 2360
rect 11655 2329 11667 2332
rect 11609 2323 11667 2329
rect 17494 2320 17500 2332
rect 17552 2320 17558 2372
rect 29089 2363 29147 2369
rect 29089 2329 29101 2363
rect 29135 2360 29147 2363
rect 29638 2360 29644 2372
rect 29135 2332 29644 2360
rect 29135 2329 29147 2332
rect 29089 2323 29147 2329
rect 29638 2320 29644 2332
rect 29696 2320 29702 2372
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 1581 2295 1639 2301
rect 1581 2292 1593 2295
rect 72 2264 1593 2292
rect 72 2252 78 2264
rect 1581 2261 1593 2264
rect 1627 2261 1639 2295
rect 1581 2255 1639 2261
rect 3418 2252 3424 2304
rect 3476 2292 3482 2304
rect 4157 2295 4215 2301
rect 4157 2292 4169 2295
rect 3476 2264 4169 2292
rect 3476 2252 3482 2264
rect 4157 2261 4169 2264
rect 4203 2261 4215 2295
rect 4157 2255 4215 2261
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7377 2295 7435 2301
rect 7377 2292 7389 2295
rect 7156 2264 7389 2292
rect 7156 2252 7162 2264
rect 7377 2261 7389 2264
rect 7423 2261 7435 2295
rect 7377 2255 7435 2261
rect 11146 2252 11152 2304
rect 11204 2292 11210 2304
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 11204 2264 11713 2292
rect 11204 2252 11210 2264
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 11701 2255 11759 2261
rect 14918 2252 14924 2304
rect 14976 2292 14982 2304
rect 15289 2295 15347 2301
rect 15289 2292 15301 2295
rect 14976 2264 15301 2292
rect 14976 2252 14982 2264
rect 15289 2261 15301 2264
rect 15335 2261 15347 2295
rect 15289 2255 15347 2261
rect 19058 2252 19064 2304
rect 19116 2292 19122 2304
rect 19429 2295 19487 2301
rect 19429 2292 19441 2295
rect 19116 2264 19441 2292
rect 19116 2252 19122 2264
rect 19429 2261 19441 2264
rect 19475 2261 19487 2295
rect 19429 2255 19487 2261
rect 22002 2252 22008 2304
rect 22060 2292 22066 2304
rect 22189 2295 22247 2301
rect 22189 2292 22201 2295
rect 22060 2264 22201 2292
rect 22060 2252 22066 2264
rect 22189 2261 22201 2264
rect 22235 2261 22247 2295
rect 22189 2255 22247 2261
rect 26142 2252 26148 2304
rect 26200 2292 26206 2304
rect 26237 2295 26295 2301
rect 26237 2292 26249 2295
rect 26200 2264 26249 2292
rect 26200 2252 26206 2264
rect 26237 2261 26249 2264
rect 26283 2261 26295 2295
rect 26237 2255 26295 2261
rect 1104 2202 29595 2224
rect 1104 2150 8032 2202
rect 8084 2150 8096 2202
rect 8148 2150 8160 2202
rect 8212 2150 8224 2202
rect 8276 2150 8288 2202
rect 8340 2150 15115 2202
rect 15167 2150 15179 2202
rect 15231 2150 15243 2202
rect 15295 2150 15307 2202
rect 15359 2150 15371 2202
rect 15423 2150 22198 2202
rect 22250 2150 22262 2202
rect 22314 2150 22326 2202
rect 22378 2150 22390 2202
rect 22442 2150 22454 2202
rect 22506 2150 29281 2202
rect 29333 2150 29345 2202
rect 29397 2150 29409 2202
rect 29461 2150 29473 2202
rect 29525 2150 29537 2202
rect 29589 2150 29595 2202
rect 1104 2128 29595 2150
<< via1 >>
rect 8032 30438 8084 30490
rect 8096 30438 8148 30490
rect 8160 30438 8212 30490
rect 8224 30438 8276 30490
rect 8288 30438 8340 30490
rect 15115 30438 15167 30490
rect 15179 30438 15231 30490
rect 15243 30438 15295 30490
rect 15307 30438 15359 30490
rect 15371 30438 15423 30490
rect 22198 30438 22250 30490
rect 22262 30438 22314 30490
rect 22326 30438 22378 30490
rect 22390 30438 22442 30490
rect 22454 30438 22506 30490
rect 29281 30438 29333 30490
rect 29345 30438 29397 30490
rect 29409 30438 29461 30490
rect 29473 30438 29525 30490
rect 29537 30438 29589 30490
rect 6736 30379 6788 30388
rect 6736 30345 6745 30379
rect 6745 30345 6779 30379
rect 6779 30345 6788 30379
rect 6736 30336 6788 30345
rect 9680 30268 9732 30320
rect 21272 30268 21324 30320
rect 25412 30268 25464 30320
rect 1584 30243 1636 30252
rect 1584 30209 1593 30243
rect 1593 30209 1627 30243
rect 1627 30209 1636 30243
rect 1584 30200 1636 30209
rect 3424 30200 3476 30252
rect 6092 30200 6144 30252
rect 9864 30243 9916 30252
rect 9864 30209 9873 30243
rect 9873 30209 9907 30243
rect 9907 30209 9916 30243
rect 9864 30200 9916 30209
rect 14188 30243 14240 30252
rect 14188 30209 14197 30243
rect 14197 30209 14231 30243
rect 14231 30209 14240 30243
rect 14188 30200 14240 30209
rect 17592 30243 17644 30252
rect 17592 30209 17601 30243
rect 17601 30209 17635 30243
rect 17635 30209 17644 30243
rect 17592 30200 17644 30209
rect 21916 30243 21968 30252
rect 21916 30209 21925 30243
rect 21925 30209 21959 30243
rect 21959 30209 21968 30243
rect 21916 30200 21968 30209
rect 25320 30243 25372 30252
rect 25320 30209 25329 30243
rect 25329 30209 25363 30243
rect 25363 30209 25372 30243
rect 25320 30200 25372 30209
rect 29000 30268 29052 30320
rect 28724 30243 28776 30252
rect 28724 30209 28733 30243
rect 28733 30209 28767 30243
rect 28767 30209 28776 30243
rect 28724 30200 28776 30209
rect 28908 30132 28960 30184
rect 2780 30064 2832 30116
rect 13820 30064 13872 30116
rect 17408 30064 17460 30116
rect 1584 29996 1636 30048
rect 28540 30039 28592 30048
rect 28540 30005 28549 30039
rect 28549 30005 28583 30039
rect 28583 30005 28592 30039
rect 28540 29996 28592 30005
rect 4491 29894 4543 29946
rect 4555 29894 4607 29946
rect 4619 29894 4671 29946
rect 4683 29894 4735 29946
rect 4747 29894 4799 29946
rect 11574 29894 11626 29946
rect 11638 29894 11690 29946
rect 11702 29894 11754 29946
rect 11766 29894 11818 29946
rect 11830 29894 11882 29946
rect 18657 29894 18709 29946
rect 18721 29894 18773 29946
rect 18785 29894 18837 29946
rect 18849 29894 18901 29946
rect 18913 29894 18965 29946
rect 25740 29894 25792 29946
rect 25804 29894 25856 29946
rect 25868 29894 25920 29946
rect 25932 29894 25984 29946
rect 25996 29894 26048 29946
rect 21916 29792 21968 29844
rect 5080 29724 5132 29776
rect 5448 29724 5500 29776
rect 5356 29588 5408 29640
rect 14096 29656 14148 29708
rect 5724 29631 5776 29640
rect 5724 29597 5733 29631
rect 5733 29597 5767 29631
rect 5767 29597 5776 29631
rect 5724 29588 5776 29597
rect 9036 29631 9088 29640
rect 9036 29597 9045 29631
rect 9045 29597 9079 29631
rect 9079 29597 9088 29631
rect 9036 29588 9088 29597
rect 11336 29588 11388 29640
rect 13268 29588 13320 29640
rect 16212 29656 16264 29708
rect 19156 29656 19208 29708
rect 6000 29520 6052 29572
rect 7380 29563 7432 29572
rect 7380 29529 7389 29563
rect 7389 29529 7423 29563
rect 7423 29529 7432 29563
rect 7380 29520 7432 29529
rect 7564 29563 7616 29572
rect 7564 29529 7573 29563
rect 7573 29529 7607 29563
rect 7607 29529 7616 29563
rect 7564 29520 7616 29529
rect 9404 29563 9456 29572
rect 9404 29529 9413 29563
rect 9413 29529 9447 29563
rect 9447 29529 9456 29563
rect 9404 29520 9456 29529
rect 12256 29520 12308 29572
rect 14280 29520 14332 29572
rect 16488 29520 16540 29572
rect 20812 29631 20864 29640
rect 20812 29597 20821 29631
rect 20821 29597 20855 29631
rect 20855 29597 20864 29631
rect 20812 29588 20864 29597
rect 25228 29588 25280 29640
rect 4896 29495 4948 29504
rect 4896 29461 4905 29495
rect 4905 29461 4939 29495
rect 4939 29461 4948 29495
rect 4896 29452 4948 29461
rect 5816 29452 5868 29504
rect 7748 29495 7800 29504
rect 7748 29461 7757 29495
rect 7757 29461 7791 29495
rect 7791 29461 7800 29495
rect 7748 29452 7800 29461
rect 11060 29452 11112 29504
rect 11244 29452 11296 29504
rect 17132 29452 17184 29504
rect 17316 29495 17368 29504
rect 17316 29461 17325 29495
rect 17325 29461 17359 29495
rect 17359 29461 17368 29495
rect 17316 29452 17368 29461
rect 19248 29452 19300 29504
rect 20444 29452 20496 29504
rect 8032 29350 8084 29402
rect 8096 29350 8148 29402
rect 8160 29350 8212 29402
rect 8224 29350 8276 29402
rect 8288 29350 8340 29402
rect 15115 29350 15167 29402
rect 15179 29350 15231 29402
rect 15243 29350 15295 29402
rect 15307 29350 15359 29402
rect 15371 29350 15423 29402
rect 22198 29350 22250 29402
rect 22262 29350 22314 29402
rect 22326 29350 22378 29402
rect 22390 29350 22442 29402
rect 22454 29350 22506 29402
rect 29281 29350 29333 29402
rect 29345 29350 29397 29402
rect 29409 29350 29461 29402
rect 29473 29350 29525 29402
rect 29537 29350 29589 29402
rect 3240 29248 3292 29300
rect 1584 29180 1636 29232
rect 3976 29180 4028 29232
rect 7104 29248 7156 29300
rect 9404 29248 9456 29300
rect 11244 29248 11296 29300
rect 3240 29155 3292 29164
rect 3240 29121 3249 29155
rect 3249 29121 3283 29155
rect 3283 29121 3292 29155
rect 3240 29112 3292 29121
rect 6828 29155 6880 29164
rect 6828 29121 6837 29155
rect 6837 29121 6871 29155
rect 6871 29121 6880 29155
rect 6828 29112 6880 29121
rect 3516 29087 3568 29096
rect 3516 29053 3525 29087
rect 3525 29053 3559 29087
rect 3559 29053 3568 29087
rect 3516 29044 3568 29053
rect 5448 29044 5500 29096
rect 7472 29180 7524 29232
rect 8484 29180 8536 29232
rect 9772 29180 9824 29232
rect 3148 29019 3200 29028
rect 3148 28985 3157 29019
rect 3157 28985 3191 29019
rect 3191 28985 3200 29019
rect 3148 28976 3200 28985
rect 4160 28908 4212 28960
rect 5172 28976 5224 29028
rect 7564 29044 7616 29096
rect 12624 29248 12676 29300
rect 13268 29291 13320 29300
rect 13268 29257 13277 29291
rect 13277 29257 13311 29291
rect 13311 29257 13320 29291
rect 13268 29248 13320 29257
rect 16488 29291 16540 29300
rect 16488 29257 16497 29291
rect 16497 29257 16531 29291
rect 16531 29257 16540 29291
rect 16488 29248 16540 29257
rect 12256 29180 12308 29232
rect 14280 29180 14332 29232
rect 16212 29155 16264 29164
rect 16212 29121 16221 29155
rect 16221 29121 16255 29155
rect 16255 29121 16264 29155
rect 16212 29112 16264 29121
rect 16672 29180 16724 29232
rect 17316 29248 17368 29300
rect 19156 29291 19208 29300
rect 19156 29257 19165 29291
rect 19165 29257 19199 29291
rect 19199 29257 19208 29291
rect 19156 29248 19208 29257
rect 19248 29248 19300 29300
rect 20444 29180 20496 29232
rect 20720 29180 20772 29232
rect 18052 29112 18104 29164
rect 11244 29044 11296 29096
rect 13452 29087 13504 29096
rect 13452 29053 13461 29087
rect 13461 29053 13495 29087
rect 13495 29053 13504 29087
rect 13452 29044 13504 29053
rect 13728 29087 13780 29096
rect 13728 29053 13737 29087
rect 13737 29053 13771 29087
rect 13771 29053 13780 29087
rect 13728 29044 13780 29053
rect 5080 28908 5132 28960
rect 5264 28908 5316 28960
rect 6920 28908 6972 28960
rect 7196 28908 7248 28960
rect 7380 28908 7432 28960
rect 7840 28908 7892 28960
rect 8760 28951 8812 28960
rect 8760 28917 8769 28951
rect 8769 28917 8803 28951
rect 8803 28917 8812 28951
rect 8760 28908 8812 28917
rect 11152 28951 11204 28960
rect 11152 28917 11161 28951
rect 11161 28917 11195 28951
rect 11195 28917 11204 28951
rect 11152 28908 11204 28917
rect 16580 29044 16632 29096
rect 18420 29044 18472 29096
rect 22836 29112 22888 29164
rect 20168 29044 20220 29096
rect 22100 29044 22152 29096
rect 23388 29087 23440 29096
rect 23388 29053 23397 29087
rect 23397 29053 23431 29087
rect 23431 29053 23440 29087
rect 23388 29044 23440 29053
rect 28540 29248 28592 29300
rect 24492 29044 24544 29096
rect 15568 28908 15620 28960
rect 15936 28951 15988 28960
rect 15936 28917 15945 28951
rect 15945 28917 15979 28951
rect 15979 28917 15988 28951
rect 15936 28908 15988 28917
rect 18328 28908 18380 28960
rect 20720 28908 20772 28960
rect 21364 28908 21416 28960
rect 22928 28908 22980 28960
rect 23204 28976 23256 29028
rect 23112 28951 23164 28960
rect 23112 28917 23121 28951
rect 23121 28917 23155 28951
rect 23155 28917 23164 28951
rect 23112 28908 23164 28917
rect 4491 28806 4543 28858
rect 4555 28806 4607 28858
rect 4619 28806 4671 28858
rect 4683 28806 4735 28858
rect 4747 28806 4799 28858
rect 11574 28806 11626 28858
rect 11638 28806 11690 28858
rect 11702 28806 11754 28858
rect 11766 28806 11818 28858
rect 11830 28806 11882 28858
rect 18657 28806 18709 28858
rect 18721 28806 18773 28858
rect 18785 28806 18837 28858
rect 18849 28806 18901 28858
rect 18913 28806 18965 28858
rect 25740 28806 25792 28858
rect 25804 28806 25856 28858
rect 25868 28806 25920 28858
rect 25932 28806 25984 28858
rect 25996 28806 26048 28858
rect 5172 28704 5224 28756
rect 5724 28704 5776 28756
rect 4252 28568 4304 28620
rect 4988 28568 5040 28620
rect 6368 28568 6420 28620
rect 4160 28500 4212 28552
rect 3608 28407 3660 28416
rect 3608 28373 3617 28407
rect 3617 28373 3651 28407
rect 3651 28373 3660 28407
rect 3608 28364 3660 28373
rect 4160 28364 4212 28416
rect 4344 28364 4396 28416
rect 4896 28432 4948 28484
rect 5264 28432 5316 28484
rect 6184 28475 6236 28484
rect 6184 28441 6193 28475
rect 6193 28441 6227 28475
rect 6227 28441 6236 28475
rect 6184 28432 6236 28441
rect 7748 28704 7800 28756
rect 6460 28543 6512 28552
rect 6460 28509 6469 28543
rect 6469 28509 6503 28543
rect 6503 28509 6512 28543
rect 6460 28500 6512 28509
rect 7288 28500 7340 28552
rect 7564 28500 7616 28552
rect 5356 28364 5408 28416
rect 7196 28475 7248 28484
rect 7196 28441 7205 28475
rect 7205 28441 7239 28475
rect 7239 28441 7248 28475
rect 7196 28432 7248 28441
rect 7012 28407 7064 28416
rect 7012 28373 7021 28407
rect 7021 28373 7055 28407
rect 7055 28373 7064 28407
rect 7012 28364 7064 28373
rect 7104 28364 7156 28416
rect 7288 28364 7340 28416
rect 7840 28475 7892 28484
rect 7840 28441 7865 28475
rect 7865 28441 7892 28475
rect 7840 28432 7892 28441
rect 8760 28568 8812 28620
rect 9772 28747 9824 28756
rect 9772 28713 9781 28747
rect 9781 28713 9815 28747
rect 9815 28713 9824 28747
rect 9772 28704 9824 28713
rect 12624 28747 12676 28756
rect 12624 28713 12633 28747
rect 12633 28713 12667 28747
rect 12667 28713 12676 28747
rect 12624 28704 12676 28713
rect 12900 28704 12952 28756
rect 13728 28704 13780 28756
rect 16212 28704 16264 28756
rect 16672 28747 16724 28756
rect 16672 28713 16681 28747
rect 16681 28713 16715 28747
rect 16715 28713 16724 28747
rect 16672 28704 16724 28713
rect 9404 28568 9456 28620
rect 11152 28568 11204 28620
rect 11244 28568 11296 28620
rect 10416 28543 10468 28552
rect 10416 28509 10425 28543
rect 10425 28509 10459 28543
rect 10459 28509 10468 28543
rect 10416 28500 10468 28509
rect 9956 28475 10008 28484
rect 9956 28441 9965 28475
rect 9965 28441 9999 28475
rect 9999 28441 10008 28475
rect 9956 28432 10008 28441
rect 8576 28364 8628 28416
rect 11152 28432 11204 28484
rect 13636 28611 13688 28620
rect 13636 28577 13645 28611
rect 13645 28577 13679 28611
rect 13679 28577 13688 28611
rect 13636 28568 13688 28577
rect 15936 28568 15988 28620
rect 13360 28543 13412 28552
rect 13360 28509 13369 28543
rect 13369 28509 13403 28543
rect 13403 28509 13412 28543
rect 13360 28500 13412 28509
rect 14004 28500 14056 28552
rect 14464 28500 14516 28552
rect 12164 28407 12216 28416
rect 12164 28373 12173 28407
rect 12173 28373 12207 28407
rect 12207 28373 12216 28407
rect 12164 28364 12216 28373
rect 13636 28432 13688 28484
rect 15568 28543 15620 28552
rect 15568 28509 15577 28543
rect 15577 28509 15611 28543
rect 15611 28509 15620 28543
rect 15568 28500 15620 28509
rect 18144 28636 18196 28688
rect 19248 28636 19300 28688
rect 19340 28636 19392 28688
rect 20812 28704 20864 28756
rect 21272 28704 21324 28756
rect 22376 28704 22428 28756
rect 22928 28704 22980 28756
rect 17132 28568 17184 28620
rect 16488 28543 16540 28552
rect 16488 28509 16497 28543
rect 16497 28509 16531 28543
rect 16531 28509 16540 28543
rect 16488 28500 16540 28509
rect 16580 28500 16632 28552
rect 16304 28475 16356 28484
rect 12348 28364 12400 28416
rect 13912 28407 13964 28416
rect 13912 28373 13921 28407
rect 13921 28373 13955 28407
rect 13955 28373 13964 28407
rect 13912 28364 13964 28373
rect 14740 28407 14792 28416
rect 14740 28373 14749 28407
rect 14749 28373 14783 28407
rect 14783 28373 14792 28407
rect 14740 28364 14792 28373
rect 15016 28364 15068 28416
rect 16304 28441 16313 28475
rect 16313 28441 16347 28475
rect 16347 28441 16356 28475
rect 16304 28432 16356 28441
rect 19432 28500 19484 28552
rect 20168 28568 20220 28620
rect 20812 28543 20864 28552
rect 20812 28509 20821 28543
rect 20821 28509 20855 28543
rect 20855 28509 20864 28543
rect 20812 28500 20864 28509
rect 21364 28543 21416 28552
rect 18052 28364 18104 28416
rect 18420 28364 18472 28416
rect 19432 28364 19484 28416
rect 20260 28364 20312 28416
rect 21364 28509 21373 28543
rect 21373 28509 21407 28543
rect 21407 28509 21416 28543
rect 21364 28500 21416 28509
rect 21640 28500 21692 28552
rect 21824 28543 21876 28552
rect 21824 28509 21857 28543
rect 21857 28509 21876 28543
rect 21824 28500 21876 28509
rect 21272 28364 21324 28416
rect 21364 28364 21416 28416
rect 22376 28543 22428 28552
rect 22376 28509 22385 28543
rect 22385 28509 22419 28543
rect 22419 28509 22428 28543
rect 22376 28500 22428 28509
rect 22100 28475 22152 28484
rect 22100 28441 22109 28475
rect 22109 28441 22143 28475
rect 22143 28441 22152 28475
rect 22100 28432 22152 28441
rect 22008 28407 22060 28416
rect 22008 28373 22017 28407
rect 22017 28373 22051 28407
rect 22051 28373 22060 28407
rect 22008 28364 22060 28373
rect 23112 28568 23164 28620
rect 24216 28679 24268 28688
rect 24216 28645 24225 28679
rect 24225 28645 24259 28679
rect 24259 28645 24268 28679
rect 24216 28636 24268 28645
rect 24032 28500 24084 28552
rect 24492 28543 24544 28552
rect 24492 28509 24501 28543
rect 24501 28509 24535 28543
rect 24535 28509 24544 28543
rect 24492 28500 24544 28509
rect 22652 28432 22704 28484
rect 23388 28364 23440 28416
rect 24676 28432 24728 28484
rect 24400 28364 24452 28416
rect 8032 28262 8084 28314
rect 8096 28262 8148 28314
rect 8160 28262 8212 28314
rect 8224 28262 8276 28314
rect 8288 28262 8340 28314
rect 15115 28262 15167 28314
rect 15179 28262 15231 28314
rect 15243 28262 15295 28314
rect 15307 28262 15359 28314
rect 15371 28262 15423 28314
rect 22198 28262 22250 28314
rect 22262 28262 22314 28314
rect 22326 28262 22378 28314
rect 22390 28262 22442 28314
rect 22454 28262 22506 28314
rect 29281 28262 29333 28314
rect 29345 28262 29397 28314
rect 29409 28262 29461 28314
rect 29473 28262 29525 28314
rect 29537 28262 29589 28314
rect 3516 28160 3568 28212
rect 3608 28160 3660 28212
rect 5264 28160 5316 28212
rect 5448 28203 5500 28212
rect 5448 28169 5457 28203
rect 5457 28169 5491 28203
rect 5491 28169 5500 28203
rect 5448 28160 5500 28169
rect 6000 28203 6052 28212
rect 6000 28169 6009 28203
rect 6009 28169 6043 28203
rect 6043 28169 6052 28203
rect 6000 28160 6052 28169
rect 7012 28160 7064 28212
rect 7288 28203 7340 28212
rect 7288 28169 7297 28203
rect 7297 28169 7331 28203
rect 7331 28169 7340 28203
rect 7288 28160 7340 28169
rect 8576 28160 8628 28212
rect 4436 28092 4488 28144
rect 6184 28092 6236 28144
rect 3608 28067 3660 28076
rect 3608 28033 3617 28067
rect 3617 28033 3651 28067
rect 3651 28033 3660 28067
rect 3608 28024 3660 28033
rect 4988 27956 5040 28008
rect 5816 27931 5868 27940
rect 5816 27897 5825 27931
rect 5825 27897 5859 27931
rect 5859 27897 5868 27931
rect 5816 27888 5868 27897
rect 6460 27956 6512 28008
rect 7104 28067 7156 28076
rect 7104 28033 7113 28067
rect 7113 28033 7147 28067
rect 7147 28033 7156 28067
rect 7104 28024 7156 28033
rect 7564 28024 7616 28076
rect 9036 28024 9088 28076
rect 9404 28203 9456 28212
rect 9404 28169 9413 28203
rect 9413 28169 9447 28203
rect 9447 28169 9456 28203
rect 9404 28160 9456 28169
rect 9956 28160 10008 28212
rect 11244 28203 11296 28212
rect 11244 28169 11253 28203
rect 11253 28169 11287 28203
rect 11287 28169 11296 28203
rect 11244 28160 11296 28169
rect 9312 28024 9364 28076
rect 7472 27956 7524 28008
rect 7656 27999 7708 28008
rect 7656 27965 7665 27999
rect 7665 27965 7699 27999
rect 7699 27965 7708 27999
rect 7656 27956 7708 27965
rect 9772 27956 9824 28008
rect 11336 28024 11388 28076
rect 11980 28024 12032 28076
rect 11428 27956 11480 28008
rect 12164 28160 12216 28212
rect 7104 27888 7156 27940
rect 5080 27820 5132 27872
rect 5448 27820 5500 27872
rect 6368 27820 6420 27872
rect 6552 27820 6604 27872
rect 11336 27888 11388 27940
rect 12900 28160 12952 28212
rect 15016 28160 15068 28212
rect 16304 28160 16356 28212
rect 13084 28092 13136 28144
rect 14280 28092 14332 28144
rect 12072 27863 12124 27872
rect 12072 27829 12081 27863
rect 12081 27829 12115 27863
rect 12115 27829 12124 27863
rect 12072 27820 12124 27829
rect 12440 27820 12492 27872
rect 13452 28067 13504 28076
rect 13452 28033 13461 28067
rect 13461 28033 13495 28067
rect 13495 28033 13504 28067
rect 13452 28024 13504 28033
rect 17868 28160 17920 28212
rect 16488 28024 16540 28076
rect 15476 27956 15528 28008
rect 17684 28024 17736 28076
rect 18420 28092 18472 28144
rect 18144 28024 18196 28076
rect 18052 27956 18104 28008
rect 18328 27999 18380 28008
rect 18328 27965 18337 27999
rect 18337 27965 18371 27999
rect 18371 27965 18380 27999
rect 18328 27956 18380 27965
rect 19248 28092 19300 28144
rect 21824 28160 21876 28212
rect 22284 28160 22336 28212
rect 24216 28160 24268 28212
rect 24676 28203 24728 28212
rect 24676 28169 24685 28203
rect 24685 28169 24719 28203
rect 24719 28169 24728 28203
rect 24676 28160 24728 28169
rect 20812 28067 20864 28076
rect 20812 28033 20821 28067
rect 20821 28033 20855 28067
rect 20855 28033 20864 28067
rect 20812 28024 20864 28033
rect 22376 28024 22428 28076
rect 22652 28024 22704 28076
rect 23204 28135 23256 28144
rect 23204 28101 23213 28135
rect 23213 28101 23247 28135
rect 23247 28101 23256 28135
rect 23204 28092 23256 28101
rect 23756 28092 23808 28144
rect 14464 27820 14516 27872
rect 17132 27820 17184 27872
rect 17960 27863 18012 27872
rect 17960 27829 17969 27863
rect 17969 27829 18003 27863
rect 18003 27829 18012 27863
rect 17960 27820 18012 27829
rect 18052 27863 18104 27872
rect 18052 27829 18061 27863
rect 18061 27829 18095 27863
rect 18095 27829 18104 27863
rect 18052 27820 18104 27829
rect 19340 27956 19392 28008
rect 21272 27956 21324 28008
rect 21640 27956 21692 28008
rect 20260 27888 20312 27940
rect 22652 27931 22704 27940
rect 22652 27897 22661 27931
rect 22661 27897 22695 27931
rect 22695 27897 22704 27931
rect 22652 27888 22704 27897
rect 19892 27820 19944 27872
rect 22192 27820 22244 27872
rect 22560 27863 22612 27872
rect 22560 27829 22569 27863
rect 22569 27829 22603 27863
rect 22603 27829 22612 27863
rect 22560 27820 22612 27829
rect 4491 27718 4543 27770
rect 4555 27718 4607 27770
rect 4619 27718 4671 27770
rect 4683 27718 4735 27770
rect 4747 27718 4799 27770
rect 11574 27718 11626 27770
rect 11638 27718 11690 27770
rect 11702 27718 11754 27770
rect 11766 27718 11818 27770
rect 11830 27718 11882 27770
rect 18657 27718 18709 27770
rect 18721 27718 18773 27770
rect 18785 27718 18837 27770
rect 18849 27718 18901 27770
rect 18913 27718 18965 27770
rect 25740 27718 25792 27770
rect 25804 27718 25856 27770
rect 25868 27718 25920 27770
rect 25932 27718 25984 27770
rect 25996 27718 26048 27770
rect 3608 27616 3660 27668
rect 9312 27659 9364 27668
rect 9312 27625 9321 27659
rect 9321 27625 9355 27659
rect 9355 27625 9364 27659
rect 9312 27616 9364 27625
rect 11060 27616 11112 27668
rect 11336 27616 11388 27668
rect 7196 27548 7248 27600
rect 3148 27480 3200 27532
rect 4252 27523 4304 27532
rect 4252 27489 4261 27523
rect 4261 27489 4295 27523
rect 4295 27489 4304 27523
rect 4252 27480 4304 27489
rect 4344 27412 4396 27464
rect 1492 27387 1544 27396
rect 1492 27353 1501 27387
rect 1501 27353 1535 27387
rect 1535 27353 1544 27387
rect 1492 27344 1544 27353
rect 4160 27344 4212 27396
rect 5448 27412 5500 27464
rect 5172 27344 5224 27396
rect 7932 27387 7984 27396
rect 7932 27353 7941 27387
rect 7941 27353 7975 27387
rect 7975 27353 7984 27387
rect 7932 27344 7984 27353
rect 9772 27412 9824 27464
rect 9956 27412 10008 27464
rect 13360 27616 13412 27668
rect 14004 27616 14056 27668
rect 14464 27616 14516 27668
rect 18144 27616 18196 27668
rect 19340 27616 19392 27668
rect 22560 27616 22612 27668
rect 940 27276 992 27328
rect 2780 27276 2832 27328
rect 8576 27319 8628 27328
rect 8576 27285 8585 27319
rect 8585 27285 8619 27319
rect 8619 27285 8628 27319
rect 8576 27276 8628 27285
rect 8944 27319 8996 27328
rect 8944 27285 8953 27319
rect 8953 27285 8987 27319
rect 8987 27285 8996 27319
rect 8944 27276 8996 27285
rect 11428 27412 11480 27464
rect 11888 27412 11940 27464
rect 12072 27412 12124 27464
rect 11520 27344 11572 27396
rect 12440 27480 12492 27532
rect 22652 27548 22704 27600
rect 22836 27548 22888 27600
rect 13084 27480 13136 27532
rect 14004 27480 14056 27532
rect 15568 27480 15620 27532
rect 16488 27523 16540 27532
rect 16488 27489 16497 27523
rect 16497 27489 16531 27523
rect 16531 27489 16540 27523
rect 16488 27480 16540 27489
rect 17132 27480 17184 27532
rect 12808 27412 12860 27464
rect 10784 27276 10836 27328
rect 11888 27276 11940 27328
rect 11980 27276 12032 27328
rect 12532 27276 12584 27328
rect 14004 27276 14056 27328
rect 14464 27276 14516 27328
rect 16396 27455 16448 27464
rect 16396 27421 16405 27455
rect 16405 27421 16439 27455
rect 16439 27421 16448 27455
rect 16396 27412 16448 27421
rect 19432 27412 19484 27464
rect 19524 27455 19576 27464
rect 19524 27421 19533 27455
rect 19533 27421 19567 27455
rect 19567 27421 19576 27455
rect 20812 27480 20864 27532
rect 19524 27412 19576 27421
rect 19892 27455 19944 27464
rect 19892 27421 19901 27455
rect 19901 27421 19935 27455
rect 19935 27421 19944 27455
rect 19892 27412 19944 27421
rect 22100 27480 22152 27532
rect 22008 27455 22060 27464
rect 22008 27421 22017 27455
rect 22017 27421 22051 27455
rect 22051 27421 22060 27455
rect 22008 27412 22060 27421
rect 22284 27455 22336 27464
rect 22284 27421 22293 27455
rect 22293 27421 22327 27455
rect 22327 27421 22336 27455
rect 22284 27412 22336 27421
rect 22376 27455 22428 27464
rect 22376 27421 22385 27455
rect 22385 27421 22419 27455
rect 22419 27421 22428 27455
rect 22376 27412 22428 27421
rect 24400 27412 24452 27464
rect 17224 27344 17276 27396
rect 20076 27344 20128 27396
rect 20260 27344 20312 27396
rect 20720 27344 20772 27396
rect 22192 27344 22244 27396
rect 20996 27276 21048 27328
rect 21640 27319 21692 27328
rect 21640 27285 21649 27319
rect 21649 27285 21683 27319
rect 21683 27285 21692 27319
rect 21640 27276 21692 27285
rect 22008 27276 22060 27328
rect 8032 27174 8084 27226
rect 8096 27174 8148 27226
rect 8160 27174 8212 27226
rect 8224 27174 8276 27226
rect 8288 27174 8340 27226
rect 15115 27174 15167 27226
rect 15179 27174 15231 27226
rect 15243 27174 15295 27226
rect 15307 27174 15359 27226
rect 15371 27174 15423 27226
rect 22198 27174 22250 27226
rect 22262 27174 22314 27226
rect 22326 27174 22378 27226
rect 22390 27174 22442 27226
rect 22454 27174 22506 27226
rect 29281 27174 29333 27226
rect 29345 27174 29397 27226
rect 29409 27174 29461 27226
rect 29473 27174 29525 27226
rect 29537 27174 29589 27226
rect 8944 27072 8996 27124
rect 9772 27072 9824 27124
rect 10784 27072 10836 27124
rect 13636 27072 13688 27124
rect 14464 27072 14516 27124
rect 16396 27072 16448 27124
rect 19524 27072 19576 27124
rect 20904 27072 20956 27124
rect 22008 27072 22060 27124
rect 11152 27004 11204 27056
rect 12716 27004 12768 27056
rect 12808 27047 12860 27056
rect 12808 27013 12817 27047
rect 12817 27013 12851 27047
rect 12851 27013 12860 27047
rect 12808 27004 12860 27013
rect 14740 27004 14792 27056
rect 17132 27047 17184 27056
rect 17132 27013 17141 27047
rect 17141 27013 17175 27047
rect 17175 27013 17184 27047
rect 17132 27004 17184 27013
rect 9220 26936 9272 26988
rect 7656 26868 7708 26920
rect 8576 26868 8628 26920
rect 11520 26868 11572 26920
rect 12256 26936 12308 26988
rect 13912 26936 13964 26988
rect 11888 26911 11940 26920
rect 11888 26877 11897 26911
rect 11897 26877 11931 26911
rect 11931 26877 11940 26911
rect 11888 26868 11940 26877
rect 12440 26868 12492 26920
rect 20812 27047 20864 27056
rect 20812 27013 20821 27047
rect 20821 27013 20855 27047
rect 20855 27013 20864 27047
rect 20812 27004 20864 27013
rect 21916 26936 21968 26988
rect 28264 26936 28316 26988
rect 13912 26800 13964 26852
rect 14280 26800 14332 26852
rect 15476 26868 15528 26920
rect 18052 26800 18104 26852
rect 11244 26732 11296 26784
rect 12808 26732 12860 26784
rect 20996 26775 21048 26784
rect 20996 26741 21005 26775
rect 21005 26741 21039 26775
rect 21039 26741 21048 26775
rect 20996 26732 21048 26741
rect 29000 26775 29052 26784
rect 29000 26741 29009 26775
rect 29009 26741 29043 26775
rect 29043 26741 29052 26775
rect 29000 26732 29052 26741
rect 4491 26630 4543 26682
rect 4555 26630 4607 26682
rect 4619 26630 4671 26682
rect 4683 26630 4735 26682
rect 4747 26630 4799 26682
rect 11574 26630 11626 26682
rect 11638 26630 11690 26682
rect 11702 26630 11754 26682
rect 11766 26630 11818 26682
rect 11830 26630 11882 26682
rect 18657 26630 18709 26682
rect 18721 26630 18773 26682
rect 18785 26630 18837 26682
rect 18849 26630 18901 26682
rect 18913 26630 18965 26682
rect 25740 26630 25792 26682
rect 25804 26630 25856 26682
rect 25868 26630 25920 26682
rect 25932 26630 25984 26682
rect 25996 26630 26048 26682
rect 1492 26528 1544 26580
rect 11244 26528 11296 26580
rect 12532 26571 12584 26580
rect 12532 26537 12541 26571
rect 12541 26537 12575 26571
rect 12575 26537 12584 26571
rect 12532 26528 12584 26537
rect 2412 26367 2464 26376
rect 2412 26333 2421 26367
rect 2421 26333 2455 26367
rect 2455 26333 2464 26367
rect 2412 26324 2464 26333
rect 7012 26392 7064 26444
rect 10416 26392 10468 26444
rect 11428 26392 11480 26444
rect 12256 26392 12308 26444
rect 6276 26367 6328 26376
rect 6276 26333 6285 26367
rect 6285 26333 6319 26367
rect 6319 26333 6328 26367
rect 6276 26324 6328 26333
rect 9220 26324 9272 26376
rect 17960 26324 18012 26376
rect 11152 26256 11204 26308
rect 5816 26231 5868 26240
rect 5816 26197 5825 26231
rect 5825 26197 5859 26231
rect 5859 26197 5868 26231
rect 5816 26188 5868 26197
rect 19432 26299 19484 26308
rect 19432 26265 19441 26299
rect 19441 26265 19475 26299
rect 19475 26265 19484 26299
rect 19432 26256 19484 26265
rect 19800 26256 19852 26308
rect 8032 26086 8084 26138
rect 8096 26086 8148 26138
rect 8160 26086 8212 26138
rect 8224 26086 8276 26138
rect 8288 26086 8340 26138
rect 15115 26086 15167 26138
rect 15179 26086 15231 26138
rect 15243 26086 15295 26138
rect 15307 26086 15359 26138
rect 15371 26086 15423 26138
rect 22198 26086 22250 26138
rect 22262 26086 22314 26138
rect 22326 26086 22378 26138
rect 22390 26086 22442 26138
rect 22454 26086 22506 26138
rect 29281 26086 29333 26138
rect 29345 26086 29397 26138
rect 29409 26086 29461 26138
rect 29473 26086 29525 26138
rect 29537 26086 29589 26138
rect 7932 25984 7984 26036
rect 5816 25916 5868 25968
rect 5172 25891 5224 25900
rect 5172 25857 5181 25891
rect 5181 25857 5215 25891
rect 5215 25857 5224 25891
rect 5172 25848 5224 25857
rect 5356 25848 5408 25900
rect 6460 25916 6512 25968
rect 5540 25780 5592 25832
rect 6552 25848 6604 25900
rect 6920 25848 6972 25900
rect 7288 25891 7340 25900
rect 7288 25857 7297 25891
rect 7297 25857 7331 25891
rect 7331 25857 7340 25891
rect 7288 25848 7340 25857
rect 8576 25916 8628 25968
rect 18236 25916 18288 25968
rect 19340 25916 19392 25968
rect 20720 25984 20772 26036
rect 6736 25780 6788 25832
rect 4344 25644 4396 25696
rect 5080 25644 5132 25696
rect 5632 25687 5684 25696
rect 5632 25653 5641 25687
rect 5641 25653 5675 25687
rect 5675 25653 5684 25687
rect 5632 25644 5684 25653
rect 5724 25687 5776 25696
rect 5724 25653 5733 25687
rect 5733 25653 5767 25687
rect 5767 25653 5776 25687
rect 5724 25644 5776 25653
rect 7196 25644 7248 25696
rect 17868 25780 17920 25832
rect 7748 25712 7800 25764
rect 8760 25644 8812 25696
rect 20720 25644 20772 25696
rect 4491 25542 4543 25594
rect 4555 25542 4607 25594
rect 4619 25542 4671 25594
rect 4683 25542 4735 25594
rect 4747 25542 4799 25594
rect 11574 25542 11626 25594
rect 11638 25542 11690 25594
rect 11702 25542 11754 25594
rect 11766 25542 11818 25594
rect 11830 25542 11882 25594
rect 18657 25542 18709 25594
rect 18721 25542 18773 25594
rect 18785 25542 18837 25594
rect 18849 25542 18901 25594
rect 18913 25542 18965 25594
rect 25740 25542 25792 25594
rect 25804 25542 25856 25594
rect 25868 25542 25920 25594
rect 25932 25542 25984 25594
rect 25996 25542 26048 25594
rect 5080 25440 5132 25492
rect 5540 25440 5592 25492
rect 6460 25483 6512 25492
rect 6460 25449 6469 25483
rect 6469 25449 6503 25483
rect 6503 25449 6512 25483
rect 6460 25440 6512 25449
rect 6736 25483 6788 25492
rect 6736 25449 6745 25483
rect 6745 25449 6779 25483
rect 6779 25449 6788 25483
rect 6736 25440 6788 25449
rect 7012 25440 7064 25492
rect 7748 25440 7800 25492
rect 8760 25483 8812 25492
rect 8760 25449 8769 25483
rect 8769 25449 8803 25483
rect 8803 25449 8812 25483
rect 8760 25440 8812 25449
rect 18880 25440 18932 25492
rect 18144 25372 18196 25424
rect 4988 25304 5040 25356
rect 5356 25304 5408 25356
rect 4344 25236 4396 25288
rect 4620 25279 4672 25288
rect 4620 25245 4629 25279
rect 4629 25245 4663 25279
rect 4663 25245 4672 25279
rect 4620 25236 4672 25245
rect 3516 25168 3568 25220
rect 2780 25100 2832 25152
rect 5264 25168 5316 25220
rect 4896 25100 4948 25152
rect 5080 25100 5132 25152
rect 8392 25236 8444 25288
rect 9312 25236 9364 25288
rect 12992 25236 13044 25288
rect 13452 25236 13504 25288
rect 15016 25279 15068 25288
rect 15016 25245 15025 25279
rect 15025 25245 15059 25279
rect 15059 25245 15068 25279
rect 15016 25236 15068 25245
rect 17224 25304 17276 25356
rect 17868 25236 17920 25288
rect 19248 25304 19300 25356
rect 18880 25279 18932 25288
rect 18880 25245 18915 25279
rect 18915 25245 18932 25279
rect 18880 25236 18932 25245
rect 19064 25279 19116 25288
rect 19064 25245 19073 25279
rect 19073 25245 19107 25279
rect 19107 25245 19116 25279
rect 19064 25236 19116 25245
rect 19892 25304 19944 25356
rect 19432 25236 19484 25288
rect 19800 25236 19852 25288
rect 7288 25168 7340 25220
rect 14924 25168 14976 25220
rect 16580 25168 16632 25220
rect 5724 25100 5776 25152
rect 7472 25100 7524 25152
rect 11888 25143 11940 25152
rect 11888 25109 11897 25143
rect 11897 25109 11931 25143
rect 11931 25109 11940 25143
rect 11888 25100 11940 25109
rect 17408 25211 17460 25220
rect 17408 25177 17417 25211
rect 17417 25177 17451 25211
rect 17451 25177 17460 25211
rect 17408 25168 17460 25177
rect 17040 25143 17092 25152
rect 17040 25109 17049 25143
rect 17049 25109 17083 25143
rect 17083 25109 17092 25143
rect 17040 25100 17092 25109
rect 18420 25143 18472 25152
rect 18420 25109 18429 25143
rect 18429 25109 18463 25143
rect 18463 25109 18472 25143
rect 18420 25100 18472 25109
rect 18788 25211 18840 25220
rect 18788 25177 18797 25211
rect 18797 25177 18831 25211
rect 18831 25177 18840 25211
rect 18788 25168 18840 25177
rect 20076 25168 20128 25220
rect 21272 25304 21324 25356
rect 20812 25168 20864 25220
rect 22652 25211 22704 25220
rect 22652 25177 22661 25211
rect 22661 25177 22695 25211
rect 22695 25177 22704 25211
rect 22652 25168 22704 25177
rect 19156 25100 19208 25152
rect 8032 24998 8084 25050
rect 8096 24998 8148 25050
rect 8160 24998 8212 25050
rect 8224 24998 8276 25050
rect 8288 24998 8340 25050
rect 15115 24998 15167 25050
rect 15179 24998 15231 25050
rect 15243 24998 15295 25050
rect 15307 24998 15359 25050
rect 15371 24998 15423 25050
rect 22198 24998 22250 25050
rect 22262 24998 22314 25050
rect 22326 24998 22378 25050
rect 22390 24998 22442 25050
rect 22454 24998 22506 25050
rect 29281 24998 29333 25050
rect 29345 24998 29397 25050
rect 29409 24998 29461 25050
rect 29473 24998 29525 25050
rect 29537 24998 29589 25050
rect 5264 24896 5316 24948
rect 5448 24896 5500 24948
rect 6460 24896 6512 24948
rect 7472 24939 7524 24948
rect 7472 24905 7481 24939
rect 7481 24905 7515 24939
rect 7515 24905 7524 24939
rect 7472 24896 7524 24905
rect 14924 24939 14976 24948
rect 14924 24905 14933 24939
rect 14933 24905 14967 24939
rect 14967 24905 14976 24939
rect 14924 24896 14976 24905
rect 3516 24828 3568 24880
rect 4896 24828 4948 24880
rect 4988 24828 5040 24880
rect 3424 24735 3476 24744
rect 3424 24701 3433 24735
rect 3433 24701 3467 24735
rect 3467 24701 3476 24735
rect 3424 24692 3476 24701
rect 4620 24692 4672 24744
rect 5632 24760 5684 24812
rect 6736 24828 6788 24880
rect 11888 24828 11940 24880
rect 6552 24760 6604 24812
rect 7656 24760 7708 24812
rect 9220 24760 9272 24812
rect 9588 24760 9640 24812
rect 9680 24803 9732 24812
rect 9680 24769 9689 24803
rect 9689 24769 9723 24803
rect 9723 24769 9732 24803
rect 9680 24760 9732 24769
rect 11428 24760 11480 24812
rect 5724 24692 5776 24744
rect 6828 24692 6880 24744
rect 5264 24624 5316 24676
rect 3516 24556 3568 24608
rect 5080 24556 5132 24608
rect 6000 24624 6052 24676
rect 6920 24624 6972 24676
rect 7288 24624 7340 24676
rect 11336 24692 11388 24744
rect 14096 24828 14148 24880
rect 14832 24828 14884 24880
rect 17132 24896 17184 24948
rect 13544 24735 13596 24744
rect 13544 24701 13553 24735
rect 13553 24701 13587 24735
rect 13587 24701 13596 24735
rect 13544 24692 13596 24701
rect 14464 24735 14516 24744
rect 14464 24701 14473 24735
rect 14473 24701 14507 24735
rect 14507 24701 14516 24735
rect 14464 24692 14516 24701
rect 14556 24735 14608 24744
rect 14556 24701 14565 24735
rect 14565 24701 14599 24735
rect 14599 24701 14608 24735
rect 14556 24692 14608 24701
rect 14740 24624 14792 24676
rect 15292 24803 15344 24812
rect 15292 24769 15301 24803
rect 15301 24769 15335 24803
rect 15335 24769 15344 24803
rect 15292 24760 15344 24769
rect 15476 24760 15528 24812
rect 15660 24803 15712 24812
rect 15660 24769 15669 24803
rect 15669 24769 15703 24803
rect 15703 24769 15712 24803
rect 15660 24760 15712 24769
rect 15752 24692 15804 24744
rect 16028 24760 16080 24812
rect 17040 24828 17092 24880
rect 17040 24692 17092 24744
rect 19064 24896 19116 24948
rect 18328 24828 18380 24880
rect 18420 24828 18472 24880
rect 19340 24828 19392 24880
rect 20260 24828 20312 24880
rect 17960 24803 18012 24812
rect 17960 24769 17969 24803
rect 17969 24769 18003 24803
rect 18003 24769 18012 24803
rect 17960 24760 18012 24769
rect 18144 24803 18196 24812
rect 18144 24769 18179 24803
rect 18179 24769 18196 24803
rect 18144 24760 18196 24769
rect 7656 24599 7708 24608
rect 7656 24565 7665 24599
rect 7665 24565 7699 24599
rect 7699 24565 7708 24599
rect 7656 24556 7708 24565
rect 10416 24556 10468 24608
rect 16120 24624 16172 24676
rect 18236 24624 18288 24676
rect 20076 24692 20128 24744
rect 20720 24760 20772 24812
rect 19432 24556 19484 24608
rect 20076 24556 20128 24608
rect 4491 24454 4543 24506
rect 4555 24454 4607 24506
rect 4619 24454 4671 24506
rect 4683 24454 4735 24506
rect 4747 24454 4799 24506
rect 11574 24454 11626 24506
rect 11638 24454 11690 24506
rect 11702 24454 11754 24506
rect 11766 24454 11818 24506
rect 11830 24454 11882 24506
rect 18657 24454 18709 24506
rect 18721 24454 18773 24506
rect 18785 24454 18837 24506
rect 18849 24454 18901 24506
rect 18913 24454 18965 24506
rect 25740 24454 25792 24506
rect 25804 24454 25856 24506
rect 25868 24454 25920 24506
rect 25932 24454 25984 24506
rect 25996 24454 26048 24506
rect 3424 24352 3476 24404
rect 5356 24352 5408 24404
rect 6552 24284 6604 24336
rect 9680 24352 9732 24404
rect 15292 24352 15344 24404
rect 16028 24352 16080 24404
rect 19248 24395 19300 24404
rect 19248 24361 19257 24395
rect 19257 24361 19291 24395
rect 19291 24361 19300 24395
rect 19248 24352 19300 24361
rect 19892 24395 19944 24404
rect 19892 24361 19901 24395
rect 19901 24361 19935 24395
rect 19935 24361 19944 24395
rect 19892 24352 19944 24361
rect 7472 24284 7524 24336
rect 14464 24284 14516 24336
rect 19432 24284 19484 24336
rect 4988 24216 5040 24268
rect 6828 24216 6880 24268
rect 15016 24216 15068 24268
rect 7012 24148 7064 24200
rect 7196 24148 7248 24200
rect 10048 24191 10100 24200
rect 10048 24157 10057 24191
rect 10057 24157 10091 24191
rect 10091 24157 10100 24191
rect 10048 24148 10100 24157
rect 6000 24080 6052 24132
rect 9496 24012 9548 24064
rect 9680 24012 9732 24064
rect 11888 24123 11940 24132
rect 11888 24089 11897 24123
rect 11897 24089 11931 24123
rect 11931 24089 11940 24123
rect 11888 24080 11940 24089
rect 13452 24080 13504 24132
rect 13912 24148 13964 24200
rect 15936 24216 15988 24268
rect 16120 24216 16172 24268
rect 16396 24259 16448 24268
rect 16396 24225 16405 24259
rect 16405 24225 16439 24259
rect 16439 24225 16448 24259
rect 16396 24216 16448 24225
rect 16304 24191 16356 24200
rect 16304 24157 16313 24191
rect 16313 24157 16347 24191
rect 16347 24157 16356 24191
rect 16304 24148 16356 24157
rect 17960 24148 18012 24200
rect 19064 24148 19116 24200
rect 15016 24080 15068 24132
rect 15936 24123 15988 24132
rect 15936 24089 15945 24123
rect 15945 24089 15979 24123
rect 15979 24089 15988 24123
rect 15936 24080 15988 24089
rect 16028 24123 16080 24132
rect 16028 24089 16037 24123
rect 16037 24089 16071 24123
rect 16071 24089 16080 24123
rect 16028 24080 16080 24089
rect 16212 24080 16264 24132
rect 14372 24012 14424 24064
rect 17224 24080 17276 24132
rect 18052 24080 18104 24132
rect 19892 24080 19944 24132
rect 20076 24191 20128 24200
rect 20076 24157 20085 24191
rect 20085 24157 20119 24191
rect 20119 24157 20128 24191
rect 20076 24148 20128 24157
rect 20260 24080 20312 24132
rect 20076 24012 20128 24064
rect 8032 23910 8084 23962
rect 8096 23910 8148 23962
rect 8160 23910 8212 23962
rect 8224 23910 8276 23962
rect 8288 23910 8340 23962
rect 15115 23910 15167 23962
rect 15179 23910 15231 23962
rect 15243 23910 15295 23962
rect 15307 23910 15359 23962
rect 15371 23910 15423 23962
rect 22198 23910 22250 23962
rect 22262 23910 22314 23962
rect 22326 23910 22378 23962
rect 22390 23910 22442 23962
rect 22454 23910 22506 23962
rect 29281 23910 29333 23962
rect 29345 23910 29397 23962
rect 29409 23910 29461 23962
rect 29473 23910 29525 23962
rect 29537 23910 29589 23962
rect 5172 23808 5224 23860
rect 7656 23808 7708 23860
rect 11888 23808 11940 23860
rect 12992 23851 13044 23860
rect 12992 23817 13001 23851
rect 13001 23817 13035 23851
rect 13035 23817 13044 23851
rect 12992 23808 13044 23817
rect 5724 23740 5776 23792
rect 9496 23740 9548 23792
rect 10784 23740 10836 23792
rect 11336 23740 11388 23792
rect 14832 23808 14884 23860
rect 15936 23808 15988 23860
rect 1492 23715 1544 23724
rect 1492 23681 1501 23715
rect 1501 23681 1535 23715
rect 1535 23681 1544 23715
rect 1492 23672 1544 23681
rect 12808 23672 12860 23724
rect 1584 23511 1636 23520
rect 1584 23477 1593 23511
rect 1593 23477 1627 23511
rect 1627 23477 1636 23511
rect 1584 23468 1636 23477
rect 9312 23468 9364 23520
rect 10784 23468 10836 23520
rect 15660 23783 15712 23792
rect 15660 23749 15669 23783
rect 15669 23749 15703 23783
rect 15703 23749 15712 23783
rect 15660 23740 15712 23749
rect 16028 23740 16080 23792
rect 16304 23740 16356 23792
rect 17500 23740 17552 23792
rect 12164 23511 12216 23520
rect 12164 23477 12173 23511
rect 12173 23477 12207 23511
rect 12207 23477 12216 23511
rect 12164 23468 12216 23477
rect 13544 23647 13596 23656
rect 13544 23613 13553 23647
rect 13553 23613 13587 23647
rect 13587 23613 13596 23647
rect 13544 23604 13596 23613
rect 14372 23604 14424 23656
rect 15384 23672 15436 23724
rect 15200 23604 15252 23656
rect 15200 23468 15252 23520
rect 15568 23715 15620 23724
rect 15568 23681 15577 23715
rect 15577 23681 15611 23715
rect 15611 23681 15620 23715
rect 15568 23672 15620 23681
rect 16120 23672 16172 23724
rect 15476 23536 15528 23588
rect 15752 23536 15804 23588
rect 15936 23579 15988 23588
rect 15936 23545 15945 23579
rect 15945 23545 15979 23579
rect 15979 23545 15988 23579
rect 15936 23536 15988 23545
rect 16212 23468 16264 23520
rect 17040 23672 17092 23724
rect 17132 23715 17184 23724
rect 17132 23681 17141 23715
rect 17141 23681 17175 23715
rect 17175 23681 17184 23715
rect 17132 23672 17184 23681
rect 19892 23808 19944 23860
rect 22652 23808 22704 23860
rect 17132 23536 17184 23588
rect 17960 23647 18012 23656
rect 17960 23613 17969 23647
rect 17969 23613 18003 23647
rect 18003 23613 18012 23647
rect 17960 23604 18012 23613
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 4491 23366 4543 23418
rect 4555 23366 4607 23418
rect 4619 23366 4671 23418
rect 4683 23366 4735 23418
rect 4747 23366 4799 23418
rect 11574 23366 11626 23418
rect 11638 23366 11690 23418
rect 11702 23366 11754 23418
rect 11766 23366 11818 23418
rect 11830 23366 11882 23418
rect 18657 23366 18709 23418
rect 18721 23366 18773 23418
rect 18785 23366 18837 23418
rect 18849 23366 18901 23418
rect 18913 23366 18965 23418
rect 25740 23366 25792 23418
rect 25804 23366 25856 23418
rect 25868 23366 25920 23418
rect 25932 23366 25984 23418
rect 25996 23366 26048 23418
rect 10048 23264 10100 23316
rect 10508 23264 10560 23316
rect 14556 23264 14608 23316
rect 14924 23307 14976 23316
rect 14924 23273 14933 23307
rect 14933 23273 14967 23307
rect 14967 23273 14976 23307
rect 14924 23264 14976 23273
rect 15016 23264 15068 23316
rect 16396 23264 16448 23316
rect 17408 23264 17460 23316
rect 25228 23307 25280 23316
rect 25228 23273 25237 23307
rect 25237 23273 25271 23307
rect 25271 23273 25280 23307
rect 25228 23264 25280 23273
rect 6828 23171 6880 23180
rect 6828 23137 6837 23171
rect 6837 23137 6871 23171
rect 6871 23137 6880 23171
rect 6828 23128 6880 23137
rect 9312 23128 9364 23180
rect 11428 23128 11480 23180
rect 6184 23060 6236 23112
rect 10692 23060 10744 23112
rect 10876 23103 10928 23112
rect 10876 23069 10885 23103
rect 10885 23069 10919 23103
rect 10919 23069 10928 23103
rect 15200 23239 15252 23248
rect 15200 23205 15209 23239
rect 15209 23205 15243 23239
rect 15243 23205 15252 23239
rect 15200 23196 15252 23205
rect 15568 23239 15620 23248
rect 15568 23205 15577 23239
rect 15577 23205 15611 23239
rect 15611 23205 15620 23239
rect 15568 23196 15620 23205
rect 15936 23196 15988 23248
rect 18144 23196 18196 23248
rect 14556 23128 14608 23180
rect 10876 23060 10928 23069
rect 13544 23060 13596 23112
rect 14004 23060 14056 23112
rect 14740 23103 14792 23112
rect 14740 23069 14749 23103
rect 14749 23069 14783 23103
rect 14783 23069 14792 23103
rect 14740 23060 14792 23069
rect 5080 22967 5132 22976
rect 5080 22933 5089 22967
rect 5089 22933 5123 22967
rect 5123 22933 5132 22967
rect 5080 22924 5132 22933
rect 5264 22924 5316 22976
rect 9220 22992 9272 23044
rect 13912 22992 13964 23044
rect 15384 23060 15436 23112
rect 16028 23171 16080 23180
rect 16028 23137 16037 23171
rect 16037 23137 16071 23171
rect 16071 23137 16080 23171
rect 16028 23128 16080 23137
rect 21640 23128 21692 23180
rect 24308 23128 24360 23180
rect 25044 23128 25096 23180
rect 15476 23035 15528 23044
rect 14280 22967 14332 22976
rect 14280 22933 14289 22967
rect 14289 22933 14323 22967
rect 14323 22933 14332 22967
rect 14280 22924 14332 22933
rect 14372 22924 14424 22976
rect 15476 23001 15485 23035
rect 15485 23001 15519 23035
rect 15519 23001 15528 23035
rect 15476 22992 15528 23001
rect 15568 22992 15620 23044
rect 14924 22924 14976 22976
rect 15108 22924 15160 22976
rect 16764 22992 16816 23044
rect 18328 23060 18380 23112
rect 20720 23103 20772 23112
rect 20720 23069 20729 23103
rect 20729 23069 20763 23103
rect 20763 23069 20772 23103
rect 20720 23060 20772 23069
rect 20812 23103 20864 23112
rect 20812 23069 20821 23103
rect 20821 23069 20855 23103
rect 20855 23069 20864 23103
rect 20812 23060 20864 23069
rect 21732 23060 21784 23112
rect 24492 23103 24544 23112
rect 24492 23069 24501 23103
rect 24501 23069 24535 23103
rect 24535 23069 24544 23103
rect 24492 23060 24544 23069
rect 21180 23035 21232 23044
rect 21180 23001 21189 23035
rect 21189 23001 21223 23035
rect 21223 23001 21232 23035
rect 21180 22992 21232 23001
rect 22560 22992 22612 23044
rect 24676 22992 24728 23044
rect 16212 22924 16264 22976
rect 17592 22924 17644 22976
rect 18052 22924 18104 22976
rect 20996 22967 21048 22976
rect 20996 22933 21005 22967
rect 21005 22933 21039 22967
rect 21039 22933 21048 22967
rect 20996 22924 21048 22933
rect 23480 22924 23532 22976
rect 24124 22924 24176 22976
rect 24768 22924 24820 22976
rect 24952 22924 25004 22976
rect 25504 22992 25556 23044
rect 8032 22822 8084 22874
rect 8096 22822 8148 22874
rect 8160 22822 8212 22874
rect 8224 22822 8276 22874
rect 8288 22822 8340 22874
rect 15115 22822 15167 22874
rect 15179 22822 15231 22874
rect 15243 22822 15295 22874
rect 15307 22822 15359 22874
rect 15371 22822 15423 22874
rect 22198 22822 22250 22874
rect 22262 22822 22314 22874
rect 22326 22822 22378 22874
rect 22390 22822 22442 22874
rect 22454 22822 22506 22874
rect 29281 22822 29333 22874
rect 29345 22822 29397 22874
rect 29409 22822 29461 22874
rect 29473 22822 29525 22874
rect 29537 22822 29589 22874
rect 6920 22720 6972 22772
rect 10232 22720 10284 22772
rect 5264 22695 5316 22704
rect 5264 22661 5273 22695
rect 5273 22661 5307 22695
rect 5307 22661 5316 22695
rect 5264 22652 5316 22661
rect 9680 22652 9732 22704
rect 12808 22763 12860 22772
rect 12808 22729 12817 22763
rect 12817 22729 12851 22763
rect 12851 22729 12860 22763
rect 12808 22720 12860 22729
rect 15016 22720 15068 22772
rect 12532 22695 12584 22704
rect 12532 22661 12541 22695
rect 12541 22661 12575 22695
rect 12575 22661 12584 22695
rect 12532 22652 12584 22661
rect 20720 22720 20772 22772
rect 5632 22516 5684 22568
rect 6000 22559 6052 22568
rect 6000 22525 6009 22559
rect 6009 22525 6043 22559
rect 6043 22525 6052 22559
rect 6000 22516 6052 22525
rect 4160 22380 4212 22432
rect 8116 22584 8168 22636
rect 8668 22627 8720 22636
rect 8668 22593 8677 22627
rect 8677 22593 8711 22627
rect 8711 22593 8720 22627
rect 8668 22584 8720 22593
rect 8852 22627 8904 22636
rect 8852 22593 8861 22627
rect 8861 22593 8895 22627
rect 8895 22593 8904 22627
rect 8852 22584 8904 22593
rect 7656 22559 7708 22568
rect 7656 22525 7665 22559
rect 7665 22525 7699 22559
rect 7699 22525 7708 22559
rect 7656 22516 7708 22525
rect 9312 22627 9364 22636
rect 9312 22593 9321 22627
rect 9321 22593 9355 22627
rect 9355 22593 9364 22627
rect 9312 22584 9364 22593
rect 10968 22584 11020 22636
rect 12164 22584 12216 22636
rect 12624 22627 12676 22636
rect 12624 22593 12633 22627
rect 12633 22593 12667 22627
rect 12667 22593 12676 22627
rect 12624 22584 12676 22593
rect 9220 22491 9272 22500
rect 9220 22457 9229 22491
rect 9229 22457 9263 22491
rect 9263 22457 9272 22491
rect 9220 22448 9272 22457
rect 9956 22516 10008 22568
rect 11428 22516 11480 22568
rect 13912 22448 13964 22500
rect 20720 22627 20772 22636
rect 20720 22593 20729 22627
rect 20729 22593 20763 22627
rect 20763 22593 20772 22627
rect 20720 22584 20772 22593
rect 20812 22584 20864 22636
rect 23480 22720 23532 22772
rect 21732 22652 21784 22704
rect 21640 22584 21692 22636
rect 22836 22652 22888 22704
rect 15660 22516 15712 22568
rect 16488 22516 16540 22568
rect 16672 22559 16724 22568
rect 16672 22525 16681 22559
rect 16681 22525 16715 22559
rect 16715 22525 16724 22559
rect 16672 22516 16724 22525
rect 20444 22516 20496 22568
rect 21364 22559 21416 22568
rect 21364 22525 21373 22559
rect 21373 22525 21407 22559
rect 21407 22525 21416 22559
rect 21364 22516 21416 22525
rect 23020 22584 23072 22636
rect 23296 22627 23348 22636
rect 23296 22593 23305 22627
rect 23305 22593 23339 22627
rect 23339 22593 23348 22627
rect 23296 22584 23348 22593
rect 23572 22584 23624 22636
rect 25320 22720 25372 22772
rect 6920 22380 6972 22432
rect 7288 22423 7340 22432
rect 7288 22389 7297 22423
rect 7297 22389 7331 22423
rect 7331 22389 7340 22423
rect 7288 22380 7340 22389
rect 7748 22380 7800 22432
rect 9404 22380 9456 22432
rect 10232 22380 10284 22432
rect 14832 22423 14884 22432
rect 14832 22389 14841 22423
rect 14841 22389 14875 22423
rect 14875 22389 14884 22423
rect 14832 22380 14884 22389
rect 15936 22448 15988 22500
rect 21180 22448 21232 22500
rect 21456 22448 21508 22500
rect 23388 22516 23440 22568
rect 21640 22448 21692 22500
rect 24124 22627 24176 22636
rect 24124 22593 24133 22627
rect 24133 22593 24167 22627
rect 24167 22593 24176 22627
rect 24124 22584 24176 22593
rect 24308 22627 24360 22636
rect 24308 22593 24317 22627
rect 24317 22593 24351 22627
rect 24351 22593 24360 22627
rect 24308 22584 24360 22593
rect 24400 22584 24452 22636
rect 24584 22627 24636 22636
rect 24584 22593 24593 22627
rect 24593 22593 24627 22627
rect 24627 22593 24636 22627
rect 24584 22584 24636 22593
rect 24952 22652 25004 22704
rect 24860 22627 24912 22636
rect 24860 22593 24869 22627
rect 24869 22593 24903 22627
rect 24903 22593 24912 22627
rect 24860 22584 24912 22593
rect 25044 22627 25096 22636
rect 25044 22593 25053 22627
rect 25053 22593 25087 22627
rect 25087 22593 25096 22627
rect 25044 22584 25096 22593
rect 25228 22627 25280 22636
rect 25228 22593 25237 22627
rect 25237 22593 25271 22627
rect 25271 22593 25280 22627
rect 25228 22584 25280 22593
rect 28816 22627 28868 22636
rect 28816 22593 28825 22627
rect 28825 22593 28859 22627
rect 28859 22593 28868 22627
rect 28816 22584 28868 22593
rect 24216 22516 24268 22568
rect 24032 22448 24084 22500
rect 15568 22380 15620 22432
rect 15844 22380 15896 22432
rect 21088 22423 21140 22432
rect 21088 22389 21097 22423
rect 21097 22389 21131 22423
rect 21131 22389 21140 22423
rect 21088 22380 21140 22389
rect 21548 22380 21600 22432
rect 22100 22380 22152 22432
rect 22744 22423 22796 22432
rect 22744 22389 22753 22423
rect 22753 22389 22787 22423
rect 22787 22389 22796 22423
rect 22744 22380 22796 22389
rect 22836 22380 22888 22432
rect 23204 22380 23256 22432
rect 24952 22448 25004 22500
rect 25596 22516 25648 22568
rect 29000 22491 29052 22500
rect 29000 22457 29009 22491
rect 29009 22457 29043 22491
rect 29043 22457 29052 22491
rect 29000 22448 29052 22457
rect 4491 22278 4543 22330
rect 4555 22278 4607 22330
rect 4619 22278 4671 22330
rect 4683 22278 4735 22330
rect 4747 22278 4799 22330
rect 11574 22278 11626 22330
rect 11638 22278 11690 22330
rect 11702 22278 11754 22330
rect 11766 22278 11818 22330
rect 11830 22278 11882 22330
rect 18657 22278 18709 22330
rect 18721 22278 18773 22330
rect 18785 22278 18837 22330
rect 18849 22278 18901 22330
rect 18913 22278 18965 22330
rect 25740 22278 25792 22330
rect 25804 22278 25856 22330
rect 25868 22278 25920 22330
rect 25932 22278 25984 22330
rect 25996 22278 26048 22330
rect 7288 22176 7340 22228
rect 7656 22176 7708 22228
rect 8668 22176 8720 22228
rect 8116 22108 8168 22160
rect 10600 22176 10652 22228
rect 11152 22176 11204 22228
rect 12624 22176 12676 22228
rect 14832 22176 14884 22228
rect 6000 22083 6052 22092
rect 6000 22049 6009 22083
rect 6009 22049 6043 22083
rect 6043 22049 6052 22083
rect 6000 22040 6052 22049
rect 6368 22040 6420 22092
rect 7288 22040 7340 22092
rect 4252 22015 4304 22024
rect 4252 21981 4261 22015
rect 4261 21981 4295 22015
rect 4295 21981 4304 22015
rect 4252 21972 4304 21981
rect 4436 21904 4488 21956
rect 5356 22015 5408 22024
rect 5356 21981 5365 22015
rect 5365 21981 5399 22015
rect 5399 21981 5408 22015
rect 5356 21972 5408 21981
rect 5448 21972 5500 22024
rect 5908 22015 5960 22024
rect 5908 21981 5917 22015
rect 5917 21981 5951 22015
rect 5951 21981 5960 22015
rect 5908 21972 5960 21981
rect 3332 21836 3384 21888
rect 4068 21879 4120 21888
rect 4068 21845 4077 21879
rect 4077 21845 4111 21879
rect 4111 21845 4120 21879
rect 4068 21836 4120 21845
rect 4528 21836 4580 21888
rect 5172 21836 5224 21888
rect 9404 22015 9456 22024
rect 9404 21981 9413 22015
rect 9413 21981 9447 22015
rect 9447 21981 9456 22015
rect 9404 21972 9456 21981
rect 8392 21904 8444 21956
rect 8852 21904 8904 21956
rect 9496 21904 9548 21956
rect 7104 21836 7156 21888
rect 7840 21836 7892 21888
rect 8484 21879 8536 21888
rect 8484 21845 8493 21879
rect 8493 21845 8527 21879
rect 8527 21845 8536 21879
rect 8484 21836 8536 21845
rect 8576 21836 8628 21888
rect 9404 21836 9456 21888
rect 9956 22040 10008 22092
rect 12532 22108 12584 22160
rect 20352 22151 20404 22160
rect 20352 22117 20361 22151
rect 20361 22117 20395 22151
rect 20395 22117 20404 22151
rect 20352 22108 20404 22117
rect 21364 22176 21416 22228
rect 21640 22219 21692 22228
rect 21640 22185 21649 22219
rect 21649 22185 21683 22219
rect 21683 22185 21692 22219
rect 21640 22176 21692 22185
rect 21732 22176 21784 22228
rect 10232 21904 10284 21956
rect 10508 22015 10560 22024
rect 10508 21981 10518 22015
rect 10518 21981 10552 22015
rect 10552 21981 10560 22015
rect 10508 21972 10560 21981
rect 14464 22083 14516 22092
rect 14464 22049 14473 22083
rect 14473 22049 14507 22083
rect 14507 22049 14516 22083
rect 14464 22040 14516 22049
rect 16488 22040 16540 22092
rect 18052 22040 18104 22092
rect 19248 22040 19300 22092
rect 21272 22108 21324 22160
rect 22560 22176 22612 22228
rect 24216 22176 24268 22228
rect 24676 22176 24728 22228
rect 24768 22219 24820 22228
rect 24768 22185 24777 22219
rect 24777 22185 24811 22219
rect 24811 22185 24820 22219
rect 24768 22176 24820 22185
rect 10784 22015 10836 22024
rect 10784 21981 10793 22015
rect 10793 21981 10827 22015
rect 10827 21981 10836 22015
rect 10784 21972 10836 21981
rect 11980 21972 12032 22024
rect 17224 21972 17276 22024
rect 18420 21972 18472 22024
rect 10600 21904 10652 21956
rect 10692 21947 10744 21956
rect 10692 21913 10701 21947
rect 10701 21913 10735 21947
rect 10735 21913 10744 21947
rect 10692 21904 10744 21913
rect 10508 21836 10560 21888
rect 10968 21836 11020 21888
rect 12072 21836 12124 21888
rect 12624 21904 12676 21956
rect 13360 21904 13412 21956
rect 20444 21972 20496 22024
rect 20720 21972 20772 22024
rect 20812 22015 20864 22024
rect 20812 21981 20821 22015
rect 20821 21981 20855 22015
rect 20855 21981 20864 22015
rect 20812 21972 20864 21981
rect 20996 21972 21048 22024
rect 21088 22015 21140 22024
rect 21088 21981 21097 22015
rect 21097 21981 21131 22015
rect 21131 21981 21140 22015
rect 21088 21972 21140 21981
rect 21456 22015 21508 22024
rect 21456 21981 21465 22015
rect 21465 21981 21499 22015
rect 21499 21981 21508 22015
rect 21456 21972 21508 21981
rect 21548 21972 21600 22024
rect 23848 22108 23900 22160
rect 24308 22108 24360 22160
rect 22560 22083 22612 22092
rect 22560 22049 22569 22083
rect 22569 22049 22603 22083
rect 22603 22049 22612 22083
rect 22560 22040 22612 22049
rect 22100 21972 22152 22024
rect 23388 22083 23440 22092
rect 23388 22049 23397 22083
rect 23397 22049 23431 22083
rect 23431 22049 23440 22083
rect 23388 22040 23440 22049
rect 23572 22040 23624 22092
rect 21640 21904 21692 21956
rect 12900 21836 12952 21888
rect 13636 21836 13688 21888
rect 16304 21836 16356 21888
rect 16672 21836 16724 21888
rect 17868 21879 17920 21888
rect 17868 21845 17877 21879
rect 17877 21845 17911 21879
rect 17911 21845 17920 21879
rect 17868 21836 17920 21845
rect 20444 21836 20496 21888
rect 22560 21836 22612 21888
rect 22928 21947 22980 21956
rect 22928 21913 22937 21947
rect 22937 21913 22971 21947
rect 22971 21913 22980 21947
rect 22928 21904 22980 21913
rect 23204 22015 23256 22024
rect 23204 21981 23222 22015
rect 23222 21981 23256 22015
rect 23204 21972 23256 21981
rect 24492 21972 24544 22024
rect 24676 21972 24728 22024
rect 25228 22040 25280 22092
rect 25044 21972 25096 22024
rect 25136 22015 25188 22024
rect 25136 21981 25145 22015
rect 25145 21981 25179 22015
rect 25179 21981 25188 22015
rect 25136 21972 25188 21981
rect 25504 21972 25556 22024
rect 23296 21836 23348 21888
rect 24216 21836 24268 21888
rect 24400 21879 24452 21888
rect 24400 21845 24409 21879
rect 24409 21845 24443 21879
rect 24443 21845 24452 21879
rect 24400 21836 24452 21845
rect 28816 21972 28868 22024
rect 25596 21836 25648 21888
rect 25688 21836 25740 21888
rect 8032 21734 8084 21786
rect 8096 21734 8148 21786
rect 8160 21734 8212 21786
rect 8224 21734 8276 21786
rect 8288 21734 8340 21786
rect 15115 21734 15167 21786
rect 15179 21734 15231 21786
rect 15243 21734 15295 21786
rect 15307 21734 15359 21786
rect 15371 21734 15423 21786
rect 22198 21734 22250 21786
rect 22262 21734 22314 21786
rect 22326 21734 22378 21786
rect 22390 21734 22442 21786
rect 22454 21734 22506 21786
rect 29281 21734 29333 21786
rect 29345 21734 29397 21786
rect 29409 21734 29461 21786
rect 29473 21734 29525 21786
rect 29537 21734 29589 21786
rect 4160 21632 4212 21684
rect 4436 21632 4488 21684
rect 5356 21632 5408 21684
rect 5908 21632 5960 21684
rect 6184 21675 6236 21684
rect 6184 21641 6193 21675
rect 6193 21641 6227 21675
rect 6227 21641 6236 21675
rect 6184 21632 6236 21641
rect 3332 21607 3384 21616
rect 3332 21573 3341 21607
rect 3341 21573 3375 21607
rect 3375 21573 3384 21607
rect 3332 21564 3384 21573
rect 3424 21539 3476 21548
rect 3424 21505 3433 21539
rect 3433 21505 3467 21539
rect 3467 21505 3476 21539
rect 3424 21496 3476 21505
rect 4528 21564 4580 21616
rect 5080 21428 5132 21480
rect 5816 21539 5868 21548
rect 5816 21505 5825 21539
rect 5825 21505 5859 21539
rect 5859 21505 5868 21539
rect 5816 21496 5868 21505
rect 6000 21539 6052 21548
rect 6000 21505 6009 21539
rect 6009 21505 6043 21539
rect 6043 21505 6052 21539
rect 6000 21496 6052 21505
rect 7932 21632 7984 21684
rect 7104 21564 7156 21616
rect 8392 21607 8444 21616
rect 8392 21573 8401 21607
rect 8401 21573 8435 21607
rect 8435 21573 8444 21607
rect 8392 21564 8444 21573
rect 8484 21607 8536 21616
rect 8484 21573 8493 21607
rect 8493 21573 8527 21607
rect 8527 21573 8536 21607
rect 8484 21564 8536 21573
rect 8208 21539 8260 21548
rect 8208 21505 8217 21539
rect 8217 21505 8251 21539
rect 8251 21505 8260 21539
rect 8208 21496 8260 21505
rect 8576 21539 8628 21548
rect 8576 21505 8585 21539
rect 8585 21505 8619 21539
rect 8619 21505 8628 21539
rect 8576 21496 8628 21505
rect 9956 21632 10008 21684
rect 10968 21564 11020 21616
rect 12072 21539 12124 21548
rect 12072 21505 12081 21539
rect 12081 21505 12115 21539
rect 12115 21505 12124 21539
rect 12072 21496 12124 21505
rect 12164 21539 12216 21548
rect 12164 21505 12174 21539
rect 12174 21505 12208 21539
rect 12208 21505 12216 21539
rect 12164 21496 12216 21505
rect 3700 21335 3752 21344
rect 3700 21301 3709 21335
rect 3709 21301 3743 21335
rect 3743 21301 3752 21335
rect 3700 21292 3752 21301
rect 3792 21292 3844 21344
rect 4068 21292 4120 21344
rect 5724 21428 5776 21480
rect 7748 21360 7800 21412
rect 8208 21360 8260 21412
rect 10324 21428 10376 21480
rect 12624 21496 12676 21548
rect 12716 21428 12768 21480
rect 6460 21292 6512 21344
rect 7380 21292 7432 21344
rect 7840 21292 7892 21344
rect 10784 21335 10836 21344
rect 10784 21301 10793 21335
rect 10793 21301 10827 21335
rect 10827 21301 10836 21335
rect 10784 21292 10836 21301
rect 12624 21292 12676 21344
rect 14464 21632 14516 21684
rect 18420 21675 18472 21684
rect 18420 21641 18429 21675
rect 18429 21641 18463 21675
rect 18463 21641 18472 21675
rect 18420 21632 18472 21641
rect 13636 21564 13688 21616
rect 17224 21564 17276 21616
rect 19616 21564 19668 21616
rect 13268 21428 13320 21480
rect 16580 21428 16632 21480
rect 16948 21471 17000 21480
rect 16948 21437 16957 21471
rect 16957 21437 16991 21471
rect 16991 21437 17000 21471
rect 16948 21428 17000 21437
rect 19064 21496 19116 21548
rect 19156 21539 19208 21548
rect 19156 21505 19165 21539
rect 19165 21505 19199 21539
rect 19199 21505 19208 21539
rect 19156 21496 19208 21505
rect 19432 21496 19484 21548
rect 20812 21675 20864 21684
rect 20812 21641 20821 21675
rect 20821 21641 20855 21675
rect 20855 21641 20864 21675
rect 20812 21632 20864 21641
rect 21456 21632 21508 21684
rect 21640 21632 21692 21684
rect 21364 21564 21416 21616
rect 12992 21292 13044 21344
rect 14740 21292 14792 21344
rect 19708 21428 19760 21480
rect 20628 21471 20680 21480
rect 20628 21437 20637 21471
rect 20637 21437 20671 21471
rect 20671 21437 20680 21471
rect 20628 21428 20680 21437
rect 21272 21471 21324 21480
rect 21272 21437 21281 21471
rect 21281 21437 21315 21471
rect 21315 21437 21324 21471
rect 21272 21428 21324 21437
rect 21364 21471 21416 21480
rect 21364 21437 21373 21471
rect 21373 21437 21407 21471
rect 21407 21437 21416 21471
rect 21364 21428 21416 21437
rect 20720 21360 20772 21412
rect 19524 21335 19576 21344
rect 19524 21301 19533 21335
rect 19533 21301 19567 21335
rect 19567 21301 19576 21335
rect 19524 21292 19576 21301
rect 20628 21292 20680 21344
rect 21364 21292 21416 21344
rect 22008 21539 22060 21548
rect 22008 21505 22017 21539
rect 22017 21505 22051 21539
rect 22051 21505 22060 21539
rect 22008 21496 22060 21505
rect 23296 21632 23348 21684
rect 23480 21632 23532 21684
rect 24124 21632 24176 21684
rect 22560 21564 22612 21616
rect 22836 21573 22888 21616
rect 22836 21564 22845 21573
rect 22845 21564 22879 21573
rect 22879 21564 22888 21573
rect 24032 21564 24084 21616
rect 24860 21564 24912 21616
rect 25136 21564 25188 21616
rect 24400 21496 24452 21548
rect 24676 21539 24728 21548
rect 24676 21505 24685 21539
rect 24685 21505 24719 21539
rect 24719 21505 24728 21539
rect 24676 21496 24728 21505
rect 24952 21539 25004 21548
rect 24952 21505 24961 21539
rect 24961 21505 24995 21539
rect 24995 21505 25004 21539
rect 24952 21496 25004 21505
rect 25320 21539 25372 21548
rect 25320 21505 25329 21539
rect 25329 21505 25363 21539
rect 25363 21505 25372 21539
rect 25320 21496 25372 21505
rect 25504 21539 25556 21548
rect 25504 21505 25513 21539
rect 25513 21505 25547 21539
rect 25547 21505 25556 21539
rect 25504 21496 25556 21505
rect 26976 21539 27028 21548
rect 26976 21505 26985 21539
rect 26985 21505 27019 21539
rect 27019 21505 27028 21539
rect 26976 21496 27028 21505
rect 27528 21539 27580 21548
rect 22560 21471 22612 21480
rect 22560 21437 22569 21471
rect 22569 21437 22603 21471
rect 22603 21437 22612 21471
rect 22560 21428 22612 21437
rect 21824 21403 21876 21412
rect 21824 21369 21833 21403
rect 21833 21369 21867 21403
rect 21867 21369 21876 21403
rect 21824 21360 21876 21369
rect 22928 21471 22980 21480
rect 22928 21437 22937 21471
rect 22937 21437 22971 21471
rect 22971 21437 22980 21471
rect 22928 21428 22980 21437
rect 23388 21428 23440 21480
rect 23480 21471 23532 21480
rect 23480 21437 23489 21471
rect 23489 21437 23523 21471
rect 23523 21437 23532 21471
rect 23480 21428 23532 21437
rect 27528 21505 27537 21539
rect 27537 21505 27571 21539
rect 27571 21505 27580 21539
rect 27528 21496 27580 21505
rect 27804 21496 27856 21548
rect 22836 21360 22888 21412
rect 23204 21403 23256 21412
rect 23204 21369 23213 21403
rect 23213 21369 23247 21403
rect 23247 21369 23256 21403
rect 23204 21360 23256 21369
rect 26240 21360 26292 21412
rect 27068 21403 27120 21412
rect 27068 21369 27077 21403
rect 27077 21369 27111 21403
rect 27111 21369 27120 21403
rect 27068 21360 27120 21369
rect 22652 21292 22704 21344
rect 23848 21335 23900 21344
rect 23848 21301 23857 21335
rect 23857 21301 23891 21335
rect 23891 21301 23900 21335
rect 23848 21292 23900 21301
rect 24584 21292 24636 21344
rect 27252 21292 27304 21344
rect 27620 21335 27672 21344
rect 27620 21301 27629 21335
rect 27629 21301 27663 21335
rect 27663 21301 27672 21335
rect 27620 21292 27672 21301
rect 4491 21190 4543 21242
rect 4555 21190 4607 21242
rect 4619 21190 4671 21242
rect 4683 21190 4735 21242
rect 4747 21190 4799 21242
rect 11574 21190 11626 21242
rect 11638 21190 11690 21242
rect 11702 21190 11754 21242
rect 11766 21190 11818 21242
rect 11830 21190 11882 21242
rect 18657 21190 18709 21242
rect 18721 21190 18773 21242
rect 18785 21190 18837 21242
rect 18849 21190 18901 21242
rect 18913 21190 18965 21242
rect 25740 21190 25792 21242
rect 25804 21190 25856 21242
rect 25868 21190 25920 21242
rect 25932 21190 25984 21242
rect 25996 21190 26048 21242
rect 3700 21088 3752 21140
rect 5632 21088 5684 21140
rect 3792 20995 3844 21004
rect 3792 20961 3801 20995
rect 3801 20961 3835 20995
rect 3835 20961 3844 20995
rect 6368 21088 6420 21140
rect 10692 21088 10744 21140
rect 3792 20952 3844 20961
rect 1860 20884 1912 20936
rect 5356 20884 5408 20936
rect 5816 20884 5868 20936
rect 6184 20884 6236 20936
rect 6736 20884 6788 20936
rect 7012 20884 7064 20936
rect 7380 20927 7432 20936
rect 7380 20893 7390 20927
rect 7390 20893 7424 20927
rect 7424 20893 7432 20927
rect 7380 20884 7432 20893
rect 3516 20748 3568 20800
rect 4344 20748 4396 20800
rect 7656 20927 7708 20936
rect 7656 20893 7665 20927
rect 7665 20893 7699 20927
rect 7699 20893 7708 20927
rect 7656 20884 7708 20893
rect 5632 20748 5684 20800
rect 6920 20748 6972 20800
rect 8484 20884 8536 20936
rect 10508 21020 10560 21072
rect 10784 20952 10836 21004
rect 10048 20884 10100 20936
rect 10876 20884 10928 20936
rect 11428 20927 11480 20936
rect 11428 20893 11437 20927
rect 11437 20893 11471 20927
rect 11471 20893 11480 20927
rect 11428 20884 11480 20893
rect 11520 20927 11572 20936
rect 11520 20893 11530 20927
rect 11530 20893 11564 20927
rect 11564 20893 11572 20927
rect 11520 20884 11572 20893
rect 12624 21088 12676 21140
rect 13452 21020 13504 21072
rect 14740 21131 14792 21140
rect 14740 21097 14749 21131
rect 14749 21097 14783 21131
rect 14783 21097 14792 21131
rect 14740 21088 14792 21097
rect 16948 21088 17000 21140
rect 17868 21088 17920 21140
rect 19156 21088 19208 21140
rect 19524 21088 19576 21140
rect 19616 21088 19668 21140
rect 11796 20952 11848 21004
rect 14280 20952 14332 21004
rect 9956 20816 10008 20868
rect 11152 20859 11204 20868
rect 11152 20825 11161 20859
rect 11161 20825 11195 20859
rect 11195 20825 11204 20859
rect 11152 20816 11204 20825
rect 8576 20748 8628 20800
rect 10140 20791 10192 20800
rect 10140 20757 10149 20791
rect 10149 20757 10183 20791
rect 10183 20757 10192 20791
rect 10140 20748 10192 20757
rect 10784 20748 10836 20800
rect 12900 20816 12952 20868
rect 11980 20748 12032 20800
rect 14188 20927 14240 20936
rect 14188 20893 14198 20927
rect 14198 20893 14232 20927
rect 14232 20893 14240 20927
rect 14188 20884 14240 20893
rect 13820 20816 13872 20868
rect 15476 20791 15528 20800
rect 15476 20757 15485 20791
rect 15485 20757 15519 20791
rect 15519 20757 15528 20791
rect 15476 20748 15528 20757
rect 16028 20884 16080 20936
rect 16488 20884 16540 20936
rect 16580 20927 16632 20936
rect 16580 20893 16589 20927
rect 16589 20893 16623 20927
rect 16623 20893 16632 20927
rect 16580 20884 16632 20893
rect 19340 20884 19392 20936
rect 20536 21020 20588 21072
rect 19708 20952 19760 21004
rect 19892 20952 19944 21004
rect 19800 20884 19852 20936
rect 16120 20859 16172 20868
rect 16120 20825 16129 20859
rect 16129 20825 16163 20859
rect 16163 20825 16172 20859
rect 16120 20816 16172 20825
rect 17132 20816 17184 20868
rect 18144 20816 18196 20868
rect 18972 20816 19024 20868
rect 18880 20748 18932 20800
rect 19064 20791 19116 20800
rect 19064 20757 19073 20791
rect 19073 20757 19107 20791
rect 19107 20757 19116 20791
rect 19064 20748 19116 20757
rect 19248 20816 19300 20868
rect 20628 20927 20680 20936
rect 20628 20893 20637 20927
rect 20637 20893 20671 20927
rect 20671 20893 20680 20927
rect 21456 21020 21508 21072
rect 21548 20952 21600 21004
rect 23388 21088 23440 21140
rect 23940 21088 23992 21140
rect 24216 21088 24268 21140
rect 26148 21088 26200 21140
rect 26976 21088 27028 21140
rect 23572 21020 23624 21072
rect 20628 20884 20680 20893
rect 21272 20927 21324 20936
rect 21272 20893 21281 20927
rect 21281 20893 21315 20927
rect 21315 20893 21324 20927
rect 21272 20884 21324 20893
rect 21364 20884 21416 20936
rect 21732 20884 21784 20936
rect 22100 20927 22152 20936
rect 22100 20893 22109 20927
rect 22109 20893 22143 20927
rect 22143 20893 22152 20927
rect 22100 20884 22152 20893
rect 22652 20927 22704 20936
rect 22652 20893 22661 20927
rect 22661 20893 22695 20927
rect 22695 20893 22704 20927
rect 22652 20884 22704 20893
rect 23020 20952 23072 21004
rect 23020 20816 23072 20868
rect 23756 20884 23808 20936
rect 19524 20748 19576 20800
rect 22652 20748 22704 20800
rect 24124 20884 24176 20936
rect 25596 20952 25648 21004
rect 25320 20816 25372 20868
rect 24032 20748 24084 20800
rect 27068 20952 27120 21004
rect 27988 21020 28040 21072
rect 26240 20884 26292 20936
rect 26608 20884 26660 20936
rect 27528 20952 27580 21004
rect 27804 20952 27856 21004
rect 28908 20952 28960 21004
rect 27988 20816 28040 20868
rect 27436 20748 27488 20800
rect 28172 20791 28224 20800
rect 28172 20757 28181 20791
rect 28181 20757 28215 20791
rect 28215 20757 28224 20791
rect 28172 20748 28224 20757
rect 28540 20748 28592 20800
rect 8032 20646 8084 20698
rect 8096 20646 8148 20698
rect 8160 20646 8212 20698
rect 8224 20646 8276 20698
rect 8288 20646 8340 20698
rect 15115 20646 15167 20698
rect 15179 20646 15231 20698
rect 15243 20646 15295 20698
rect 15307 20646 15359 20698
rect 15371 20646 15423 20698
rect 22198 20646 22250 20698
rect 22262 20646 22314 20698
rect 22326 20646 22378 20698
rect 22390 20646 22442 20698
rect 22454 20646 22506 20698
rect 29281 20646 29333 20698
rect 29345 20646 29397 20698
rect 29409 20646 29461 20698
rect 29473 20646 29525 20698
rect 29537 20646 29589 20698
rect 3976 20544 4028 20596
rect 6184 20544 6236 20596
rect 7012 20544 7064 20596
rect 3424 20476 3476 20528
rect 4068 20476 4120 20528
rect 4252 20476 4304 20528
rect 5356 20408 5408 20460
rect 4896 20340 4948 20392
rect 3884 20247 3936 20256
rect 3884 20213 3893 20247
rect 3893 20213 3927 20247
rect 3927 20213 3936 20247
rect 3884 20204 3936 20213
rect 7104 20476 7156 20528
rect 8392 20544 8444 20596
rect 8484 20476 8536 20528
rect 11244 20544 11296 20596
rect 14280 20544 14332 20596
rect 16948 20587 17000 20596
rect 16948 20553 16957 20587
rect 16957 20553 16991 20587
rect 16991 20553 17000 20587
rect 16948 20544 17000 20553
rect 10232 20476 10284 20528
rect 10600 20519 10652 20528
rect 10600 20485 10609 20519
rect 10609 20485 10643 20519
rect 10643 20485 10652 20519
rect 10600 20476 10652 20485
rect 12348 20476 12400 20528
rect 12808 20476 12860 20528
rect 9680 20451 9732 20460
rect 9680 20417 9689 20451
rect 9689 20417 9723 20451
rect 9723 20417 9732 20451
rect 9680 20408 9732 20417
rect 9864 20451 9916 20460
rect 9864 20417 9873 20451
rect 9873 20417 9907 20451
rect 9907 20417 9916 20451
rect 9864 20408 9916 20417
rect 6368 20383 6420 20392
rect 6368 20349 6377 20383
rect 6377 20349 6411 20383
rect 6411 20349 6420 20383
rect 6368 20340 6420 20349
rect 6644 20383 6696 20392
rect 6644 20349 6653 20383
rect 6653 20349 6687 20383
rect 6687 20349 6696 20383
rect 6644 20340 6696 20349
rect 7104 20204 7156 20256
rect 7196 20204 7248 20256
rect 10140 20408 10192 20460
rect 10416 20408 10468 20460
rect 10968 20408 11020 20460
rect 11152 20408 11204 20460
rect 11796 20451 11848 20460
rect 11796 20417 11805 20451
rect 11805 20417 11839 20451
rect 11839 20417 11848 20451
rect 11796 20408 11848 20417
rect 8484 20272 8536 20324
rect 10324 20272 10376 20324
rect 8208 20204 8260 20256
rect 12072 20383 12124 20392
rect 12072 20349 12081 20383
rect 12081 20349 12115 20383
rect 12115 20349 12124 20383
rect 12072 20340 12124 20349
rect 12440 20340 12492 20392
rect 14188 20408 14240 20460
rect 14556 20451 14608 20460
rect 14556 20417 14565 20451
rect 14565 20417 14599 20451
rect 14599 20417 14608 20451
rect 14556 20408 14608 20417
rect 14648 20451 14700 20460
rect 14648 20417 14657 20451
rect 14657 20417 14691 20451
rect 14691 20417 14700 20451
rect 14648 20408 14700 20417
rect 14740 20451 14792 20460
rect 14740 20417 14749 20451
rect 14749 20417 14783 20451
rect 14783 20417 14792 20451
rect 14740 20408 14792 20417
rect 15476 20408 15528 20460
rect 16488 20408 16540 20460
rect 16856 20451 16908 20460
rect 16856 20417 16865 20451
rect 16865 20417 16899 20451
rect 16899 20417 16908 20451
rect 16856 20408 16908 20417
rect 17040 20408 17092 20460
rect 17224 20451 17276 20460
rect 17224 20417 17233 20451
rect 17233 20417 17267 20451
rect 17267 20417 17276 20451
rect 17224 20408 17276 20417
rect 19064 20544 19116 20596
rect 22560 20544 22612 20596
rect 22652 20544 22704 20596
rect 22836 20544 22888 20596
rect 23296 20544 23348 20596
rect 24676 20544 24728 20596
rect 27068 20544 27120 20596
rect 17500 20451 17552 20460
rect 17500 20417 17509 20451
rect 17509 20417 17543 20451
rect 17543 20417 17552 20451
rect 17500 20408 17552 20417
rect 17592 20451 17644 20460
rect 17592 20417 17601 20451
rect 17601 20417 17635 20451
rect 17635 20417 17644 20451
rect 17592 20408 17644 20417
rect 18144 20451 18196 20460
rect 18144 20417 18153 20451
rect 18153 20417 18187 20451
rect 18187 20417 18196 20451
rect 18144 20408 18196 20417
rect 18328 20451 18380 20460
rect 18328 20417 18337 20451
rect 18337 20417 18371 20451
rect 18371 20417 18380 20451
rect 18328 20408 18380 20417
rect 17960 20340 18012 20392
rect 18880 20408 18932 20460
rect 21548 20476 21600 20528
rect 21088 20408 21140 20460
rect 18512 20272 18564 20324
rect 13176 20204 13228 20256
rect 14280 20247 14332 20256
rect 14280 20213 14289 20247
rect 14289 20213 14323 20247
rect 14323 20213 14332 20247
rect 14280 20204 14332 20213
rect 14648 20204 14700 20256
rect 17132 20204 17184 20256
rect 20536 20340 20588 20392
rect 21548 20340 21600 20392
rect 19248 20272 19300 20324
rect 21272 20272 21324 20324
rect 23756 20408 23808 20460
rect 22008 20340 22060 20392
rect 23112 20272 23164 20324
rect 23940 20451 23992 20460
rect 23940 20417 23949 20451
rect 23949 20417 23983 20451
rect 23983 20417 23992 20451
rect 23940 20408 23992 20417
rect 24032 20451 24084 20460
rect 24032 20417 24041 20451
rect 24041 20417 24075 20451
rect 24075 20417 24084 20451
rect 24032 20408 24084 20417
rect 24124 20451 24176 20460
rect 24124 20417 24133 20451
rect 24133 20417 24167 20451
rect 24167 20417 24176 20451
rect 24124 20408 24176 20417
rect 25320 20408 25372 20460
rect 26608 20451 26660 20460
rect 26608 20417 26617 20451
rect 26617 20417 26651 20451
rect 26651 20417 26660 20451
rect 26608 20408 26660 20417
rect 27344 20408 27396 20460
rect 27436 20451 27488 20460
rect 27436 20417 27445 20451
rect 27445 20417 27479 20451
rect 27479 20417 27488 20451
rect 27436 20408 27488 20417
rect 28540 20476 28592 20528
rect 28080 20408 28132 20460
rect 28908 20451 28960 20460
rect 28908 20417 28917 20451
rect 28917 20417 28951 20451
rect 28951 20417 28960 20451
rect 28908 20408 28960 20417
rect 19432 20204 19484 20256
rect 23756 20204 23808 20256
rect 27252 20272 27304 20324
rect 27344 20247 27396 20256
rect 27344 20213 27353 20247
rect 27353 20213 27387 20247
rect 27387 20213 27396 20247
rect 27344 20204 27396 20213
rect 27528 20204 27580 20256
rect 27712 20247 27764 20256
rect 27712 20213 27721 20247
rect 27721 20213 27755 20247
rect 27755 20213 27764 20247
rect 27712 20204 27764 20213
rect 28356 20247 28408 20256
rect 28356 20213 28365 20247
rect 28365 20213 28399 20247
rect 28399 20213 28408 20247
rect 28356 20204 28408 20213
rect 4491 20102 4543 20154
rect 4555 20102 4607 20154
rect 4619 20102 4671 20154
rect 4683 20102 4735 20154
rect 4747 20102 4799 20154
rect 11574 20102 11626 20154
rect 11638 20102 11690 20154
rect 11702 20102 11754 20154
rect 11766 20102 11818 20154
rect 11830 20102 11882 20154
rect 18657 20102 18709 20154
rect 18721 20102 18773 20154
rect 18785 20102 18837 20154
rect 18849 20102 18901 20154
rect 18913 20102 18965 20154
rect 25740 20102 25792 20154
rect 25804 20102 25856 20154
rect 25868 20102 25920 20154
rect 25932 20102 25984 20154
rect 25996 20102 26048 20154
rect 3884 20000 3936 20052
rect 3976 20000 4028 20052
rect 6644 20000 6696 20052
rect 8208 20000 8260 20052
rect 9680 20000 9732 20052
rect 12072 20000 12124 20052
rect 16856 20000 16908 20052
rect 17040 20000 17092 20052
rect 18144 20000 18196 20052
rect 18512 20000 18564 20052
rect 22652 20000 22704 20052
rect 28080 20000 28132 20052
rect 1860 19839 1912 19848
rect 1860 19805 1869 19839
rect 1869 19805 1903 19839
rect 1903 19805 1912 19839
rect 1860 19796 1912 19805
rect 3424 19728 3476 19780
rect 6460 19796 6512 19848
rect 6828 19796 6880 19848
rect 6920 19796 6972 19848
rect 7196 19839 7248 19848
rect 7196 19805 7203 19839
rect 7203 19805 7248 19839
rect 7196 19796 7248 19805
rect 9404 19932 9456 19984
rect 7840 19796 7892 19848
rect 8852 19796 8904 19848
rect 8944 19839 8996 19848
rect 8944 19805 8953 19839
rect 8953 19805 8987 19839
rect 8987 19805 8996 19839
rect 8944 19796 8996 19805
rect 10048 19839 10100 19848
rect 10048 19805 10057 19839
rect 10057 19805 10091 19839
rect 10091 19805 10100 19839
rect 10048 19796 10100 19805
rect 6552 19771 6604 19780
rect 6552 19737 6561 19771
rect 6561 19737 6595 19771
rect 6595 19737 6604 19771
rect 6552 19728 6604 19737
rect 7288 19771 7340 19780
rect 7288 19737 7297 19771
rect 7297 19737 7331 19771
rect 7331 19737 7340 19771
rect 7288 19728 7340 19737
rect 10416 19728 10468 19780
rect 9588 19703 9640 19712
rect 9588 19669 9597 19703
rect 9597 19669 9631 19703
rect 9631 19669 9640 19703
rect 9588 19660 9640 19669
rect 10140 19703 10192 19712
rect 10140 19669 10149 19703
rect 10149 19669 10183 19703
rect 10183 19669 10192 19703
rect 10140 19660 10192 19669
rect 10876 19771 10928 19780
rect 10876 19737 10885 19771
rect 10885 19737 10919 19771
rect 10919 19737 10928 19771
rect 10876 19728 10928 19737
rect 11060 19660 11112 19712
rect 11152 19703 11204 19712
rect 11152 19669 11161 19703
rect 11161 19669 11195 19703
rect 11195 19669 11204 19703
rect 11152 19660 11204 19669
rect 12072 19839 12124 19848
rect 12072 19805 12081 19839
rect 12081 19805 12115 19839
rect 12115 19805 12124 19839
rect 12072 19796 12124 19805
rect 12440 19932 12492 19984
rect 12348 19839 12400 19848
rect 12348 19805 12357 19839
rect 12357 19805 12391 19839
rect 12391 19805 12400 19839
rect 12348 19796 12400 19805
rect 12532 19796 12584 19848
rect 12992 19839 13044 19848
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 12992 19796 13044 19805
rect 13176 19796 13228 19848
rect 14004 19796 14056 19848
rect 14740 19796 14792 19848
rect 17960 19796 18012 19848
rect 27252 19839 27304 19848
rect 27252 19805 27261 19839
rect 27261 19805 27295 19839
rect 27295 19805 27304 19839
rect 27252 19796 27304 19805
rect 27344 19796 27396 19848
rect 27528 19839 27580 19848
rect 14924 19728 14976 19780
rect 15844 19728 15896 19780
rect 16856 19728 16908 19780
rect 23388 19728 23440 19780
rect 27528 19805 27537 19839
rect 27537 19805 27571 19839
rect 27571 19805 27580 19839
rect 27528 19796 27580 19805
rect 27988 19796 28040 19848
rect 28172 19796 28224 19848
rect 12256 19660 12308 19712
rect 12900 19660 12952 19712
rect 14648 19660 14700 19712
rect 17592 19660 17644 19712
rect 19340 19660 19392 19712
rect 19524 19660 19576 19712
rect 19616 19660 19668 19712
rect 19708 19660 19760 19712
rect 26976 19660 27028 19712
rect 27068 19703 27120 19712
rect 27068 19669 27077 19703
rect 27077 19669 27111 19703
rect 27111 19669 27120 19703
rect 27068 19660 27120 19669
rect 27620 19660 27672 19712
rect 28724 19660 28776 19712
rect 8032 19558 8084 19610
rect 8096 19558 8148 19610
rect 8160 19558 8212 19610
rect 8224 19558 8276 19610
rect 8288 19558 8340 19610
rect 15115 19558 15167 19610
rect 15179 19558 15231 19610
rect 15243 19558 15295 19610
rect 15307 19558 15359 19610
rect 15371 19558 15423 19610
rect 22198 19558 22250 19610
rect 22262 19558 22314 19610
rect 22326 19558 22378 19610
rect 22390 19558 22442 19610
rect 22454 19558 22506 19610
rect 29281 19558 29333 19610
rect 29345 19558 29397 19610
rect 29409 19558 29461 19610
rect 29473 19558 29525 19610
rect 29537 19558 29589 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 1492 19363 1544 19372
rect 1492 19329 1501 19363
rect 1501 19329 1535 19363
rect 1535 19329 1544 19363
rect 1492 19320 1544 19329
rect 6552 19320 6604 19372
rect 7012 19320 7064 19372
rect 9588 19456 9640 19508
rect 11060 19456 11112 19508
rect 12256 19456 12308 19508
rect 12532 19456 12584 19508
rect 7748 19388 7800 19440
rect 8484 19388 8536 19440
rect 9772 19388 9824 19440
rect 10876 19388 10928 19440
rect 12624 19388 12676 19440
rect 7656 19363 7708 19372
rect 7656 19329 7665 19363
rect 7665 19329 7699 19363
rect 7699 19329 7708 19363
rect 7656 19320 7708 19329
rect 7932 19363 7984 19372
rect 7932 19329 7941 19363
rect 7941 19329 7975 19363
rect 7975 19329 7984 19363
rect 7932 19320 7984 19329
rect 9864 19320 9916 19372
rect 7840 19252 7892 19304
rect 8852 19252 8904 19304
rect 9220 19252 9272 19304
rect 12164 19252 12216 19304
rect 12900 19320 12952 19372
rect 13268 19456 13320 19508
rect 14556 19456 14608 19508
rect 15200 19456 15252 19508
rect 16120 19456 16172 19508
rect 16856 19456 16908 19508
rect 17224 19499 17276 19508
rect 17224 19465 17233 19499
rect 17233 19465 17267 19499
rect 17267 19465 17276 19499
rect 17224 19456 17276 19465
rect 17960 19456 18012 19508
rect 19064 19499 19116 19508
rect 19064 19465 19073 19499
rect 19073 19465 19107 19499
rect 19107 19465 19116 19499
rect 19064 19456 19116 19465
rect 13176 19363 13228 19372
rect 13176 19329 13185 19363
rect 13185 19329 13219 19363
rect 13219 19329 13228 19363
rect 13176 19320 13228 19329
rect 15108 19363 15160 19372
rect 15108 19329 15117 19363
rect 15117 19329 15151 19363
rect 15151 19329 15160 19363
rect 15108 19320 15160 19329
rect 15292 19363 15344 19372
rect 15292 19329 15301 19363
rect 15301 19329 15335 19363
rect 15335 19329 15344 19363
rect 15292 19320 15344 19329
rect 15568 19320 15620 19372
rect 19708 19456 19760 19508
rect 19892 19499 19944 19508
rect 19892 19465 19901 19499
rect 19901 19465 19935 19499
rect 19935 19465 19944 19499
rect 19892 19456 19944 19465
rect 20536 19499 20588 19508
rect 20536 19465 20545 19499
rect 20545 19465 20579 19499
rect 20579 19465 20588 19499
rect 20536 19456 20588 19465
rect 28080 19456 28132 19508
rect 19432 19388 19484 19440
rect 19616 19431 19668 19440
rect 19616 19397 19625 19431
rect 19625 19397 19659 19431
rect 19659 19397 19668 19431
rect 19616 19388 19668 19397
rect 22560 19388 22612 19440
rect 15936 19252 15988 19304
rect 6460 19184 6512 19236
rect 7840 19159 7892 19168
rect 7840 19125 7849 19159
rect 7849 19125 7883 19159
rect 7883 19125 7892 19159
rect 7840 19116 7892 19125
rect 9588 19184 9640 19236
rect 17960 19184 18012 19236
rect 19340 19363 19392 19372
rect 19340 19329 19349 19363
rect 19349 19329 19383 19363
rect 19383 19329 19392 19363
rect 19340 19320 19392 19329
rect 19524 19363 19576 19372
rect 19524 19329 19533 19363
rect 19533 19329 19567 19363
rect 19567 19329 19576 19363
rect 19524 19320 19576 19329
rect 19616 19252 19668 19304
rect 20076 19320 20128 19372
rect 20168 19363 20220 19372
rect 20168 19329 20177 19363
rect 20177 19329 20211 19363
rect 20211 19329 20220 19363
rect 20168 19320 20220 19329
rect 27436 19320 27488 19372
rect 12624 19116 12676 19168
rect 12716 19116 12768 19168
rect 12900 19116 12952 19168
rect 13728 19116 13780 19168
rect 13820 19116 13872 19168
rect 15016 19116 15068 19168
rect 15476 19159 15528 19168
rect 15476 19125 15485 19159
rect 15485 19125 15519 19159
rect 15519 19125 15528 19159
rect 15476 19116 15528 19125
rect 19800 19184 19852 19236
rect 27804 19295 27856 19304
rect 27804 19261 27813 19295
rect 27813 19261 27847 19295
rect 27847 19261 27856 19295
rect 27804 19252 27856 19261
rect 21272 19116 21324 19168
rect 4491 19014 4543 19066
rect 4555 19014 4607 19066
rect 4619 19014 4671 19066
rect 4683 19014 4735 19066
rect 4747 19014 4799 19066
rect 11574 19014 11626 19066
rect 11638 19014 11690 19066
rect 11702 19014 11754 19066
rect 11766 19014 11818 19066
rect 11830 19014 11882 19066
rect 18657 19014 18709 19066
rect 18721 19014 18773 19066
rect 18785 19014 18837 19066
rect 18849 19014 18901 19066
rect 18913 19014 18965 19066
rect 25740 19014 25792 19066
rect 25804 19014 25856 19066
rect 25868 19014 25920 19066
rect 25932 19014 25984 19066
rect 25996 19014 26048 19066
rect 8944 18912 8996 18964
rect 9588 18955 9640 18964
rect 9588 18921 9597 18955
rect 9597 18921 9631 18955
rect 9631 18921 9640 18955
rect 9588 18912 9640 18921
rect 12164 18912 12216 18964
rect 6368 18776 6420 18828
rect 7840 18776 7892 18828
rect 3516 18708 3568 18760
rect 6460 18751 6512 18760
rect 6460 18717 6469 18751
rect 6469 18717 6503 18751
rect 6503 18717 6512 18751
rect 6460 18708 6512 18717
rect 6920 18708 6972 18760
rect 8576 18708 8628 18760
rect 9220 18776 9272 18828
rect 9956 18776 10008 18828
rect 11152 18776 11204 18828
rect 12808 18912 12860 18964
rect 13176 18912 13228 18964
rect 13820 18912 13872 18964
rect 13912 18912 13964 18964
rect 12624 18844 12676 18896
rect 15476 18844 15528 18896
rect 15568 18844 15620 18896
rect 15936 18955 15988 18964
rect 15936 18921 15945 18955
rect 15945 18921 15979 18955
rect 15979 18921 15988 18955
rect 15936 18912 15988 18921
rect 19432 18912 19484 18964
rect 19892 18912 19944 18964
rect 17684 18844 17736 18896
rect 19156 18844 19208 18896
rect 9404 18751 9456 18760
rect 9404 18717 9418 18751
rect 9418 18717 9452 18751
rect 9452 18717 9456 18751
rect 9404 18708 9456 18717
rect 6276 18640 6328 18692
rect 7012 18640 7064 18692
rect 7288 18640 7340 18692
rect 7748 18640 7800 18692
rect 3976 18572 4028 18624
rect 5264 18572 5316 18624
rect 5816 18572 5868 18624
rect 9312 18572 9364 18624
rect 10692 18572 10744 18624
rect 11060 18572 11112 18624
rect 12532 18776 12584 18828
rect 12716 18708 12768 18760
rect 12348 18640 12400 18692
rect 16488 18708 16540 18760
rect 12716 18572 12768 18624
rect 12808 18615 12860 18624
rect 12808 18581 12817 18615
rect 12817 18581 12851 18615
rect 12851 18581 12860 18615
rect 12808 18572 12860 18581
rect 14372 18640 14424 18692
rect 14556 18640 14608 18692
rect 15476 18640 15528 18692
rect 16764 18708 16816 18760
rect 18788 18708 18840 18760
rect 14740 18572 14792 18624
rect 16120 18615 16172 18624
rect 16120 18581 16129 18615
rect 16129 18581 16163 18615
rect 16163 18581 16172 18615
rect 16120 18572 16172 18581
rect 17500 18572 17552 18624
rect 17684 18683 17736 18692
rect 17684 18649 17693 18683
rect 17693 18649 17727 18683
rect 17727 18649 17736 18683
rect 19800 18708 19852 18760
rect 29460 18844 29512 18896
rect 27712 18708 27764 18760
rect 17684 18640 17736 18649
rect 19432 18683 19484 18692
rect 19432 18649 19441 18683
rect 19441 18649 19475 18683
rect 19475 18649 19484 18683
rect 19432 18640 19484 18649
rect 23296 18640 23348 18692
rect 17960 18615 18012 18624
rect 17960 18581 17969 18615
rect 17969 18581 18003 18615
rect 18003 18581 18012 18615
rect 17960 18572 18012 18581
rect 23940 18572 23992 18624
rect 24492 18572 24544 18624
rect 8032 18470 8084 18522
rect 8096 18470 8148 18522
rect 8160 18470 8212 18522
rect 8224 18470 8276 18522
rect 8288 18470 8340 18522
rect 15115 18470 15167 18522
rect 15179 18470 15231 18522
rect 15243 18470 15295 18522
rect 15307 18470 15359 18522
rect 15371 18470 15423 18522
rect 22198 18470 22250 18522
rect 22262 18470 22314 18522
rect 22326 18470 22378 18522
rect 22390 18470 22442 18522
rect 22454 18470 22506 18522
rect 29281 18470 29333 18522
rect 29345 18470 29397 18522
rect 29409 18470 29461 18522
rect 29473 18470 29525 18522
rect 29537 18470 29589 18522
rect 1860 18368 1912 18420
rect 3700 18368 3752 18420
rect 6276 18368 6328 18420
rect 9312 18368 9364 18420
rect 9680 18368 9732 18420
rect 5264 18300 5316 18352
rect 3240 18232 3292 18284
rect 3700 18275 3752 18284
rect 3700 18241 3709 18275
rect 3709 18241 3743 18275
rect 3743 18241 3752 18275
rect 3700 18232 3752 18241
rect 3424 18164 3476 18216
rect 3516 18164 3568 18216
rect 5264 18164 5316 18216
rect 5080 18096 5132 18148
rect 5172 18028 5224 18080
rect 5724 18232 5776 18284
rect 6276 18232 6328 18284
rect 6736 18232 6788 18284
rect 6552 18164 6604 18216
rect 6920 18232 6972 18284
rect 7656 18232 7708 18284
rect 7840 18232 7892 18284
rect 7012 18164 7064 18216
rect 7564 18207 7616 18216
rect 7564 18173 7573 18207
rect 7573 18173 7607 18207
rect 7607 18173 7616 18207
rect 7564 18164 7616 18173
rect 7104 18096 7156 18148
rect 12624 18368 12676 18420
rect 12716 18368 12768 18420
rect 14372 18368 14424 18420
rect 13912 18300 13964 18352
rect 9680 18275 9732 18284
rect 9680 18241 9689 18275
rect 9689 18241 9723 18275
rect 9723 18241 9732 18275
rect 9680 18232 9732 18241
rect 9772 18275 9824 18284
rect 9772 18241 9781 18275
rect 9781 18241 9815 18275
rect 9815 18241 9824 18275
rect 9772 18232 9824 18241
rect 9496 18096 9548 18148
rect 10232 18275 10284 18284
rect 10232 18241 10241 18275
rect 10241 18241 10275 18275
rect 10275 18241 10284 18275
rect 10232 18232 10284 18241
rect 12624 18275 12676 18284
rect 12624 18241 12633 18275
rect 12633 18241 12667 18275
rect 12667 18241 12676 18275
rect 12624 18232 12676 18241
rect 10324 18164 10376 18216
rect 11244 18164 11296 18216
rect 11336 18164 11388 18216
rect 12900 18275 12952 18284
rect 12900 18241 12909 18275
rect 12909 18241 12943 18275
rect 12943 18241 12952 18275
rect 12900 18232 12952 18241
rect 13360 18232 13412 18284
rect 16580 18368 16632 18420
rect 15476 18300 15528 18352
rect 17960 18368 18012 18420
rect 18144 18368 18196 18420
rect 18788 18411 18840 18420
rect 18788 18377 18797 18411
rect 18797 18377 18831 18411
rect 18831 18377 18840 18411
rect 18788 18368 18840 18377
rect 19984 18368 20036 18420
rect 20168 18300 20220 18352
rect 13820 18164 13872 18216
rect 15476 18164 15528 18216
rect 15568 18164 15620 18216
rect 18052 18164 18104 18216
rect 19064 18232 19116 18284
rect 19432 18275 19484 18284
rect 19432 18241 19441 18275
rect 19441 18241 19475 18275
rect 19475 18241 19484 18275
rect 19432 18232 19484 18241
rect 19524 18232 19576 18284
rect 19800 18275 19852 18284
rect 19800 18241 19809 18275
rect 19809 18241 19843 18275
rect 19843 18241 19852 18275
rect 19800 18232 19852 18241
rect 18512 18164 18564 18216
rect 19248 18207 19300 18216
rect 19248 18173 19257 18207
rect 19257 18173 19291 18207
rect 19291 18173 19300 18207
rect 19248 18164 19300 18173
rect 20444 18275 20496 18284
rect 20444 18241 20454 18275
rect 20454 18241 20488 18275
rect 20488 18241 20496 18275
rect 20444 18232 20496 18241
rect 20720 18275 20772 18284
rect 20720 18241 20729 18275
rect 20729 18241 20763 18275
rect 20763 18241 20772 18275
rect 20720 18232 20772 18241
rect 25320 18368 25372 18420
rect 23480 18300 23532 18352
rect 24492 18300 24544 18352
rect 24952 18300 25004 18352
rect 28632 18232 28684 18284
rect 7656 18028 7708 18080
rect 9864 18028 9916 18080
rect 10048 18028 10100 18080
rect 10140 18028 10192 18080
rect 10692 18028 10744 18080
rect 12072 18028 12124 18080
rect 14740 18096 14792 18148
rect 16764 18096 16816 18148
rect 18328 18096 18380 18148
rect 23204 18207 23256 18216
rect 23204 18173 23213 18207
rect 23213 18173 23247 18207
rect 23247 18173 23256 18207
rect 23204 18164 23256 18173
rect 23664 18164 23716 18216
rect 25504 18164 25556 18216
rect 26884 18164 26936 18216
rect 27252 18207 27304 18216
rect 27252 18173 27261 18207
rect 27261 18173 27295 18207
rect 27295 18173 27304 18207
rect 27252 18164 27304 18173
rect 29000 18207 29052 18216
rect 29000 18173 29009 18207
rect 29009 18173 29043 18207
rect 29043 18173 29052 18207
rect 29000 18164 29052 18173
rect 21088 18096 21140 18148
rect 25228 18096 25280 18148
rect 26424 18096 26476 18148
rect 16120 18028 16172 18080
rect 24860 18028 24912 18080
rect 4491 17926 4543 17978
rect 4555 17926 4607 17978
rect 4619 17926 4671 17978
rect 4683 17926 4735 17978
rect 4747 17926 4799 17978
rect 11574 17926 11626 17978
rect 11638 17926 11690 17978
rect 11702 17926 11754 17978
rect 11766 17926 11818 17978
rect 11830 17926 11882 17978
rect 18657 17926 18709 17978
rect 18721 17926 18773 17978
rect 18785 17926 18837 17978
rect 18849 17926 18901 17978
rect 18913 17926 18965 17978
rect 25740 17926 25792 17978
rect 25804 17926 25856 17978
rect 25868 17926 25920 17978
rect 25932 17926 25984 17978
rect 25996 17926 26048 17978
rect 3240 17824 3292 17876
rect 5264 17824 5316 17876
rect 3700 17688 3752 17740
rect 5172 17620 5224 17672
rect 7748 17824 7800 17876
rect 11060 17824 11112 17876
rect 11336 17867 11388 17876
rect 11336 17833 11345 17867
rect 11345 17833 11379 17867
rect 11379 17833 11388 17867
rect 11336 17824 11388 17833
rect 12624 17824 12676 17876
rect 13912 17867 13964 17876
rect 13912 17833 13921 17867
rect 13921 17833 13955 17867
rect 13955 17833 13964 17867
rect 13912 17824 13964 17833
rect 19800 17867 19852 17876
rect 19800 17833 19809 17867
rect 19809 17833 19843 17867
rect 19843 17833 19852 17867
rect 19800 17824 19852 17833
rect 20720 17824 20772 17876
rect 21824 17867 21876 17876
rect 21824 17833 21833 17867
rect 21833 17833 21867 17867
rect 21867 17833 21876 17867
rect 21824 17824 21876 17833
rect 22468 17824 22520 17876
rect 22652 17824 22704 17876
rect 22836 17824 22888 17876
rect 23204 17824 23256 17876
rect 23388 17824 23440 17876
rect 25136 17824 25188 17876
rect 25872 17824 25924 17876
rect 26792 17824 26844 17876
rect 27252 17824 27304 17876
rect 7564 17756 7616 17808
rect 7288 17663 7340 17672
rect 7288 17629 7297 17663
rect 7297 17629 7331 17663
rect 7331 17629 7340 17663
rect 7288 17620 7340 17629
rect 9956 17688 10008 17740
rect 3424 17552 3476 17604
rect 4528 17552 4580 17604
rect 4804 17552 4856 17604
rect 5816 17552 5868 17604
rect 7104 17595 7156 17604
rect 7104 17561 7113 17595
rect 7113 17561 7147 17595
rect 7147 17561 7156 17595
rect 7104 17552 7156 17561
rect 5172 17484 5224 17536
rect 5448 17484 5500 17536
rect 6368 17484 6420 17536
rect 7656 17663 7708 17672
rect 7656 17629 7665 17663
rect 7665 17629 7699 17663
rect 7699 17629 7708 17663
rect 7656 17620 7708 17629
rect 18604 17756 18656 17808
rect 11244 17620 11296 17672
rect 11428 17663 11480 17672
rect 11428 17629 11437 17663
rect 11437 17629 11471 17663
rect 11471 17629 11480 17663
rect 11428 17620 11480 17629
rect 19340 17688 19392 17740
rect 10140 17552 10192 17604
rect 11152 17552 11204 17604
rect 11980 17620 12032 17672
rect 16120 17663 16172 17672
rect 16120 17629 16129 17663
rect 16129 17629 16163 17663
rect 16163 17629 16172 17663
rect 16120 17620 16172 17629
rect 18604 17620 18656 17672
rect 13176 17552 13228 17604
rect 14188 17595 14240 17604
rect 14188 17561 14197 17595
rect 14197 17561 14231 17595
rect 14231 17561 14240 17595
rect 14188 17552 14240 17561
rect 17592 17595 17644 17604
rect 17592 17561 17601 17595
rect 17601 17561 17635 17595
rect 17635 17561 17644 17595
rect 17592 17552 17644 17561
rect 14648 17484 14700 17536
rect 16396 17484 16448 17536
rect 16672 17527 16724 17536
rect 16672 17493 16681 17527
rect 16681 17493 16715 17527
rect 16715 17493 16724 17527
rect 16672 17484 16724 17493
rect 17132 17484 17184 17536
rect 17868 17484 17920 17536
rect 18420 17484 18472 17536
rect 19984 17620 20036 17672
rect 22652 17688 22704 17740
rect 22468 17620 22520 17672
rect 22560 17620 22612 17672
rect 20260 17552 20312 17604
rect 20352 17595 20404 17604
rect 20352 17561 20361 17595
rect 20361 17561 20395 17595
rect 20395 17561 20404 17595
rect 20352 17552 20404 17561
rect 21824 17552 21876 17604
rect 23296 17620 23348 17672
rect 23756 17688 23808 17740
rect 25504 17756 25556 17808
rect 24860 17688 24912 17740
rect 26240 17756 26292 17808
rect 26700 17756 26752 17808
rect 26976 17756 27028 17808
rect 26424 17731 26476 17740
rect 26424 17697 26433 17731
rect 26433 17697 26467 17731
rect 26467 17697 26476 17731
rect 26424 17688 26476 17697
rect 26516 17731 26568 17740
rect 26516 17697 26525 17731
rect 26525 17697 26559 17731
rect 26559 17697 26568 17731
rect 27896 17756 27948 17808
rect 26516 17688 26568 17697
rect 24768 17620 24820 17672
rect 25136 17663 25188 17672
rect 25136 17629 25145 17663
rect 25145 17629 25179 17663
rect 25179 17629 25188 17663
rect 25136 17620 25188 17629
rect 25320 17663 25372 17672
rect 25320 17629 25329 17663
rect 25329 17629 25363 17663
rect 25363 17629 25372 17663
rect 25320 17620 25372 17629
rect 25872 17620 25924 17672
rect 25964 17620 26016 17672
rect 26608 17663 26660 17672
rect 26608 17629 26617 17663
rect 26617 17629 26651 17663
rect 26651 17629 26660 17663
rect 26608 17620 26660 17629
rect 23572 17595 23624 17604
rect 23572 17561 23581 17595
rect 23581 17561 23615 17595
rect 23615 17561 23624 17595
rect 23572 17552 23624 17561
rect 19064 17527 19116 17536
rect 19064 17493 19073 17527
rect 19073 17493 19107 17527
rect 19107 17493 19116 17527
rect 19064 17484 19116 17493
rect 19432 17484 19484 17536
rect 23112 17484 23164 17536
rect 24032 17552 24084 17604
rect 24860 17484 24912 17536
rect 25412 17595 25464 17604
rect 25412 17561 25421 17595
rect 25421 17561 25455 17595
rect 25455 17561 25464 17595
rect 25412 17552 25464 17561
rect 26792 17595 26844 17604
rect 26792 17561 26801 17595
rect 26801 17561 26835 17595
rect 26835 17561 26844 17595
rect 26792 17552 26844 17561
rect 27160 17620 27212 17672
rect 28448 17688 28500 17740
rect 29000 17688 29052 17740
rect 26148 17484 26200 17536
rect 26240 17527 26292 17536
rect 26240 17493 26249 17527
rect 26249 17493 26283 17527
rect 26283 17493 26292 17527
rect 26240 17484 26292 17493
rect 26424 17484 26476 17536
rect 27528 17552 27580 17604
rect 27712 17484 27764 17536
rect 27988 17527 28040 17536
rect 27988 17493 27997 17527
rect 27997 17493 28031 17527
rect 28031 17493 28040 17527
rect 27988 17484 28040 17493
rect 28080 17484 28132 17536
rect 28356 17484 28408 17536
rect 8032 17382 8084 17434
rect 8096 17382 8148 17434
rect 8160 17382 8212 17434
rect 8224 17382 8276 17434
rect 8288 17382 8340 17434
rect 15115 17382 15167 17434
rect 15179 17382 15231 17434
rect 15243 17382 15295 17434
rect 15307 17382 15359 17434
rect 15371 17382 15423 17434
rect 22198 17382 22250 17434
rect 22262 17382 22314 17434
rect 22326 17382 22378 17434
rect 22390 17382 22442 17434
rect 22454 17382 22506 17434
rect 29281 17382 29333 17434
rect 29345 17382 29397 17434
rect 29409 17382 29461 17434
rect 29473 17382 29525 17434
rect 29537 17382 29589 17434
rect 3700 17280 3752 17332
rect 4344 17280 4396 17332
rect 4528 17323 4580 17332
rect 4528 17289 4537 17323
rect 4537 17289 4571 17323
rect 4571 17289 4580 17323
rect 4528 17280 4580 17289
rect 5080 17280 5132 17332
rect 4804 17255 4856 17264
rect 4804 17221 4813 17255
rect 4813 17221 4847 17255
rect 4847 17221 4856 17255
rect 4804 17212 4856 17221
rect 3516 17076 3568 17128
rect 3792 17144 3844 17196
rect 3976 17187 4028 17196
rect 3976 17153 3985 17187
rect 3985 17153 4019 17187
rect 4019 17153 4028 17187
rect 3976 17144 4028 17153
rect 4068 17144 4120 17196
rect 4252 17187 4304 17196
rect 4252 17153 4261 17187
rect 4261 17153 4295 17187
rect 4295 17153 4304 17187
rect 4252 17144 4304 17153
rect 4344 17187 4396 17196
rect 4344 17153 4377 17187
rect 4377 17153 4396 17187
rect 4344 17144 4396 17153
rect 4528 17144 4580 17196
rect 5448 17255 5500 17264
rect 5448 17221 5457 17255
rect 5457 17221 5491 17255
rect 5491 17221 5500 17255
rect 5448 17212 5500 17221
rect 9956 17280 10008 17332
rect 4804 17076 4856 17128
rect 5264 17187 5316 17196
rect 5264 17153 5273 17187
rect 5273 17153 5307 17187
rect 5307 17153 5316 17187
rect 5264 17144 5316 17153
rect 5540 17187 5592 17196
rect 5540 17153 5549 17187
rect 5549 17153 5583 17187
rect 5583 17153 5592 17187
rect 5540 17144 5592 17153
rect 5908 17144 5960 17196
rect 6000 17144 6052 17196
rect 11336 17212 11388 17264
rect 11888 17212 11940 17264
rect 12808 17280 12860 17332
rect 13820 17280 13872 17332
rect 13176 17212 13228 17264
rect 9864 17119 9916 17128
rect 9864 17085 9873 17119
rect 9873 17085 9907 17119
rect 9907 17085 9916 17119
rect 9864 17076 9916 17085
rect 13912 17144 13964 17196
rect 16672 17280 16724 17332
rect 16764 17280 16816 17332
rect 16028 17212 16080 17264
rect 16120 17212 16172 17264
rect 15108 17144 15160 17196
rect 11060 17076 11112 17128
rect 5172 17008 5224 17060
rect 5264 17008 5316 17060
rect 11244 17008 11296 17060
rect 3332 16940 3384 16992
rect 4988 16940 5040 16992
rect 5816 16983 5868 16992
rect 5816 16949 5825 16983
rect 5825 16949 5859 16983
rect 5859 16949 5868 16983
rect 5816 16940 5868 16949
rect 7748 16940 7800 16992
rect 14096 16940 14148 16992
rect 15844 17144 15896 17196
rect 15476 17076 15528 17128
rect 17132 17187 17184 17196
rect 17132 17153 17141 17187
rect 17141 17153 17175 17187
rect 17175 17153 17184 17187
rect 17132 17144 17184 17153
rect 17592 17280 17644 17332
rect 19064 17280 19116 17332
rect 19248 17323 19300 17332
rect 19248 17289 19257 17323
rect 19257 17289 19291 17323
rect 19291 17289 19300 17323
rect 19248 17280 19300 17289
rect 20352 17280 20404 17332
rect 18328 17144 18380 17196
rect 16580 17076 16632 17128
rect 18512 17187 18564 17196
rect 18512 17153 18521 17187
rect 18521 17153 18555 17187
rect 18555 17153 18564 17187
rect 18512 17144 18564 17153
rect 16488 16940 16540 16992
rect 19064 17187 19116 17196
rect 19064 17153 19073 17187
rect 19073 17153 19107 17187
rect 19107 17153 19116 17187
rect 19064 17144 19116 17153
rect 21824 17144 21876 17196
rect 22192 17187 22244 17196
rect 22192 17153 22201 17187
rect 22201 17153 22235 17187
rect 22235 17153 22244 17187
rect 22192 17144 22244 17153
rect 22836 17280 22888 17332
rect 23572 17280 23624 17332
rect 22560 17212 22612 17264
rect 23664 17212 23716 17264
rect 25136 17280 25188 17332
rect 25412 17280 25464 17332
rect 26240 17280 26292 17332
rect 26608 17280 26660 17332
rect 25504 17212 25556 17264
rect 22836 17187 22888 17196
rect 22836 17153 22845 17187
rect 22845 17153 22879 17187
rect 22879 17153 22888 17187
rect 22836 17144 22888 17153
rect 23480 17187 23532 17196
rect 23480 17153 23489 17187
rect 23489 17153 23523 17187
rect 23523 17153 23532 17187
rect 23480 17144 23532 17153
rect 24768 17144 24820 17196
rect 22284 17008 22336 17060
rect 23388 17076 23440 17128
rect 25228 17144 25280 17196
rect 25412 17187 25464 17196
rect 25412 17153 25421 17187
rect 25421 17153 25455 17187
rect 25455 17153 25464 17187
rect 25412 17144 25464 17153
rect 26056 17187 26108 17196
rect 26056 17153 26065 17187
rect 26065 17153 26099 17187
rect 26099 17153 26108 17187
rect 26056 17144 26108 17153
rect 24952 17076 25004 17128
rect 25964 17076 26016 17128
rect 23112 16983 23164 16992
rect 23112 16949 23121 16983
rect 23121 16949 23155 16983
rect 23155 16949 23164 16983
rect 23112 16940 23164 16949
rect 23572 16940 23624 16992
rect 24860 16940 24912 16992
rect 25872 17008 25924 17060
rect 27252 17144 27304 17196
rect 27528 17212 27580 17264
rect 27804 17144 27856 17196
rect 27896 17187 27948 17196
rect 27896 17153 27905 17187
rect 27905 17153 27939 17187
rect 27939 17153 27948 17187
rect 27896 17144 27948 17153
rect 28448 17255 28500 17264
rect 28448 17221 28457 17255
rect 28457 17221 28491 17255
rect 28491 17221 28500 17255
rect 28448 17212 28500 17221
rect 26700 17076 26752 17128
rect 26976 17076 27028 17128
rect 27160 17008 27212 17060
rect 27528 17076 27580 17128
rect 28356 17144 28408 17196
rect 26424 16940 26476 16992
rect 26516 16983 26568 16992
rect 26516 16949 26525 16983
rect 26525 16949 26559 16983
rect 26559 16949 26568 16983
rect 26516 16940 26568 16949
rect 28448 17076 28500 17128
rect 28632 17076 28684 17128
rect 27988 16940 28040 16992
rect 28356 16940 28408 16992
rect 28632 16983 28684 16992
rect 28632 16949 28641 16983
rect 28641 16949 28675 16983
rect 28675 16949 28684 16983
rect 28632 16940 28684 16949
rect 4491 16838 4543 16890
rect 4555 16838 4607 16890
rect 4619 16838 4671 16890
rect 4683 16838 4735 16890
rect 4747 16838 4799 16890
rect 11574 16838 11626 16890
rect 11638 16838 11690 16890
rect 11702 16838 11754 16890
rect 11766 16838 11818 16890
rect 11830 16838 11882 16890
rect 18657 16838 18709 16890
rect 18721 16838 18773 16890
rect 18785 16838 18837 16890
rect 18849 16838 18901 16890
rect 18913 16838 18965 16890
rect 25740 16838 25792 16890
rect 25804 16838 25856 16890
rect 25868 16838 25920 16890
rect 25932 16838 25984 16890
rect 25996 16838 26048 16890
rect 5540 16736 5592 16788
rect 14648 16779 14700 16788
rect 14648 16745 14657 16779
rect 14657 16745 14691 16779
rect 14691 16745 14700 16779
rect 14648 16736 14700 16745
rect 15108 16736 15160 16788
rect 20444 16736 20496 16788
rect 22192 16736 22244 16788
rect 22284 16736 22336 16788
rect 22560 16736 22612 16788
rect 22836 16736 22888 16788
rect 23756 16779 23808 16788
rect 23756 16745 23765 16779
rect 23765 16745 23799 16779
rect 23799 16745 23808 16779
rect 23756 16736 23808 16745
rect 25320 16736 25372 16788
rect 26792 16736 26844 16788
rect 26976 16736 27028 16788
rect 27528 16736 27580 16788
rect 27804 16779 27856 16788
rect 27804 16745 27813 16779
rect 27813 16745 27847 16779
rect 27847 16745 27856 16779
rect 27804 16736 27856 16745
rect 27896 16736 27948 16788
rect 5080 16668 5132 16720
rect 6920 16668 6972 16720
rect 14372 16668 14424 16720
rect 14556 16668 14608 16720
rect 23296 16711 23348 16720
rect 23296 16677 23305 16711
rect 23305 16677 23339 16711
rect 23339 16677 23348 16711
rect 23296 16668 23348 16677
rect 4252 16600 4304 16652
rect 4896 16600 4948 16652
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 1676 16507 1728 16516
rect 1676 16473 1685 16507
rect 1685 16473 1719 16507
rect 1719 16473 1728 16507
rect 1676 16464 1728 16473
rect 3884 16464 3936 16516
rect 4436 16439 4488 16448
rect 4436 16405 4445 16439
rect 4445 16405 4479 16439
rect 4479 16405 4488 16439
rect 4436 16396 4488 16405
rect 5080 16532 5132 16584
rect 5356 16575 5408 16584
rect 5356 16541 5365 16575
rect 5365 16541 5399 16575
rect 5399 16541 5408 16575
rect 5356 16532 5408 16541
rect 5724 16575 5776 16584
rect 5724 16541 5733 16575
rect 5733 16541 5767 16575
rect 5767 16541 5776 16575
rect 5724 16532 5776 16541
rect 6460 16532 6512 16584
rect 9680 16532 9732 16584
rect 9864 16575 9916 16584
rect 9864 16541 9873 16575
rect 9873 16541 9907 16575
rect 9907 16541 9916 16575
rect 9864 16532 9916 16541
rect 10968 16600 11020 16652
rect 14004 16600 14056 16652
rect 12256 16532 12308 16584
rect 14096 16575 14148 16584
rect 14096 16541 14105 16575
rect 14105 16541 14139 16575
rect 14139 16541 14148 16575
rect 14096 16532 14148 16541
rect 14648 16532 14700 16584
rect 15016 16532 15068 16584
rect 16580 16600 16632 16652
rect 19064 16600 19116 16652
rect 21824 16600 21876 16652
rect 7472 16464 7524 16516
rect 10048 16507 10100 16516
rect 10048 16473 10057 16507
rect 10057 16473 10091 16507
rect 10091 16473 10100 16507
rect 10048 16464 10100 16473
rect 5448 16396 5500 16448
rect 5540 16439 5592 16448
rect 5540 16405 5549 16439
rect 5549 16405 5583 16439
rect 5583 16405 5592 16439
rect 5540 16396 5592 16405
rect 9956 16396 10008 16448
rect 10232 16396 10284 16448
rect 10416 16439 10468 16448
rect 10416 16405 10425 16439
rect 10425 16405 10459 16439
rect 10459 16405 10468 16439
rect 10416 16396 10468 16405
rect 10508 16396 10560 16448
rect 12348 16396 12400 16448
rect 12716 16396 12768 16448
rect 14372 16507 14424 16516
rect 14372 16473 14381 16507
rect 14381 16473 14415 16507
rect 14415 16473 14424 16507
rect 14372 16464 14424 16473
rect 14924 16464 14976 16516
rect 15660 16532 15712 16584
rect 15752 16464 15804 16516
rect 17132 16464 17184 16516
rect 14832 16439 14884 16448
rect 14832 16405 14841 16439
rect 14841 16405 14875 16439
rect 14875 16405 14884 16439
rect 14832 16396 14884 16405
rect 15016 16396 15068 16448
rect 22652 16532 22704 16584
rect 23112 16396 23164 16448
rect 23204 16439 23256 16448
rect 23204 16405 23213 16439
rect 23213 16405 23247 16439
rect 23247 16405 23256 16439
rect 23204 16396 23256 16405
rect 23664 16532 23716 16584
rect 23940 16532 23992 16584
rect 24676 16532 24728 16584
rect 25596 16600 25648 16652
rect 26424 16668 26476 16720
rect 23756 16464 23808 16516
rect 25504 16575 25556 16584
rect 25504 16541 25513 16575
rect 25513 16541 25547 16575
rect 25547 16541 25556 16575
rect 25504 16532 25556 16541
rect 26148 16532 26200 16584
rect 27988 16600 28040 16652
rect 26700 16507 26752 16516
rect 26700 16473 26709 16507
rect 26709 16473 26743 16507
rect 26743 16473 26752 16507
rect 26700 16464 26752 16473
rect 27620 16575 27672 16584
rect 27620 16541 27629 16575
rect 27629 16541 27663 16575
rect 27663 16541 27672 16575
rect 27620 16532 27672 16541
rect 27896 16532 27948 16584
rect 28356 16575 28408 16584
rect 28356 16541 28373 16575
rect 28373 16541 28407 16575
rect 28407 16541 28408 16575
rect 28356 16532 28408 16541
rect 28632 16532 28684 16584
rect 26056 16396 26108 16448
rect 26424 16396 26476 16448
rect 26608 16396 26660 16448
rect 27252 16439 27304 16448
rect 27252 16405 27261 16439
rect 27261 16405 27295 16439
rect 27295 16405 27304 16439
rect 27252 16396 27304 16405
rect 27988 16439 28040 16448
rect 27988 16405 27997 16439
rect 27997 16405 28031 16439
rect 28031 16405 28040 16439
rect 27988 16396 28040 16405
rect 8032 16294 8084 16346
rect 8096 16294 8148 16346
rect 8160 16294 8212 16346
rect 8224 16294 8276 16346
rect 8288 16294 8340 16346
rect 15115 16294 15167 16346
rect 15179 16294 15231 16346
rect 15243 16294 15295 16346
rect 15307 16294 15359 16346
rect 15371 16294 15423 16346
rect 22198 16294 22250 16346
rect 22262 16294 22314 16346
rect 22326 16294 22378 16346
rect 22390 16294 22442 16346
rect 22454 16294 22506 16346
rect 29281 16294 29333 16346
rect 29345 16294 29397 16346
rect 29409 16294 29461 16346
rect 29473 16294 29525 16346
rect 29537 16294 29589 16346
rect 1676 16192 1728 16244
rect 4436 16192 4488 16244
rect 4988 16235 5040 16244
rect 4988 16201 4997 16235
rect 4997 16201 5031 16235
rect 5031 16201 5040 16235
rect 4988 16192 5040 16201
rect 5448 16192 5500 16244
rect 6276 16192 6328 16244
rect 940 16056 992 16108
rect 3884 16056 3936 16108
rect 5448 16056 5500 16108
rect 5632 16056 5684 16108
rect 5724 16056 5776 16108
rect 6184 16056 6236 16108
rect 6552 16124 6604 16176
rect 7564 16192 7616 16244
rect 6920 16124 6972 16176
rect 7748 16124 7800 16176
rect 1400 15988 1452 16040
rect 4344 15920 4396 15972
rect 7472 16099 7524 16108
rect 7472 16065 7481 16099
rect 7481 16065 7515 16099
rect 7515 16065 7524 16099
rect 7472 16056 7524 16065
rect 7932 16099 7984 16108
rect 7932 16065 7941 16099
rect 7941 16065 7975 16099
rect 7975 16065 7984 16099
rect 7932 16056 7984 16065
rect 22836 16192 22888 16244
rect 10048 16099 10100 16108
rect 10048 16065 10057 16099
rect 10057 16065 10091 16099
rect 10091 16065 10100 16099
rect 10048 16056 10100 16065
rect 10140 16099 10192 16108
rect 10140 16065 10149 16099
rect 10149 16065 10183 16099
rect 10183 16065 10192 16099
rect 10140 16056 10192 16065
rect 10324 16056 10376 16108
rect 8208 16031 8260 16040
rect 8208 15997 8217 16031
rect 8217 15997 8251 16031
rect 8251 15997 8260 16031
rect 8208 15988 8260 15997
rect 8668 16031 8720 16040
rect 8668 15997 8677 16031
rect 8677 15997 8711 16031
rect 8711 15997 8720 16031
rect 8668 15988 8720 15997
rect 10508 16031 10560 16040
rect 8392 15920 8444 15972
rect 10508 15997 10517 16031
rect 10517 15997 10551 16031
rect 10551 15997 10560 16031
rect 10508 15988 10560 15997
rect 11060 15988 11112 16040
rect 12900 16124 12952 16176
rect 12624 16056 12676 16108
rect 13176 16099 13228 16108
rect 13176 16065 13185 16099
rect 13185 16065 13219 16099
rect 13219 16065 13228 16099
rect 13176 16056 13228 16065
rect 13360 16099 13412 16108
rect 13360 16065 13369 16099
rect 13369 16065 13403 16099
rect 13403 16065 13412 16099
rect 13360 16056 13412 16065
rect 13912 16056 13964 16108
rect 13636 15988 13688 16040
rect 23204 16124 23256 16176
rect 26700 16192 26752 16244
rect 27344 16192 27396 16244
rect 27804 16192 27856 16244
rect 14832 16056 14884 16108
rect 15476 16056 15528 16108
rect 15844 16056 15896 16108
rect 16488 16056 16540 16108
rect 23940 16056 23992 16108
rect 15016 15988 15068 16040
rect 9864 15920 9916 15972
rect 10140 15920 10192 15972
rect 9956 15852 10008 15904
rect 12348 15920 12400 15972
rect 13084 15920 13136 15972
rect 25504 15988 25556 16040
rect 26608 16056 26660 16108
rect 23388 15920 23440 15972
rect 23664 15963 23716 15972
rect 23664 15929 23673 15963
rect 23673 15929 23707 15963
rect 23707 15929 23716 15963
rect 23664 15920 23716 15929
rect 13820 15852 13872 15904
rect 15476 15852 15528 15904
rect 15752 15852 15804 15904
rect 15936 15852 15988 15904
rect 16120 15852 16172 15904
rect 16304 15895 16356 15904
rect 16304 15861 16313 15895
rect 16313 15861 16347 15895
rect 16347 15861 16356 15895
rect 16304 15852 16356 15861
rect 26148 15852 26200 15904
rect 4491 15750 4543 15802
rect 4555 15750 4607 15802
rect 4619 15750 4671 15802
rect 4683 15750 4735 15802
rect 4747 15750 4799 15802
rect 11574 15750 11626 15802
rect 11638 15750 11690 15802
rect 11702 15750 11754 15802
rect 11766 15750 11818 15802
rect 11830 15750 11882 15802
rect 18657 15750 18709 15802
rect 18721 15750 18773 15802
rect 18785 15750 18837 15802
rect 18849 15750 18901 15802
rect 18913 15750 18965 15802
rect 25740 15750 25792 15802
rect 25804 15750 25856 15802
rect 25868 15750 25920 15802
rect 25932 15750 25984 15802
rect 25996 15750 26048 15802
rect 4344 15648 4396 15700
rect 5724 15648 5776 15700
rect 7932 15648 7984 15700
rect 1400 15512 1452 15564
rect 3332 15512 3384 15564
rect 3240 15444 3292 15496
rect 3884 15444 3936 15496
rect 4068 15444 4120 15496
rect 7564 15512 7616 15564
rect 5816 15444 5868 15496
rect 6644 15487 6696 15496
rect 6644 15453 6653 15487
rect 6653 15453 6687 15487
rect 6687 15453 6696 15487
rect 6644 15444 6696 15453
rect 7932 15444 7984 15496
rect 8208 15444 8260 15496
rect 8668 15648 8720 15700
rect 9956 15648 10008 15700
rect 10784 15648 10836 15700
rect 11060 15648 11112 15700
rect 11704 15648 11756 15700
rect 12164 15648 12216 15700
rect 16120 15691 16172 15700
rect 16120 15657 16129 15691
rect 16129 15657 16163 15691
rect 16163 15657 16172 15691
rect 16120 15648 16172 15657
rect 16304 15648 16356 15700
rect 10140 15512 10192 15564
rect 9220 15487 9272 15496
rect 9220 15453 9229 15487
rect 9229 15453 9263 15487
rect 9263 15453 9272 15487
rect 9220 15444 9272 15453
rect 12624 15555 12676 15564
rect 12624 15521 12633 15555
rect 12633 15521 12667 15555
rect 12667 15521 12676 15555
rect 12624 15512 12676 15521
rect 13084 15512 13136 15564
rect 9588 15376 9640 15428
rect 9956 15376 10008 15428
rect 11796 15376 11848 15428
rect 12256 15487 12308 15496
rect 12256 15453 12265 15487
rect 12265 15453 12299 15487
rect 12299 15453 12308 15487
rect 12256 15444 12308 15453
rect 12716 15444 12768 15496
rect 13912 15444 13964 15496
rect 14372 15487 14424 15496
rect 14372 15453 14381 15487
rect 14381 15453 14415 15487
rect 14415 15453 14424 15487
rect 14372 15444 14424 15453
rect 15752 15444 15804 15496
rect 16120 15444 16172 15496
rect 17408 15512 17460 15564
rect 23572 15691 23624 15700
rect 23572 15657 23581 15691
rect 23581 15657 23615 15691
rect 23615 15657 23624 15691
rect 23572 15648 23624 15657
rect 26148 15648 26200 15700
rect 26976 15691 27028 15700
rect 18512 15580 18564 15632
rect 19984 15580 20036 15632
rect 17960 15512 18012 15564
rect 18144 15444 18196 15496
rect 23296 15580 23348 15632
rect 22652 15512 22704 15564
rect 23112 15512 23164 15564
rect 6920 15308 6972 15360
rect 12440 15351 12492 15360
rect 12440 15317 12449 15351
rect 12449 15317 12483 15351
rect 12483 15317 12492 15351
rect 12440 15308 12492 15317
rect 13176 15351 13228 15360
rect 13176 15317 13185 15351
rect 13185 15317 13219 15351
rect 13219 15317 13228 15351
rect 13176 15308 13228 15317
rect 15936 15376 15988 15428
rect 19064 15376 19116 15428
rect 19432 15419 19484 15428
rect 19432 15385 19441 15419
rect 19441 15385 19475 15419
rect 19475 15385 19484 15419
rect 19432 15376 19484 15385
rect 23204 15487 23256 15496
rect 23204 15453 23213 15487
rect 23213 15453 23247 15487
rect 23247 15453 23256 15487
rect 23204 15444 23256 15453
rect 23756 15555 23808 15564
rect 23756 15521 23765 15555
rect 23765 15521 23799 15555
rect 23799 15521 23808 15555
rect 23756 15512 23808 15521
rect 24032 15555 24084 15564
rect 24032 15521 24041 15555
rect 24041 15521 24075 15555
rect 24075 15521 24084 15555
rect 24032 15512 24084 15521
rect 24676 15512 24728 15564
rect 23940 15487 23992 15496
rect 23940 15453 23949 15487
rect 23949 15453 23983 15487
rect 23983 15453 23992 15487
rect 23940 15444 23992 15453
rect 24124 15376 24176 15428
rect 18144 15308 18196 15360
rect 19524 15308 19576 15360
rect 20076 15351 20128 15360
rect 20076 15317 20085 15351
rect 20085 15317 20119 15351
rect 20119 15317 20128 15351
rect 20076 15308 20128 15317
rect 26240 15512 26292 15564
rect 26148 15308 26200 15360
rect 26976 15657 26985 15691
rect 26985 15657 27019 15691
rect 27019 15657 27028 15691
rect 26976 15648 27028 15657
rect 27344 15648 27396 15700
rect 26516 15623 26568 15632
rect 26516 15589 26525 15623
rect 26525 15589 26559 15623
rect 26559 15589 26568 15623
rect 26516 15580 26568 15589
rect 26792 15580 26844 15632
rect 28172 15580 28224 15632
rect 28356 15580 28408 15632
rect 27712 15512 27764 15564
rect 27252 15487 27304 15496
rect 27252 15453 27261 15487
rect 27261 15453 27295 15487
rect 27295 15453 27304 15487
rect 27252 15444 27304 15453
rect 26516 15308 26568 15360
rect 27160 15351 27212 15360
rect 27160 15317 27169 15351
rect 27169 15317 27203 15351
rect 27203 15317 27212 15351
rect 27160 15308 27212 15317
rect 27252 15308 27304 15360
rect 8032 15206 8084 15258
rect 8096 15206 8148 15258
rect 8160 15206 8212 15258
rect 8224 15206 8276 15258
rect 8288 15206 8340 15258
rect 15115 15206 15167 15258
rect 15179 15206 15231 15258
rect 15243 15206 15295 15258
rect 15307 15206 15359 15258
rect 15371 15206 15423 15258
rect 22198 15206 22250 15258
rect 22262 15206 22314 15258
rect 22326 15206 22378 15258
rect 22390 15206 22442 15258
rect 22454 15206 22506 15258
rect 29281 15206 29333 15258
rect 29345 15206 29397 15258
rect 29409 15206 29461 15258
rect 29473 15206 29525 15258
rect 29537 15206 29589 15258
rect 5724 15104 5776 15156
rect 6644 15104 6696 15156
rect 7472 15104 7524 15156
rect 8668 15104 8720 15156
rect 9404 15104 9456 15156
rect 5448 14968 5500 15020
rect 10416 15104 10468 15156
rect 10968 15147 11020 15156
rect 10968 15113 10977 15147
rect 10977 15113 11011 15147
rect 11011 15113 11020 15147
rect 10968 15104 11020 15113
rect 1400 14900 1452 14952
rect 4068 14943 4120 14952
rect 4068 14909 4077 14943
rect 4077 14909 4111 14943
rect 4111 14909 4120 14943
rect 4068 14900 4120 14909
rect 5540 14900 5592 14952
rect 7932 14968 7984 15020
rect 8392 15011 8444 15020
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 8576 14968 8628 15020
rect 9956 15036 10008 15088
rect 8116 14764 8168 14816
rect 9220 14943 9272 14952
rect 9220 14909 9229 14943
rect 9229 14909 9263 14943
rect 9263 14909 9272 14943
rect 9220 14900 9272 14909
rect 10508 14900 10560 14952
rect 11428 14968 11480 15020
rect 13176 15104 13228 15156
rect 13912 15147 13964 15156
rect 13912 15113 13921 15147
rect 13921 15113 13955 15147
rect 13955 15113 13964 15147
rect 13912 15104 13964 15113
rect 11704 15079 11756 15088
rect 11704 15045 11713 15079
rect 11713 15045 11747 15079
rect 11747 15045 11756 15079
rect 11704 15036 11756 15045
rect 11796 15079 11848 15088
rect 11796 15045 11805 15079
rect 11805 15045 11839 15079
rect 11839 15045 11848 15079
rect 11796 15036 11848 15045
rect 12348 15036 12400 15088
rect 12440 15079 12492 15088
rect 12440 15045 12449 15079
rect 12449 15045 12483 15079
rect 12483 15045 12492 15079
rect 12440 15036 12492 15045
rect 13452 14968 13504 15020
rect 11336 14900 11388 14952
rect 15660 15104 15712 15156
rect 16212 15104 16264 15156
rect 15752 15036 15804 15088
rect 16396 15036 16448 15088
rect 20812 15104 20864 15156
rect 24768 15104 24820 15156
rect 24860 15104 24912 15156
rect 19340 15036 19392 15088
rect 18144 14968 18196 15020
rect 19524 14968 19576 15020
rect 11428 14832 11480 14884
rect 14372 14900 14424 14952
rect 15476 14900 15528 14952
rect 17408 14943 17460 14952
rect 17408 14909 17417 14943
rect 17417 14909 17451 14943
rect 17451 14909 17460 14943
rect 17408 14900 17460 14909
rect 19708 15011 19760 15020
rect 19708 14977 19717 15011
rect 19717 14977 19751 15011
rect 19751 14977 19760 15011
rect 19708 14968 19760 14977
rect 24032 15079 24084 15088
rect 24032 15045 24041 15079
rect 24041 15045 24075 15079
rect 24075 15045 24084 15079
rect 27160 15104 27212 15156
rect 27344 15104 27396 15156
rect 24032 15036 24084 15045
rect 21456 14968 21508 15020
rect 19800 14900 19852 14952
rect 20168 14943 20220 14952
rect 20168 14909 20177 14943
rect 20177 14909 20211 14943
rect 20211 14909 20220 14943
rect 20168 14900 20220 14909
rect 22928 15011 22980 15020
rect 22928 14977 22937 15011
rect 22937 14977 22971 15011
rect 22971 14977 22980 15011
rect 22928 14968 22980 14977
rect 23296 15011 23348 15020
rect 23296 14977 23305 15011
rect 23305 14977 23339 15011
rect 23339 14977 23348 15011
rect 23296 14968 23348 14977
rect 23388 14968 23440 15020
rect 24676 15011 24728 15020
rect 24676 14977 24685 15011
rect 24685 14977 24719 15011
rect 24719 14977 24728 15011
rect 24676 14968 24728 14977
rect 24768 15011 24820 15020
rect 24768 14977 24777 15011
rect 24777 14977 24811 15011
rect 24811 14977 24820 15011
rect 24768 14968 24820 14977
rect 17960 14875 18012 14884
rect 17960 14841 17969 14875
rect 17969 14841 18003 14875
rect 18003 14841 18012 14875
rect 17960 14832 18012 14841
rect 19340 14832 19392 14884
rect 14740 14764 14792 14816
rect 15108 14764 15160 14816
rect 16580 14764 16632 14816
rect 18144 14807 18196 14816
rect 18144 14773 18153 14807
rect 18153 14773 18187 14807
rect 18187 14773 18196 14807
rect 18144 14764 18196 14773
rect 19616 14764 19668 14816
rect 21548 14764 21600 14816
rect 25504 14943 25556 14952
rect 25504 14909 25513 14943
rect 25513 14909 25547 14943
rect 25547 14909 25556 14943
rect 25504 14900 25556 14909
rect 23940 14832 23992 14884
rect 27804 15036 27856 15088
rect 27160 15011 27212 15020
rect 27160 14977 27169 15011
rect 27169 14977 27203 15011
rect 27203 14977 27212 15011
rect 27160 14968 27212 14977
rect 28172 14968 28224 15020
rect 27712 14875 27764 14884
rect 27712 14841 27721 14875
rect 27721 14841 27755 14875
rect 27755 14841 27764 14875
rect 27712 14832 27764 14841
rect 23020 14764 23072 14816
rect 24492 14807 24544 14816
rect 24492 14773 24501 14807
rect 24501 14773 24535 14807
rect 24535 14773 24544 14807
rect 24492 14764 24544 14773
rect 27068 14764 27120 14816
rect 4491 14662 4543 14714
rect 4555 14662 4607 14714
rect 4619 14662 4671 14714
rect 4683 14662 4735 14714
rect 4747 14662 4799 14714
rect 11574 14662 11626 14714
rect 11638 14662 11690 14714
rect 11702 14662 11754 14714
rect 11766 14662 11818 14714
rect 11830 14662 11882 14714
rect 18657 14662 18709 14714
rect 18721 14662 18773 14714
rect 18785 14662 18837 14714
rect 18849 14662 18901 14714
rect 18913 14662 18965 14714
rect 25740 14662 25792 14714
rect 25804 14662 25856 14714
rect 25868 14662 25920 14714
rect 25932 14662 25984 14714
rect 25996 14662 26048 14714
rect 6828 14560 6880 14612
rect 11428 14560 11480 14612
rect 10140 14492 10192 14544
rect 7012 14424 7064 14476
rect 7380 14424 7432 14476
rect 8116 14467 8168 14476
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 8116 14424 8168 14433
rect 11336 14424 11388 14476
rect 12624 14560 12676 14612
rect 15108 14560 15160 14612
rect 15384 14560 15436 14612
rect 15660 14560 15712 14612
rect 13452 14424 13504 14476
rect 16212 14603 16264 14612
rect 16212 14569 16221 14603
rect 16221 14569 16255 14603
rect 16255 14569 16264 14603
rect 16212 14560 16264 14569
rect 18144 14560 18196 14612
rect 19524 14560 19576 14612
rect 19616 14560 19668 14612
rect 20168 14560 20220 14612
rect 23388 14560 23440 14612
rect 23572 14603 23624 14612
rect 23572 14569 23581 14603
rect 23581 14569 23615 14603
rect 23615 14569 23624 14603
rect 23572 14560 23624 14569
rect 24492 14560 24544 14612
rect 26884 14560 26936 14612
rect 19340 14492 19392 14544
rect 7840 14356 7892 14408
rect 9220 14356 9272 14408
rect 10416 14399 10468 14408
rect 10416 14365 10425 14399
rect 10425 14365 10459 14399
rect 10459 14365 10468 14399
rect 10416 14356 10468 14365
rect 7748 14288 7800 14340
rect 10784 14399 10836 14408
rect 10784 14365 10793 14399
rect 10793 14365 10827 14399
rect 10827 14365 10836 14399
rect 10784 14356 10836 14365
rect 11244 14356 11296 14408
rect 12992 14356 13044 14408
rect 14280 14356 14332 14408
rect 14648 14356 14700 14408
rect 15752 14399 15804 14408
rect 15752 14365 15761 14399
rect 15761 14365 15795 14399
rect 15795 14365 15804 14399
rect 15752 14356 15804 14365
rect 10692 14331 10744 14340
rect 10692 14297 10701 14331
rect 10701 14297 10735 14331
rect 10735 14297 10744 14331
rect 10692 14288 10744 14297
rect 11152 14288 11204 14340
rect 16304 14424 16356 14476
rect 16580 14399 16632 14408
rect 16580 14365 16589 14399
rect 16589 14365 16623 14399
rect 16623 14365 16632 14399
rect 16580 14356 16632 14365
rect 18604 14399 18656 14408
rect 18604 14365 18613 14399
rect 18613 14365 18647 14399
rect 18647 14365 18656 14399
rect 18604 14356 18656 14365
rect 19064 14356 19116 14408
rect 19708 14492 19760 14544
rect 19984 14492 20036 14544
rect 17040 14288 17092 14340
rect 10968 14220 11020 14272
rect 11060 14263 11112 14272
rect 11060 14229 11069 14263
rect 11069 14229 11103 14263
rect 11103 14229 11112 14263
rect 11060 14220 11112 14229
rect 14832 14220 14884 14272
rect 16764 14263 16816 14272
rect 16764 14229 16773 14263
rect 16773 14229 16807 14263
rect 16807 14229 16816 14263
rect 16764 14220 16816 14229
rect 18328 14263 18380 14272
rect 18328 14229 18337 14263
rect 18337 14229 18371 14263
rect 18371 14229 18380 14263
rect 18328 14220 18380 14229
rect 19248 14263 19300 14272
rect 19248 14229 19257 14263
rect 19257 14229 19291 14263
rect 19291 14229 19300 14263
rect 19248 14220 19300 14229
rect 19524 14331 19576 14340
rect 19524 14297 19533 14331
rect 19533 14297 19567 14331
rect 19567 14297 19576 14331
rect 19524 14288 19576 14297
rect 19892 14288 19944 14340
rect 19984 14331 20036 14340
rect 19984 14297 19993 14331
rect 19993 14297 20027 14331
rect 20027 14297 20036 14331
rect 19984 14288 20036 14297
rect 20076 14220 20128 14272
rect 20536 14356 20588 14408
rect 22652 14492 22704 14544
rect 21548 14399 21600 14408
rect 21548 14365 21557 14399
rect 21557 14365 21591 14399
rect 21591 14365 21600 14399
rect 21548 14356 21600 14365
rect 21640 14399 21692 14408
rect 21640 14365 21649 14399
rect 21649 14365 21683 14399
rect 21683 14365 21692 14399
rect 21640 14356 21692 14365
rect 22836 14424 22888 14476
rect 23940 14424 23992 14476
rect 24492 14467 24544 14476
rect 24492 14433 24501 14467
rect 24501 14433 24535 14467
rect 24535 14433 24544 14467
rect 24492 14424 24544 14433
rect 28172 14492 28224 14544
rect 27068 14467 27120 14476
rect 27068 14433 27077 14467
rect 27077 14433 27111 14467
rect 27111 14433 27120 14467
rect 27068 14424 27120 14433
rect 21916 14331 21968 14340
rect 21916 14297 21925 14331
rect 21925 14297 21959 14331
rect 21959 14297 21968 14331
rect 21916 14288 21968 14297
rect 22560 14399 22612 14408
rect 22560 14365 22569 14399
rect 22569 14365 22603 14399
rect 22603 14365 22612 14399
rect 22560 14356 22612 14365
rect 22652 14399 22704 14408
rect 22652 14365 22661 14399
rect 22661 14365 22695 14399
rect 22695 14365 22704 14399
rect 22652 14356 22704 14365
rect 22928 14399 22980 14408
rect 22928 14365 22937 14399
rect 22937 14365 22971 14399
rect 22971 14365 22980 14399
rect 22928 14356 22980 14365
rect 23664 14356 23716 14408
rect 25872 14356 25924 14408
rect 23112 14288 23164 14340
rect 23848 14220 23900 14272
rect 23940 14263 23992 14272
rect 23940 14229 23949 14263
rect 23949 14229 23983 14263
rect 23983 14229 23992 14263
rect 23940 14220 23992 14229
rect 25504 14220 25556 14272
rect 28080 14288 28132 14340
rect 8032 14118 8084 14170
rect 8096 14118 8148 14170
rect 8160 14118 8212 14170
rect 8224 14118 8276 14170
rect 8288 14118 8340 14170
rect 15115 14118 15167 14170
rect 15179 14118 15231 14170
rect 15243 14118 15295 14170
rect 15307 14118 15359 14170
rect 15371 14118 15423 14170
rect 22198 14118 22250 14170
rect 22262 14118 22314 14170
rect 22326 14118 22378 14170
rect 22390 14118 22442 14170
rect 22454 14118 22506 14170
rect 29281 14118 29333 14170
rect 29345 14118 29397 14170
rect 29409 14118 29461 14170
rect 29473 14118 29525 14170
rect 29537 14118 29589 14170
rect 6368 14059 6420 14068
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 7840 14016 7892 14068
rect 3240 13948 3292 14000
rect 3516 13948 3568 14000
rect 11980 14016 12032 14068
rect 1400 13880 1452 13932
rect 5724 13880 5776 13932
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 6184 13812 6236 13864
rect 6644 13855 6696 13864
rect 6644 13821 6653 13855
rect 6653 13821 6687 13855
rect 6687 13821 6696 13855
rect 6644 13812 6696 13821
rect 6368 13744 6420 13796
rect 7472 13812 7524 13864
rect 9956 13812 10008 13864
rect 10324 13880 10376 13932
rect 10600 13880 10652 13932
rect 7564 13744 7616 13796
rect 10784 13855 10836 13864
rect 10784 13821 10793 13855
rect 10793 13821 10827 13855
rect 10827 13821 10836 13855
rect 10784 13812 10836 13821
rect 12624 13948 12676 14000
rect 13820 13948 13872 14000
rect 18328 14016 18380 14068
rect 19432 14016 19484 14068
rect 19524 14016 19576 14068
rect 19984 14016 20036 14068
rect 20628 14016 20680 14068
rect 11060 13880 11112 13932
rect 15384 13948 15436 14000
rect 14648 13880 14700 13932
rect 14832 13880 14884 13932
rect 15016 13880 15068 13932
rect 5908 13676 5960 13728
rect 6552 13676 6604 13728
rect 10232 13676 10284 13728
rect 10416 13719 10468 13728
rect 10416 13685 10425 13719
rect 10425 13685 10459 13719
rect 10459 13685 10468 13719
rect 10416 13676 10468 13685
rect 11428 13744 11480 13796
rect 12992 13812 13044 13864
rect 12072 13744 12124 13796
rect 14096 13744 14148 13796
rect 16488 13880 16540 13932
rect 15936 13812 15988 13864
rect 16856 13812 16908 13864
rect 15476 13787 15528 13796
rect 15476 13753 15485 13787
rect 15485 13753 15519 13787
rect 15519 13753 15528 13787
rect 15476 13744 15528 13753
rect 18696 13923 18748 13932
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 19156 13880 19208 13932
rect 19340 13923 19392 13932
rect 19340 13889 19349 13923
rect 19349 13889 19383 13923
rect 19383 13889 19392 13923
rect 19340 13880 19392 13889
rect 22560 14016 22612 14068
rect 23112 14016 23164 14068
rect 23848 14016 23900 14068
rect 25136 14016 25188 14068
rect 23572 13948 23624 14000
rect 24124 13948 24176 14000
rect 19524 13923 19576 13932
rect 19524 13889 19533 13923
rect 19533 13889 19567 13923
rect 19567 13889 19576 13923
rect 19524 13880 19576 13889
rect 19616 13923 19668 13932
rect 19616 13889 19625 13923
rect 19625 13889 19659 13923
rect 19659 13889 19668 13923
rect 19616 13880 19668 13889
rect 19708 13923 19760 13932
rect 19708 13889 19717 13923
rect 19717 13889 19751 13923
rect 19751 13889 19760 13923
rect 19708 13880 19760 13889
rect 19800 13880 19852 13932
rect 20720 13880 20772 13932
rect 20812 13880 20864 13932
rect 23480 13923 23532 13932
rect 23480 13889 23489 13923
rect 23489 13889 23523 13923
rect 23523 13889 23532 13923
rect 24492 13923 24544 13932
rect 23480 13880 23532 13889
rect 24492 13889 24501 13923
rect 24501 13889 24535 13923
rect 24535 13889 24544 13923
rect 24492 13880 24544 13889
rect 25872 13880 25924 13932
rect 28448 13880 28500 13932
rect 17132 13744 17184 13796
rect 18144 13744 18196 13796
rect 22192 13812 22244 13864
rect 16764 13676 16816 13728
rect 18420 13719 18472 13728
rect 18420 13685 18429 13719
rect 18429 13685 18463 13719
rect 18463 13685 18472 13719
rect 18420 13676 18472 13685
rect 19340 13676 19392 13728
rect 20168 13719 20220 13728
rect 20168 13685 20177 13719
rect 20177 13685 20211 13719
rect 20211 13685 20220 13719
rect 20168 13676 20220 13685
rect 21732 13676 21784 13728
rect 24124 13855 24176 13864
rect 24124 13821 24133 13855
rect 24133 13821 24167 13855
rect 24167 13821 24176 13855
rect 24124 13812 24176 13821
rect 26332 13812 26384 13864
rect 28080 13812 28132 13864
rect 25320 13676 25372 13728
rect 26240 13719 26292 13728
rect 26240 13685 26249 13719
rect 26249 13685 26283 13719
rect 26283 13685 26292 13719
rect 26240 13676 26292 13685
rect 4491 13574 4543 13626
rect 4555 13574 4607 13626
rect 4619 13574 4671 13626
rect 4683 13574 4735 13626
rect 4747 13574 4799 13626
rect 11574 13574 11626 13626
rect 11638 13574 11690 13626
rect 11702 13574 11754 13626
rect 11766 13574 11818 13626
rect 11830 13574 11882 13626
rect 18657 13574 18709 13626
rect 18721 13574 18773 13626
rect 18785 13574 18837 13626
rect 18849 13574 18901 13626
rect 18913 13574 18965 13626
rect 25740 13574 25792 13626
rect 25804 13574 25856 13626
rect 25868 13574 25920 13626
rect 25932 13574 25984 13626
rect 25996 13574 26048 13626
rect 1860 13472 1912 13524
rect 6644 13472 6696 13524
rect 13268 13472 13320 13524
rect 6000 13404 6052 13456
rect 6460 13404 6512 13456
rect 9680 13404 9732 13456
rect 9772 13404 9824 13456
rect 12532 13404 12584 13456
rect 16396 13472 16448 13524
rect 18512 13472 18564 13524
rect 15752 13404 15804 13456
rect 17868 13404 17920 13456
rect 19524 13515 19576 13524
rect 19524 13481 19533 13515
rect 19533 13481 19567 13515
rect 19567 13481 19576 13515
rect 19524 13472 19576 13481
rect 20444 13472 20496 13524
rect 22928 13472 22980 13524
rect 25320 13472 25372 13524
rect 29000 13515 29052 13524
rect 29000 13481 29009 13515
rect 29009 13481 29043 13515
rect 29043 13481 29052 13515
rect 29000 13472 29052 13481
rect 3516 13336 3568 13388
rect 3056 13268 3108 13320
rect 7288 13336 7340 13388
rect 6920 13268 6972 13320
rect 7196 13268 7248 13320
rect 3240 13132 3292 13184
rect 7104 13175 7156 13184
rect 7104 13141 7113 13175
rect 7113 13141 7147 13175
rect 7147 13141 7156 13175
rect 7104 13132 7156 13141
rect 7196 13132 7248 13184
rect 7564 13311 7616 13320
rect 7564 13277 7573 13311
rect 7573 13277 7607 13311
rect 7607 13277 7616 13311
rect 7564 13268 7616 13277
rect 8576 13268 8628 13320
rect 7472 13132 7524 13184
rect 13360 13336 13412 13388
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 10324 13268 10376 13320
rect 10508 13311 10560 13320
rect 10508 13277 10518 13311
rect 10518 13277 10552 13311
rect 10552 13277 10560 13311
rect 10508 13268 10560 13277
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 11244 13268 11296 13320
rect 11428 13268 11480 13320
rect 11612 13268 11664 13320
rect 14648 13336 14700 13388
rect 10048 13200 10100 13252
rect 10692 13243 10744 13252
rect 10692 13209 10701 13243
rect 10701 13209 10735 13243
rect 10735 13209 10744 13243
rect 10692 13200 10744 13209
rect 9404 13132 9456 13184
rect 10232 13132 10284 13184
rect 11796 13243 11848 13252
rect 11796 13209 11805 13243
rect 11805 13209 11839 13243
rect 11839 13209 11848 13243
rect 11796 13200 11848 13209
rect 14464 13200 14516 13252
rect 16488 13268 16540 13320
rect 17040 13268 17092 13320
rect 18144 13268 18196 13320
rect 16304 13132 16356 13184
rect 16580 13132 16632 13184
rect 18328 13200 18380 13252
rect 19248 13311 19300 13320
rect 19248 13277 19257 13311
rect 19257 13277 19291 13311
rect 19291 13277 19300 13311
rect 19248 13268 19300 13277
rect 19340 13200 19392 13252
rect 17316 13132 17368 13184
rect 20260 13404 20312 13456
rect 19524 13311 19576 13320
rect 19524 13277 19533 13311
rect 19533 13277 19567 13311
rect 19567 13277 19576 13311
rect 19524 13268 19576 13277
rect 21732 13311 21784 13320
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 22192 13336 22244 13388
rect 22652 13336 22704 13388
rect 25136 13336 25188 13388
rect 26240 13336 26292 13388
rect 23296 13311 23348 13320
rect 23296 13277 23305 13311
rect 23305 13277 23339 13311
rect 23339 13277 23348 13311
rect 23296 13268 23348 13277
rect 23756 13268 23808 13320
rect 19708 13175 19760 13184
rect 19708 13141 19717 13175
rect 19717 13141 19751 13175
rect 19751 13141 19760 13175
rect 19708 13132 19760 13141
rect 21824 13175 21876 13184
rect 21824 13141 21833 13175
rect 21833 13141 21867 13175
rect 21867 13141 21876 13175
rect 21824 13132 21876 13141
rect 8032 13030 8084 13082
rect 8096 13030 8148 13082
rect 8160 13030 8212 13082
rect 8224 13030 8276 13082
rect 8288 13030 8340 13082
rect 15115 13030 15167 13082
rect 15179 13030 15231 13082
rect 15243 13030 15295 13082
rect 15307 13030 15359 13082
rect 15371 13030 15423 13082
rect 22198 13030 22250 13082
rect 22262 13030 22314 13082
rect 22326 13030 22378 13082
rect 22390 13030 22442 13082
rect 22454 13030 22506 13082
rect 29281 13030 29333 13082
rect 29345 13030 29397 13082
rect 29409 13030 29461 13082
rect 29473 13030 29525 13082
rect 29537 13030 29589 13082
rect 1400 12792 1452 12844
rect 5172 12928 5224 12980
rect 3516 12860 3568 12912
rect 7104 12928 7156 12980
rect 7196 12928 7248 12980
rect 6736 12860 6788 12912
rect 3148 12792 3200 12844
rect 2044 12767 2096 12776
rect 2044 12733 2053 12767
rect 2053 12733 2087 12767
rect 2087 12733 2096 12767
rect 2044 12724 2096 12733
rect 4896 12792 4948 12844
rect 6460 12792 6512 12844
rect 6552 12724 6604 12776
rect 10416 12928 10468 12980
rect 10784 12928 10836 12980
rect 11796 12928 11848 12980
rect 13268 12928 13320 12980
rect 9956 12860 10008 12912
rect 11428 12860 11480 12912
rect 14648 12971 14700 12980
rect 14648 12937 14657 12971
rect 14657 12937 14691 12971
rect 14691 12937 14700 12971
rect 14648 12928 14700 12937
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 7564 12835 7616 12844
rect 7564 12801 7573 12835
rect 7573 12801 7607 12835
rect 7607 12801 7616 12835
rect 7564 12792 7616 12801
rect 16488 12860 16540 12912
rect 16580 12860 16632 12912
rect 6000 12656 6052 12708
rect 6276 12656 6328 12708
rect 3884 12588 3936 12640
rect 4252 12631 4304 12640
rect 4252 12597 4261 12631
rect 4261 12597 4295 12631
rect 4295 12597 4304 12631
rect 4252 12588 4304 12597
rect 6184 12631 6236 12640
rect 6184 12597 6193 12631
rect 6193 12597 6227 12631
rect 6227 12597 6236 12631
rect 6184 12588 6236 12597
rect 9220 12767 9272 12776
rect 9220 12733 9229 12767
rect 9229 12733 9263 12767
rect 9263 12733 9272 12767
rect 9220 12724 9272 12733
rect 10048 12724 10100 12776
rect 10232 12724 10284 12776
rect 10508 12724 10560 12776
rect 12348 12792 12400 12844
rect 12624 12835 12676 12844
rect 12624 12801 12633 12835
rect 12633 12801 12667 12835
rect 12667 12801 12676 12835
rect 12624 12792 12676 12801
rect 13820 12792 13872 12844
rect 14372 12835 14424 12844
rect 14372 12801 14381 12835
rect 14381 12801 14415 12835
rect 14415 12801 14424 12835
rect 14372 12792 14424 12801
rect 14464 12835 14516 12844
rect 14464 12801 14473 12835
rect 14473 12801 14507 12835
rect 14507 12801 14516 12835
rect 14464 12792 14516 12801
rect 16120 12792 16172 12844
rect 14004 12724 14056 12776
rect 14648 12724 14700 12776
rect 14740 12767 14792 12776
rect 14740 12733 14749 12767
rect 14749 12733 14783 12767
rect 14783 12733 14792 12767
rect 14740 12724 14792 12733
rect 16580 12724 16632 12776
rect 17408 12860 17460 12912
rect 18420 12928 18472 12980
rect 19616 12928 19668 12980
rect 19984 12928 20036 12980
rect 21640 12928 21692 12980
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 16948 12835 17000 12844
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 17132 12792 17184 12844
rect 20812 12860 20864 12912
rect 10508 12588 10560 12640
rect 11244 12588 11296 12640
rect 12808 12631 12860 12640
rect 12808 12597 12817 12631
rect 12817 12597 12851 12631
rect 12851 12597 12860 12631
rect 12808 12588 12860 12597
rect 13912 12588 13964 12640
rect 14372 12588 14424 12640
rect 16120 12588 16172 12640
rect 17960 12588 18012 12640
rect 20720 12792 20772 12844
rect 21548 12835 21600 12844
rect 21548 12801 21557 12835
rect 21557 12801 21591 12835
rect 21591 12801 21600 12835
rect 21548 12792 21600 12801
rect 21824 12792 21876 12844
rect 20260 12724 20312 12776
rect 22192 12724 22244 12776
rect 22744 12767 22796 12776
rect 22744 12733 22753 12767
rect 22753 12733 22787 12767
rect 22787 12733 22796 12767
rect 22744 12724 22796 12733
rect 22928 12724 22980 12776
rect 23388 12792 23440 12844
rect 22652 12656 22704 12708
rect 21548 12588 21600 12640
rect 21640 12588 21692 12640
rect 23388 12631 23440 12640
rect 23388 12597 23397 12631
rect 23397 12597 23431 12631
rect 23431 12597 23440 12631
rect 23388 12588 23440 12597
rect 4491 12486 4543 12538
rect 4555 12486 4607 12538
rect 4619 12486 4671 12538
rect 4683 12486 4735 12538
rect 4747 12486 4799 12538
rect 11574 12486 11626 12538
rect 11638 12486 11690 12538
rect 11702 12486 11754 12538
rect 11766 12486 11818 12538
rect 11830 12486 11882 12538
rect 18657 12486 18709 12538
rect 18721 12486 18773 12538
rect 18785 12486 18837 12538
rect 18849 12486 18901 12538
rect 18913 12486 18965 12538
rect 25740 12486 25792 12538
rect 25804 12486 25856 12538
rect 25868 12486 25920 12538
rect 25932 12486 25984 12538
rect 25996 12486 26048 12538
rect 2044 12384 2096 12436
rect 6920 12427 6972 12436
rect 6920 12393 6929 12427
rect 6929 12393 6963 12427
rect 6963 12393 6972 12427
rect 6920 12384 6972 12393
rect 7564 12384 7616 12436
rect 10232 12384 10284 12436
rect 12256 12384 12308 12436
rect 4252 12316 4304 12368
rect 3516 12248 3568 12300
rect 4988 12248 5040 12300
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5172 12248 5224 12257
rect 6184 12248 6236 12300
rect 7196 12316 7248 12368
rect 7472 12248 7524 12300
rect 3056 12223 3108 12232
rect 3056 12189 3065 12223
rect 3065 12189 3099 12223
rect 3099 12189 3108 12223
rect 3056 12180 3108 12189
rect 3240 12180 3292 12232
rect 4436 12223 4488 12232
rect 4436 12189 4445 12223
rect 4445 12189 4479 12223
rect 4479 12189 4488 12223
rect 4436 12180 4488 12189
rect 4620 12223 4672 12232
rect 4620 12189 4629 12223
rect 4629 12189 4663 12223
rect 4663 12189 4672 12223
rect 4620 12180 4672 12189
rect 7196 12223 7248 12232
rect 7196 12189 7205 12223
rect 7205 12189 7239 12223
rect 7239 12189 7248 12223
rect 7196 12180 7248 12189
rect 9220 12291 9272 12300
rect 9220 12257 9229 12291
rect 9229 12257 9263 12291
rect 9263 12257 9272 12291
rect 9220 12248 9272 12257
rect 12072 12248 12124 12300
rect 15108 12316 15160 12368
rect 13912 12180 13964 12232
rect 14648 12180 14700 12232
rect 14924 12180 14976 12232
rect 15292 12316 15344 12368
rect 15752 12316 15804 12368
rect 22928 12316 22980 12368
rect 23296 12316 23348 12368
rect 16764 12291 16816 12300
rect 16764 12257 16773 12291
rect 16773 12257 16807 12291
rect 16807 12257 16816 12291
rect 16764 12248 16816 12257
rect 23020 12291 23072 12300
rect 23020 12257 23029 12291
rect 23029 12257 23063 12291
rect 23063 12257 23072 12291
rect 23020 12248 23072 12257
rect 23388 12248 23440 12300
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 16672 12223 16724 12232
rect 16672 12189 16681 12223
rect 16681 12189 16715 12223
rect 16715 12189 16724 12223
rect 16672 12180 16724 12189
rect 19708 12180 19760 12232
rect 22192 12180 22244 12232
rect 5356 12112 5408 12164
rect 3884 12044 3936 12096
rect 5540 12044 5592 12096
rect 6368 12044 6420 12096
rect 7012 12087 7064 12096
rect 7012 12053 7021 12087
rect 7021 12053 7055 12087
rect 7055 12053 7064 12087
rect 7012 12044 7064 12053
rect 9772 12112 9824 12164
rect 10048 12112 10100 12164
rect 10968 12112 11020 12164
rect 12532 12112 12584 12164
rect 13728 12112 13780 12164
rect 9588 12044 9640 12096
rect 9864 12044 9916 12096
rect 16948 12112 17000 12164
rect 22652 12180 22704 12232
rect 23296 12180 23348 12232
rect 23020 12112 23072 12164
rect 23756 12155 23808 12164
rect 23756 12121 23765 12155
rect 23765 12121 23799 12155
rect 23799 12121 23808 12155
rect 23756 12112 23808 12121
rect 16764 12044 16816 12096
rect 19800 12087 19852 12096
rect 19800 12053 19809 12087
rect 19809 12053 19843 12087
rect 19843 12053 19852 12087
rect 19800 12044 19852 12053
rect 22652 12044 22704 12096
rect 22836 12044 22888 12096
rect 23480 12044 23532 12096
rect 23848 12087 23900 12096
rect 23848 12053 23857 12087
rect 23857 12053 23891 12087
rect 23891 12053 23900 12087
rect 23848 12044 23900 12053
rect 24308 12044 24360 12096
rect 8032 11942 8084 11994
rect 8096 11942 8148 11994
rect 8160 11942 8212 11994
rect 8224 11942 8276 11994
rect 8288 11942 8340 11994
rect 15115 11942 15167 11994
rect 15179 11942 15231 11994
rect 15243 11942 15295 11994
rect 15307 11942 15359 11994
rect 15371 11942 15423 11994
rect 22198 11942 22250 11994
rect 22262 11942 22314 11994
rect 22326 11942 22378 11994
rect 22390 11942 22442 11994
rect 22454 11942 22506 11994
rect 29281 11942 29333 11994
rect 29345 11942 29397 11994
rect 29409 11942 29461 11994
rect 29473 11942 29525 11994
rect 29537 11942 29589 11994
rect 4436 11840 4488 11892
rect 4988 11840 5040 11892
rect 7196 11840 7248 11892
rect 7472 11840 7524 11892
rect 10232 11840 10284 11892
rect 3148 11772 3200 11824
rect 940 11704 992 11756
rect 2228 11747 2280 11756
rect 2228 11713 2237 11747
rect 2237 11713 2271 11747
rect 2271 11713 2280 11747
rect 2228 11704 2280 11713
rect 4896 11815 4948 11824
rect 4896 11781 4905 11815
rect 4905 11781 4939 11815
rect 4939 11781 4948 11815
rect 4896 11772 4948 11781
rect 6368 11772 6420 11824
rect 2228 11500 2280 11552
rect 4344 11636 4396 11688
rect 5448 11636 5500 11688
rect 4712 11568 4764 11620
rect 6460 11611 6512 11620
rect 6460 11577 6469 11611
rect 6469 11577 6503 11611
rect 6503 11577 6512 11611
rect 9864 11772 9916 11824
rect 12716 11840 12768 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 14280 11772 14332 11824
rect 19984 11883 20036 11892
rect 19984 11849 19993 11883
rect 19993 11849 20027 11883
rect 20027 11849 20036 11883
rect 19984 11840 20036 11849
rect 23296 11840 23348 11892
rect 21732 11772 21784 11824
rect 7288 11704 7340 11756
rect 12072 11747 12124 11756
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 8944 11636 8996 11688
rect 9772 11636 9824 11688
rect 12992 11636 13044 11688
rect 13728 11704 13780 11756
rect 14096 11747 14148 11756
rect 14096 11713 14105 11747
rect 14105 11713 14139 11747
rect 14139 11713 14148 11747
rect 14096 11704 14148 11713
rect 14648 11704 14700 11756
rect 15476 11704 15528 11756
rect 15752 11704 15804 11756
rect 15844 11636 15896 11688
rect 16304 11747 16356 11756
rect 16304 11713 16313 11747
rect 16313 11713 16347 11747
rect 16347 11713 16356 11747
rect 16304 11704 16356 11713
rect 16396 11636 16448 11688
rect 18052 11636 18104 11688
rect 18512 11747 18564 11756
rect 18512 11713 18521 11747
rect 18521 11713 18555 11747
rect 18555 11713 18564 11747
rect 18512 11704 18564 11713
rect 19340 11747 19392 11756
rect 19340 11713 19349 11747
rect 19349 11713 19383 11747
rect 19383 11713 19392 11747
rect 19340 11704 19392 11713
rect 6460 11568 6512 11577
rect 4252 11500 4304 11552
rect 7196 11543 7248 11552
rect 7196 11509 7205 11543
rect 7205 11509 7239 11543
rect 7239 11509 7248 11543
rect 7196 11500 7248 11509
rect 7380 11500 7432 11552
rect 11152 11500 11204 11552
rect 14280 11543 14332 11552
rect 14280 11509 14289 11543
rect 14289 11509 14323 11543
rect 14323 11509 14332 11543
rect 14280 11500 14332 11509
rect 14740 11500 14792 11552
rect 16120 11500 16172 11552
rect 16672 11568 16724 11620
rect 20352 11704 20404 11756
rect 20076 11568 20128 11620
rect 20260 11568 20312 11620
rect 24124 11772 24176 11824
rect 22100 11704 22152 11756
rect 22560 11747 22612 11756
rect 22560 11713 22569 11747
rect 22569 11713 22603 11747
rect 22603 11713 22612 11747
rect 22560 11704 22612 11713
rect 22652 11704 22704 11756
rect 23296 11704 23348 11756
rect 24032 11704 24084 11756
rect 22560 11568 22612 11620
rect 22928 11636 22980 11688
rect 23664 11636 23716 11688
rect 24308 11636 24360 11688
rect 26700 11568 26752 11620
rect 16948 11500 17000 11552
rect 17592 11543 17644 11552
rect 17592 11509 17601 11543
rect 17601 11509 17635 11543
rect 17635 11509 17644 11543
rect 17592 11500 17644 11509
rect 19432 11500 19484 11552
rect 21456 11500 21508 11552
rect 24124 11543 24176 11552
rect 24124 11509 24133 11543
rect 24133 11509 24167 11543
rect 24167 11509 24176 11543
rect 24124 11500 24176 11509
rect 25596 11500 25648 11552
rect 26240 11500 26292 11552
rect 4491 11398 4543 11450
rect 4555 11398 4607 11450
rect 4619 11398 4671 11450
rect 4683 11398 4735 11450
rect 4747 11398 4799 11450
rect 11574 11398 11626 11450
rect 11638 11398 11690 11450
rect 11702 11398 11754 11450
rect 11766 11398 11818 11450
rect 11830 11398 11882 11450
rect 18657 11398 18709 11450
rect 18721 11398 18773 11450
rect 18785 11398 18837 11450
rect 18849 11398 18901 11450
rect 18913 11398 18965 11450
rect 25740 11398 25792 11450
rect 25804 11398 25856 11450
rect 25868 11398 25920 11450
rect 25932 11398 25984 11450
rect 25996 11398 26048 11450
rect 4160 11296 4212 11348
rect 4344 11339 4396 11348
rect 4344 11305 4353 11339
rect 4353 11305 4387 11339
rect 4387 11305 4396 11339
rect 4344 11296 4396 11305
rect 4896 11296 4948 11348
rect 4252 11228 4304 11280
rect 2228 11160 2280 11212
rect 3148 11092 3200 11144
rect 4068 11160 4120 11212
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 4804 11228 4856 11280
rect 5172 11228 5224 11280
rect 5080 11160 5132 11212
rect 5448 11203 5500 11212
rect 5448 11169 5457 11203
rect 5457 11169 5491 11203
rect 5491 11169 5500 11203
rect 5448 11160 5500 11169
rect 7288 11228 7340 11280
rect 9680 11228 9732 11280
rect 10508 11228 10560 11280
rect 3884 11024 3936 11076
rect 4252 11024 4304 11076
rect 4804 11092 4856 11144
rect 7380 11092 7432 11144
rect 7472 11135 7524 11144
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 7840 11092 7892 11144
rect 10968 11092 11020 11144
rect 17592 11296 17644 11348
rect 18052 11339 18104 11348
rect 18052 11305 18061 11339
rect 18061 11305 18095 11339
rect 18095 11305 18104 11339
rect 18052 11296 18104 11305
rect 19800 11296 19852 11348
rect 21640 11296 21692 11348
rect 21916 11296 21968 11348
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 7104 11024 7156 11076
rect 8944 11024 8996 11076
rect 13636 11024 13688 11076
rect 14372 11024 14424 11076
rect 4620 10956 4672 11008
rect 4712 10956 4764 11008
rect 5908 10956 5960 11008
rect 7656 10956 7708 11008
rect 12440 10956 12492 11008
rect 15936 11067 15988 11076
rect 15936 11033 15945 11067
rect 15945 11033 15979 11067
rect 15979 11033 15988 11067
rect 15936 11024 15988 11033
rect 16580 11160 16632 11212
rect 16948 11160 17000 11212
rect 19524 11228 19576 11280
rect 26700 11339 26752 11348
rect 26700 11305 26709 11339
rect 26709 11305 26743 11339
rect 26743 11305 26752 11339
rect 26700 11296 26752 11305
rect 17868 11092 17920 11144
rect 18420 11092 18472 11144
rect 18696 11135 18748 11144
rect 18696 11101 18705 11135
rect 18705 11101 18739 11135
rect 18739 11101 18748 11135
rect 18696 11092 18748 11101
rect 19248 11092 19300 11144
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 19616 11092 19668 11144
rect 21548 11092 21600 11144
rect 16672 11024 16724 11076
rect 16856 11024 16908 11076
rect 19984 11024 20036 11076
rect 17868 10956 17920 11008
rect 19340 10956 19392 11008
rect 20536 10956 20588 11008
rect 23664 11160 23716 11212
rect 24400 11160 24452 11212
rect 22100 11135 22152 11144
rect 22100 11101 22133 11135
rect 22133 11101 22152 11135
rect 22100 11092 22152 11101
rect 22008 11067 22060 11076
rect 22008 11033 22017 11067
rect 22017 11033 22051 11067
rect 22051 11033 22060 11067
rect 22560 11092 22612 11144
rect 23296 11092 23348 11144
rect 22008 11024 22060 11033
rect 22744 11024 22796 11076
rect 22836 11024 22888 11076
rect 23572 11024 23624 11076
rect 23480 10956 23532 11008
rect 24124 11024 24176 11076
rect 24768 11024 24820 11076
rect 24952 11135 25004 11144
rect 24952 11101 24961 11135
rect 24961 11101 24995 11135
rect 24995 11101 25004 11135
rect 24952 11092 25004 11101
rect 26332 11092 26384 11144
rect 27068 11092 27120 11144
rect 28724 11135 28776 11144
rect 28724 11101 28733 11135
rect 28733 11101 28767 11135
rect 28767 11101 28776 11135
rect 28724 11092 28776 11101
rect 25228 11067 25280 11076
rect 25228 11033 25237 11067
rect 25237 11033 25271 11067
rect 25271 11033 25280 11067
rect 25228 11024 25280 11033
rect 26056 10956 26108 11008
rect 29092 11067 29144 11076
rect 29092 11033 29101 11067
rect 29101 11033 29135 11067
rect 29135 11033 29144 11067
rect 29092 11024 29144 11033
rect 8032 10854 8084 10906
rect 8096 10854 8148 10906
rect 8160 10854 8212 10906
rect 8224 10854 8276 10906
rect 8288 10854 8340 10906
rect 15115 10854 15167 10906
rect 15179 10854 15231 10906
rect 15243 10854 15295 10906
rect 15307 10854 15359 10906
rect 15371 10854 15423 10906
rect 22198 10854 22250 10906
rect 22262 10854 22314 10906
rect 22326 10854 22378 10906
rect 22390 10854 22442 10906
rect 22454 10854 22506 10906
rect 29281 10854 29333 10906
rect 29345 10854 29397 10906
rect 29409 10854 29461 10906
rect 29473 10854 29525 10906
rect 29537 10854 29589 10906
rect 4160 10752 4212 10804
rect 5908 10795 5960 10804
rect 5908 10761 5917 10795
rect 5917 10761 5951 10795
rect 5951 10761 5960 10795
rect 5908 10752 5960 10761
rect 6460 10752 6512 10804
rect 4804 10727 4856 10736
rect 4804 10693 4813 10727
rect 4813 10693 4847 10727
rect 4847 10693 4856 10727
rect 4804 10684 4856 10693
rect 3976 10548 4028 10600
rect 4068 10412 4120 10464
rect 4160 10412 4212 10464
rect 4712 10616 4764 10668
rect 4620 10480 4672 10532
rect 5356 10684 5408 10736
rect 5540 10684 5592 10736
rect 7656 10684 7708 10736
rect 9772 10752 9824 10804
rect 9956 10752 10008 10804
rect 14096 10752 14148 10804
rect 14740 10752 14792 10804
rect 18512 10752 18564 10804
rect 21456 10795 21508 10804
rect 21456 10761 21465 10795
rect 21465 10761 21499 10795
rect 21499 10761 21508 10795
rect 21456 10752 21508 10761
rect 22008 10752 22060 10804
rect 23020 10752 23072 10804
rect 7196 10616 7248 10668
rect 9772 10616 9824 10668
rect 5264 10548 5316 10600
rect 4988 10480 5040 10532
rect 7012 10548 7064 10600
rect 10140 10659 10192 10668
rect 10140 10625 10149 10659
rect 10149 10625 10183 10659
rect 10183 10625 10192 10659
rect 10140 10616 10192 10625
rect 10324 10659 10376 10668
rect 10324 10625 10351 10659
rect 10351 10625 10376 10659
rect 10508 10727 10560 10736
rect 10508 10693 10515 10727
rect 10515 10693 10549 10727
rect 10549 10693 10560 10727
rect 10508 10684 10560 10693
rect 11152 10684 11204 10736
rect 19892 10684 19944 10736
rect 10324 10616 10376 10625
rect 13636 10616 13688 10668
rect 14280 10616 14332 10668
rect 14372 10659 14424 10668
rect 14372 10625 14381 10659
rect 14381 10625 14415 10659
rect 14415 10625 14424 10659
rect 14372 10616 14424 10625
rect 16396 10616 16448 10668
rect 10508 10548 10560 10600
rect 11428 10548 11480 10600
rect 12440 10548 12492 10600
rect 10600 10480 10652 10532
rect 14096 10548 14148 10600
rect 15936 10548 15988 10600
rect 17316 10659 17368 10668
rect 17316 10625 17330 10659
rect 17330 10625 17364 10659
rect 17364 10625 17368 10659
rect 17316 10616 17368 10625
rect 17684 10616 17736 10668
rect 17868 10659 17920 10668
rect 17868 10625 17874 10659
rect 17874 10625 17908 10659
rect 17908 10625 17920 10659
rect 17868 10616 17920 10625
rect 18052 10616 18104 10668
rect 18328 10659 18380 10668
rect 18328 10625 18337 10659
rect 18337 10625 18371 10659
rect 18371 10625 18380 10659
rect 18328 10616 18380 10625
rect 18696 10616 18748 10668
rect 19156 10659 19208 10668
rect 19156 10625 19165 10659
rect 19165 10625 19199 10659
rect 19199 10625 19208 10659
rect 19156 10616 19208 10625
rect 20076 10684 20128 10736
rect 23848 10752 23900 10804
rect 25228 10752 25280 10804
rect 20260 10616 20312 10668
rect 22100 10659 22152 10668
rect 10232 10412 10284 10464
rect 10508 10412 10560 10464
rect 13544 10455 13596 10464
rect 13544 10421 13553 10455
rect 13553 10421 13587 10455
rect 13587 10421 13596 10455
rect 13544 10412 13596 10421
rect 15292 10480 15344 10532
rect 20352 10548 20404 10600
rect 22100 10625 22109 10659
rect 22109 10625 22143 10659
rect 22143 10625 22152 10659
rect 22100 10616 22152 10625
rect 24400 10684 24452 10736
rect 26056 10727 26108 10736
rect 26056 10693 26065 10727
rect 26065 10693 26099 10727
rect 26099 10693 26108 10727
rect 26056 10684 26108 10693
rect 26240 10684 26292 10736
rect 14464 10412 14516 10464
rect 15660 10412 15712 10464
rect 16396 10412 16448 10464
rect 16948 10412 17000 10464
rect 22652 10548 22704 10600
rect 26424 10659 26476 10668
rect 26424 10625 26433 10659
rect 26433 10625 26467 10659
rect 26467 10625 26476 10659
rect 26424 10616 26476 10625
rect 26516 10659 26568 10668
rect 26516 10625 26525 10659
rect 26525 10625 26559 10659
rect 26559 10625 26568 10659
rect 26516 10616 26568 10625
rect 22836 10480 22888 10532
rect 18052 10412 18104 10464
rect 19064 10412 19116 10464
rect 20260 10412 20312 10464
rect 22100 10412 22152 10464
rect 22376 10412 22428 10464
rect 22560 10455 22612 10464
rect 22560 10421 22569 10455
rect 22569 10421 22603 10455
rect 22603 10421 22612 10455
rect 22560 10412 22612 10421
rect 22652 10412 22704 10464
rect 23664 10548 23716 10600
rect 25596 10591 25648 10600
rect 25596 10557 25605 10591
rect 25605 10557 25639 10591
rect 25639 10557 25648 10591
rect 25596 10548 25648 10557
rect 25872 10548 25924 10600
rect 26148 10548 26200 10600
rect 24768 10480 24820 10532
rect 22928 10412 22980 10464
rect 24952 10412 25004 10464
rect 4491 10310 4543 10362
rect 4555 10310 4607 10362
rect 4619 10310 4671 10362
rect 4683 10310 4735 10362
rect 4747 10310 4799 10362
rect 11574 10310 11626 10362
rect 11638 10310 11690 10362
rect 11702 10310 11754 10362
rect 11766 10310 11818 10362
rect 11830 10310 11882 10362
rect 18657 10310 18709 10362
rect 18721 10310 18773 10362
rect 18785 10310 18837 10362
rect 18849 10310 18901 10362
rect 18913 10310 18965 10362
rect 25740 10310 25792 10362
rect 25804 10310 25856 10362
rect 25868 10310 25920 10362
rect 25932 10310 25984 10362
rect 25996 10310 26048 10362
rect 4068 10208 4120 10260
rect 9772 10208 9824 10260
rect 10140 10208 10192 10260
rect 12348 10208 12400 10260
rect 13544 10251 13596 10260
rect 13544 10217 13553 10251
rect 13553 10217 13587 10251
rect 13587 10217 13596 10251
rect 13544 10208 13596 10217
rect 13912 10208 13964 10260
rect 3976 10140 4028 10192
rect 5264 10140 5316 10192
rect 10968 10140 11020 10192
rect 18052 10208 18104 10260
rect 20536 10251 20588 10260
rect 20536 10217 20545 10251
rect 20545 10217 20579 10251
rect 20579 10217 20588 10251
rect 20536 10208 20588 10217
rect 22100 10208 22152 10260
rect 22652 10208 22704 10260
rect 9588 10115 9640 10124
rect 9588 10081 9597 10115
rect 9597 10081 9631 10115
rect 9631 10081 9640 10115
rect 9588 10072 9640 10081
rect 9772 10072 9824 10124
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 9956 10004 10008 10056
rect 10232 10115 10284 10124
rect 10232 10081 10241 10115
rect 10241 10081 10275 10115
rect 10275 10081 10284 10115
rect 10232 10072 10284 10081
rect 10324 10004 10376 10056
rect 10784 10004 10836 10056
rect 10968 10004 11020 10056
rect 11060 10004 11112 10056
rect 11244 10047 11296 10056
rect 11244 10013 11253 10047
rect 11253 10013 11287 10047
rect 11287 10013 11296 10047
rect 11244 10004 11296 10013
rect 11428 10047 11480 10056
rect 11428 10013 11437 10047
rect 11437 10013 11471 10047
rect 11471 10013 11480 10047
rect 11428 10004 11480 10013
rect 16580 10115 16632 10124
rect 16580 10081 16589 10115
rect 16589 10081 16623 10115
rect 16623 10081 16632 10115
rect 16580 10072 16632 10081
rect 18420 10140 18472 10192
rect 19156 10072 19208 10124
rect 22376 10140 22428 10192
rect 22560 10140 22612 10192
rect 23112 10208 23164 10260
rect 23204 10208 23256 10260
rect 25596 10208 25648 10260
rect 20260 10072 20312 10124
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 13912 10004 13964 10056
rect 15384 10047 15436 10056
rect 15384 10013 15393 10047
rect 15393 10013 15427 10047
rect 15427 10013 15436 10047
rect 15384 10004 15436 10013
rect 13360 9979 13412 9988
rect 13360 9945 13369 9979
rect 13369 9945 13403 9979
rect 13403 9945 13412 9979
rect 13360 9936 13412 9945
rect 15292 9936 15344 9988
rect 9036 9911 9088 9920
rect 9036 9877 9045 9911
rect 9045 9877 9079 9911
rect 9079 9877 9088 9911
rect 9036 9868 9088 9877
rect 9864 9868 9916 9920
rect 10416 9868 10468 9920
rect 10692 9911 10744 9920
rect 10692 9877 10701 9911
rect 10701 9877 10735 9911
rect 10735 9877 10744 9911
rect 10692 9868 10744 9877
rect 11152 9868 11204 9920
rect 11980 9868 12032 9920
rect 13084 9868 13136 9920
rect 13820 9868 13872 9920
rect 14372 9868 14424 9920
rect 15660 10047 15712 10056
rect 15660 10013 15669 10047
rect 15669 10013 15703 10047
rect 15703 10013 15712 10047
rect 15660 10004 15712 10013
rect 16304 10004 16356 10056
rect 17960 10004 18012 10056
rect 18328 10004 18380 10056
rect 20076 10004 20128 10056
rect 20352 10004 20404 10056
rect 21640 10004 21692 10056
rect 15568 9868 15620 9920
rect 16856 9979 16908 9988
rect 16856 9945 16865 9979
rect 16865 9945 16899 9979
rect 16899 9945 16908 9979
rect 16856 9936 16908 9945
rect 22652 10004 22704 10056
rect 23112 10047 23164 10056
rect 23112 10013 23121 10047
rect 23121 10013 23155 10047
rect 23155 10013 23164 10047
rect 23112 10004 23164 10013
rect 26424 10004 26476 10056
rect 22560 9936 22612 9988
rect 22836 9979 22888 9988
rect 22836 9945 22845 9979
rect 22845 9945 22879 9979
rect 22879 9945 22888 9979
rect 22836 9936 22888 9945
rect 26240 9936 26292 9988
rect 18328 9911 18380 9920
rect 18328 9877 18337 9911
rect 18337 9877 18371 9911
rect 18371 9877 18380 9911
rect 18328 9868 18380 9877
rect 19064 9911 19116 9920
rect 19064 9877 19073 9911
rect 19073 9877 19107 9911
rect 19107 9877 19116 9911
rect 19064 9868 19116 9877
rect 22100 9868 22152 9920
rect 26516 9868 26568 9920
rect 8032 9766 8084 9818
rect 8096 9766 8148 9818
rect 8160 9766 8212 9818
rect 8224 9766 8276 9818
rect 8288 9766 8340 9818
rect 15115 9766 15167 9818
rect 15179 9766 15231 9818
rect 15243 9766 15295 9818
rect 15307 9766 15359 9818
rect 15371 9766 15423 9818
rect 22198 9766 22250 9818
rect 22262 9766 22314 9818
rect 22326 9766 22378 9818
rect 22390 9766 22442 9818
rect 22454 9766 22506 9818
rect 29281 9766 29333 9818
rect 29345 9766 29397 9818
rect 29409 9766 29461 9818
rect 29473 9766 29525 9818
rect 29537 9766 29589 9818
rect 6552 9664 6604 9716
rect 2228 9596 2280 9648
rect 4068 9596 4120 9648
rect 6276 9596 6328 9648
rect 9956 9664 10008 9716
rect 10508 9664 10560 9716
rect 10600 9707 10652 9716
rect 10600 9673 10609 9707
rect 10609 9673 10643 9707
rect 10643 9673 10652 9707
rect 10600 9664 10652 9673
rect 3332 9528 3384 9580
rect 3792 9528 3844 9580
rect 5172 9528 5224 9580
rect 4160 9460 4212 9512
rect 5540 9528 5592 9580
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 10232 9639 10284 9648
rect 10232 9605 10241 9639
rect 10241 9605 10275 9639
rect 10275 9605 10284 9639
rect 10232 9596 10284 9605
rect 10692 9596 10744 9648
rect 10968 9664 11020 9716
rect 16856 9664 16908 9716
rect 18512 9707 18564 9716
rect 18512 9673 18521 9707
rect 18521 9673 18555 9707
rect 18555 9673 18564 9707
rect 18512 9664 18564 9673
rect 21732 9664 21784 9716
rect 9036 9528 9088 9580
rect 9864 9528 9916 9580
rect 4344 9324 4396 9376
rect 4988 9392 5040 9444
rect 5908 9392 5960 9444
rect 5080 9324 5132 9376
rect 5632 9367 5684 9376
rect 5632 9333 5641 9367
rect 5641 9333 5675 9367
rect 5675 9333 5684 9367
rect 5632 9324 5684 9333
rect 6552 9392 6604 9444
rect 6644 9324 6696 9376
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7196 9324 7248 9333
rect 8852 9503 8904 9512
rect 8852 9469 8861 9503
rect 8861 9469 8895 9503
rect 8895 9469 8904 9503
rect 8852 9460 8904 9469
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 9680 9460 9732 9512
rect 9772 9503 9824 9512
rect 9772 9469 9781 9503
rect 9781 9469 9815 9503
rect 9815 9469 9824 9503
rect 9772 9460 9824 9469
rect 10416 9460 10468 9512
rect 10232 9392 10284 9444
rect 11336 9596 11388 9648
rect 13176 9639 13228 9648
rect 13176 9605 13185 9639
rect 13185 9605 13219 9639
rect 13219 9605 13228 9639
rect 13176 9596 13228 9605
rect 12348 9528 12400 9580
rect 13452 9596 13504 9648
rect 13820 9596 13872 9648
rect 14280 9596 14332 9648
rect 10692 9503 10744 9512
rect 10692 9469 10701 9503
rect 10701 9469 10735 9503
rect 10735 9469 10744 9503
rect 10692 9460 10744 9469
rect 11060 9460 11112 9512
rect 10508 9324 10560 9376
rect 11428 9324 11480 9376
rect 14096 9460 14148 9512
rect 16764 9460 16816 9512
rect 17040 9571 17092 9580
rect 17040 9537 17049 9571
rect 17049 9537 17083 9571
rect 17083 9537 17092 9571
rect 17040 9528 17092 9537
rect 17868 9528 17920 9580
rect 18052 9528 18104 9580
rect 18328 9528 18380 9580
rect 18420 9571 18472 9580
rect 18420 9537 18462 9571
rect 18462 9537 18472 9571
rect 18420 9528 18472 9537
rect 19064 9528 19116 9580
rect 25596 9596 25648 9648
rect 22652 9528 22704 9580
rect 23388 9528 23440 9580
rect 25504 9528 25556 9580
rect 17132 9392 17184 9444
rect 26884 9460 26936 9512
rect 26148 9392 26200 9444
rect 27896 9392 27948 9444
rect 13728 9324 13780 9376
rect 14280 9324 14332 9376
rect 17592 9367 17644 9376
rect 17592 9333 17601 9367
rect 17601 9333 17635 9367
rect 17635 9333 17644 9367
rect 17592 9324 17644 9333
rect 17960 9324 18012 9376
rect 19340 9324 19392 9376
rect 26608 9324 26660 9376
rect 28172 9571 28224 9580
rect 28172 9537 28181 9571
rect 28181 9537 28215 9571
rect 28215 9537 28224 9571
rect 28172 9528 28224 9537
rect 28080 9460 28132 9512
rect 4491 9222 4543 9274
rect 4555 9222 4607 9274
rect 4619 9222 4671 9274
rect 4683 9222 4735 9274
rect 4747 9222 4799 9274
rect 11574 9222 11626 9274
rect 11638 9222 11690 9274
rect 11702 9222 11754 9274
rect 11766 9222 11818 9274
rect 11830 9222 11882 9274
rect 18657 9222 18709 9274
rect 18721 9222 18773 9274
rect 18785 9222 18837 9274
rect 18849 9222 18901 9274
rect 18913 9222 18965 9274
rect 25740 9222 25792 9274
rect 25804 9222 25856 9274
rect 25868 9222 25920 9274
rect 25932 9222 25984 9274
rect 25996 9222 26048 9274
rect 5632 9120 5684 9172
rect 4160 9052 4212 9104
rect 4988 9052 5040 9104
rect 5448 9052 5500 9104
rect 10232 9052 10284 9104
rect 13084 9163 13136 9172
rect 13084 9129 13093 9163
rect 13093 9129 13127 9163
rect 13127 9129 13136 9163
rect 13084 9120 13136 9129
rect 17500 9120 17552 9172
rect 2228 8984 2280 9036
rect 4344 8984 4396 9036
rect 9128 8984 9180 9036
rect 9864 8984 9916 9036
rect 10140 8984 10192 9036
rect 3792 8848 3844 8900
rect 6000 8916 6052 8968
rect 6460 8916 6512 8968
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 10784 8984 10836 9036
rect 11152 9027 11204 9036
rect 11152 8993 11161 9027
rect 11161 8993 11195 9027
rect 11195 8993 11204 9027
rect 11152 8984 11204 8993
rect 17316 9052 17368 9104
rect 22836 9120 22888 9172
rect 26884 9120 26936 9172
rect 24032 9052 24084 9104
rect 11980 8984 12032 9036
rect 15752 8984 15804 9036
rect 16672 8984 16724 9036
rect 6276 8848 6328 8900
rect 7104 8848 7156 8900
rect 10048 8848 10100 8900
rect 11336 8848 11388 8900
rect 4344 8780 4396 8832
rect 6092 8823 6144 8832
rect 6092 8789 6101 8823
rect 6101 8789 6135 8823
rect 6135 8789 6144 8823
rect 6092 8780 6144 8789
rect 9956 8780 10008 8832
rect 12256 8916 12308 8968
rect 13728 8916 13780 8968
rect 22376 9027 22428 9036
rect 22376 8993 22385 9027
rect 22385 8993 22419 9027
rect 22419 8993 22428 9027
rect 22376 8984 22428 8993
rect 22560 8984 22612 9036
rect 22652 9027 22704 9036
rect 22652 8993 22661 9027
rect 22661 8993 22695 9027
rect 22695 8993 22704 9027
rect 22652 8984 22704 8993
rect 13268 8848 13320 8900
rect 13912 8848 13964 8900
rect 13636 8823 13688 8832
rect 13636 8789 13651 8823
rect 13651 8789 13685 8823
rect 13685 8789 13688 8823
rect 13636 8780 13688 8789
rect 18328 8959 18380 8968
rect 18328 8925 18337 8959
rect 18337 8925 18371 8959
rect 18371 8925 18380 8959
rect 18328 8916 18380 8925
rect 19340 8959 19392 8968
rect 19340 8925 19349 8959
rect 19349 8925 19383 8959
rect 19383 8925 19392 8959
rect 19340 8916 19392 8925
rect 18236 8891 18288 8900
rect 18236 8857 18241 8891
rect 18241 8857 18275 8891
rect 18275 8857 18288 8891
rect 18236 8848 18288 8857
rect 22100 8959 22152 8968
rect 22100 8925 22109 8959
rect 22109 8925 22143 8959
rect 22143 8925 22152 8959
rect 22100 8916 22152 8925
rect 27252 8984 27304 9036
rect 22836 8959 22888 8968
rect 22836 8925 22845 8959
rect 22845 8925 22879 8959
rect 22879 8925 22888 8959
rect 22836 8916 22888 8925
rect 24952 8916 25004 8968
rect 25596 8916 25648 8968
rect 26148 8959 26200 8968
rect 26148 8925 26157 8959
rect 26157 8925 26191 8959
rect 26191 8925 26200 8959
rect 26148 8916 26200 8925
rect 27896 8916 27948 8968
rect 23388 8848 23440 8900
rect 25780 8891 25832 8900
rect 25780 8857 25789 8891
rect 25789 8857 25823 8891
rect 25823 8857 25832 8891
rect 25780 8848 25832 8857
rect 25872 8891 25924 8900
rect 25872 8857 25881 8891
rect 25881 8857 25915 8891
rect 25915 8857 25924 8891
rect 25872 8848 25924 8857
rect 26240 8848 26292 8900
rect 26424 8848 26476 8900
rect 18512 8823 18564 8832
rect 18512 8789 18521 8823
rect 18521 8789 18555 8823
rect 18555 8789 18564 8823
rect 18512 8780 18564 8789
rect 20628 8780 20680 8832
rect 21732 8823 21784 8832
rect 21732 8789 21741 8823
rect 21741 8789 21775 8823
rect 21775 8789 21784 8823
rect 21732 8780 21784 8789
rect 22100 8780 22152 8832
rect 22376 8780 22428 8832
rect 24308 8780 24360 8832
rect 27068 8848 27120 8900
rect 27804 8848 27856 8900
rect 8032 8678 8084 8730
rect 8096 8678 8148 8730
rect 8160 8678 8212 8730
rect 8224 8678 8276 8730
rect 8288 8678 8340 8730
rect 15115 8678 15167 8730
rect 15179 8678 15231 8730
rect 15243 8678 15295 8730
rect 15307 8678 15359 8730
rect 15371 8678 15423 8730
rect 22198 8678 22250 8730
rect 22262 8678 22314 8730
rect 22326 8678 22378 8730
rect 22390 8678 22442 8730
rect 22454 8678 22506 8730
rect 29281 8678 29333 8730
rect 29345 8678 29397 8730
rect 29409 8678 29461 8730
rect 29473 8678 29525 8730
rect 29537 8678 29589 8730
rect 2228 8576 2280 8628
rect 4160 8576 4212 8628
rect 5448 8619 5500 8628
rect 5448 8585 5457 8619
rect 5457 8585 5491 8619
rect 5491 8585 5500 8619
rect 5448 8576 5500 8585
rect 1676 8440 1728 8492
rect 2688 8508 2740 8560
rect 3792 8440 3844 8492
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 4804 8440 4856 8492
rect 6092 8576 6144 8628
rect 6460 8576 6512 8628
rect 6736 8576 6788 8628
rect 5816 8508 5868 8560
rect 6000 8508 6052 8560
rect 5448 8440 5500 8492
rect 4344 8304 4396 8356
rect 5080 8372 5132 8424
rect 5908 8415 5960 8424
rect 5908 8381 5917 8415
rect 5917 8381 5951 8415
rect 5951 8381 5960 8415
rect 5908 8372 5960 8381
rect 6000 8415 6052 8424
rect 6000 8381 6009 8415
rect 6009 8381 6043 8415
rect 6043 8381 6052 8415
rect 6000 8372 6052 8381
rect 6276 8440 6328 8492
rect 6828 8483 6880 8492
rect 6828 8449 6837 8483
rect 6837 8449 6871 8483
rect 6871 8449 6880 8483
rect 6828 8440 6880 8449
rect 9036 8551 9088 8560
rect 9036 8517 9045 8551
rect 9045 8517 9079 8551
rect 9079 8517 9088 8551
rect 9036 8508 9088 8517
rect 9956 8576 10008 8628
rect 13268 8576 13320 8628
rect 9680 8440 9732 8492
rect 10508 8440 10560 8492
rect 13636 8508 13688 8560
rect 14280 8508 14332 8560
rect 16580 8576 16632 8628
rect 17592 8576 17644 8628
rect 18512 8576 18564 8628
rect 20628 8619 20680 8628
rect 20628 8585 20637 8619
rect 20637 8585 20671 8619
rect 20671 8585 20680 8619
rect 20628 8576 20680 8585
rect 21732 8576 21784 8628
rect 22836 8576 22888 8628
rect 26240 8576 26292 8628
rect 15752 8508 15804 8560
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 17500 8483 17552 8492
rect 17500 8449 17509 8483
rect 17509 8449 17543 8483
rect 17543 8449 17552 8483
rect 17500 8440 17552 8449
rect 17684 8440 17736 8492
rect 6644 8415 6696 8424
rect 6644 8381 6653 8415
rect 6653 8381 6687 8415
rect 6687 8381 6696 8415
rect 6644 8372 6696 8381
rect 6736 8415 6788 8424
rect 6736 8381 6745 8415
rect 6745 8381 6779 8415
rect 6779 8381 6788 8415
rect 6736 8372 6788 8381
rect 7932 8372 7984 8424
rect 5264 8279 5316 8288
rect 5264 8245 5273 8279
rect 5273 8245 5307 8279
rect 5307 8245 5316 8279
rect 5264 8236 5316 8245
rect 5540 8236 5592 8288
rect 6184 8236 6236 8288
rect 9588 8372 9640 8424
rect 13360 8415 13412 8424
rect 13360 8381 13369 8415
rect 13369 8381 13403 8415
rect 13403 8381 13412 8415
rect 13360 8372 13412 8381
rect 13452 8415 13504 8424
rect 13452 8381 13461 8415
rect 13461 8381 13495 8415
rect 13495 8381 13504 8415
rect 13452 8372 13504 8381
rect 14096 8372 14148 8424
rect 19248 8508 19300 8560
rect 12716 8304 12768 8356
rect 18236 8304 18288 8356
rect 23572 8508 23624 8560
rect 25780 8508 25832 8560
rect 26332 8508 26384 8560
rect 22560 8440 22612 8492
rect 23020 8483 23072 8492
rect 23020 8449 23029 8483
rect 23029 8449 23063 8483
rect 23063 8449 23072 8483
rect 23020 8440 23072 8449
rect 23296 8440 23348 8492
rect 23480 8483 23532 8492
rect 23480 8449 23489 8483
rect 23489 8449 23523 8483
rect 23523 8449 23532 8483
rect 23480 8440 23532 8449
rect 23112 8372 23164 8424
rect 23388 8372 23440 8424
rect 23756 8415 23808 8424
rect 23756 8381 23765 8415
rect 23765 8381 23799 8415
rect 23799 8381 23808 8415
rect 23756 8372 23808 8381
rect 24032 8440 24084 8492
rect 24584 8372 24636 8424
rect 13912 8236 13964 8288
rect 16396 8236 16448 8288
rect 17776 8279 17828 8288
rect 17776 8245 17785 8279
rect 17785 8245 17819 8279
rect 17819 8245 17828 8279
rect 17776 8236 17828 8245
rect 23664 8347 23716 8356
rect 23664 8313 23673 8347
rect 23673 8313 23707 8347
rect 23707 8313 23716 8347
rect 23664 8304 23716 8313
rect 25504 8440 25556 8492
rect 26148 8440 26200 8492
rect 26608 8440 26660 8492
rect 27252 8483 27304 8492
rect 27252 8449 27261 8483
rect 27261 8449 27295 8483
rect 27295 8449 27304 8483
rect 27252 8440 27304 8449
rect 28172 8576 28224 8628
rect 28080 8508 28132 8560
rect 26240 8372 26292 8424
rect 27528 8372 27580 8424
rect 25228 8304 25280 8356
rect 26608 8347 26660 8356
rect 26608 8313 26617 8347
rect 26617 8313 26651 8347
rect 26651 8313 26660 8347
rect 26608 8304 26660 8313
rect 20812 8236 20864 8288
rect 20904 8279 20956 8288
rect 20904 8245 20913 8279
rect 20913 8245 20947 8279
rect 20947 8245 20956 8279
rect 20904 8236 20956 8245
rect 22468 8236 22520 8288
rect 22928 8236 22980 8288
rect 24676 8236 24728 8288
rect 27344 8236 27396 8288
rect 4491 8134 4543 8186
rect 4555 8134 4607 8186
rect 4619 8134 4671 8186
rect 4683 8134 4735 8186
rect 4747 8134 4799 8186
rect 11574 8134 11626 8186
rect 11638 8134 11690 8186
rect 11702 8134 11754 8186
rect 11766 8134 11818 8186
rect 11830 8134 11882 8186
rect 18657 8134 18709 8186
rect 18721 8134 18773 8186
rect 18785 8134 18837 8186
rect 18849 8134 18901 8186
rect 18913 8134 18965 8186
rect 25740 8134 25792 8186
rect 25804 8134 25856 8186
rect 25868 8134 25920 8186
rect 25932 8134 25984 8186
rect 25996 8134 26048 8186
rect 4068 7964 4120 8016
rect 6736 8007 6788 8016
rect 6736 7973 6745 8007
rect 6745 7973 6779 8007
rect 6779 7973 6788 8007
rect 6736 7964 6788 7973
rect 14004 8032 14056 8084
rect 14188 7964 14240 8016
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 5448 7896 5500 7948
rect 6000 7896 6052 7948
rect 7196 7896 7248 7948
rect 12808 7896 12860 7948
rect 17408 8032 17460 8084
rect 16580 7964 16632 8016
rect 3792 7760 3844 7812
rect 4988 7871 5040 7880
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 4252 7760 4304 7812
rect 4896 7803 4948 7812
rect 4896 7769 4905 7803
rect 4905 7769 4939 7803
rect 4939 7769 4948 7803
rect 4896 7760 4948 7769
rect 5172 7760 5224 7812
rect 6184 7760 6236 7812
rect 14004 7828 14056 7880
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 6828 7760 6880 7812
rect 13636 7760 13688 7812
rect 13728 7803 13780 7812
rect 13728 7769 13769 7803
rect 13769 7769 13780 7803
rect 14372 7828 14424 7880
rect 13728 7760 13780 7769
rect 7196 7735 7248 7744
rect 7196 7701 7205 7735
rect 7205 7701 7239 7735
rect 7239 7701 7248 7735
rect 7196 7692 7248 7701
rect 13360 7692 13412 7744
rect 14648 7828 14700 7880
rect 15016 7828 15068 7880
rect 15476 7828 15528 7880
rect 16396 7871 16448 7880
rect 16396 7837 16405 7871
rect 16405 7837 16439 7871
rect 16439 7837 16448 7871
rect 16396 7828 16448 7837
rect 16580 7871 16632 7880
rect 16580 7837 16589 7871
rect 16589 7837 16623 7871
rect 16623 7837 16632 7871
rect 16580 7828 16632 7837
rect 17316 7828 17368 7880
rect 17408 7871 17460 7880
rect 17408 7837 17417 7871
rect 17417 7837 17451 7871
rect 17451 7837 17460 7871
rect 17408 7828 17460 7837
rect 17684 8032 17736 8084
rect 17592 7964 17644 8016
rect 17224 7803 17276 7812
rect 17224 7769 17233 7803
rect 17233 7769 17267 7803
rect 17267 7769 17276 7803
rect 17224 7760 17276 7769
rect 13912 7735 13964 7744
rect 13912 7701 13921 7735
rect 13921 7701 13955 7735
rect 13955 7701 13964 7735
rect 13912 7692 13964 7701
rect 14464 7735 14516 7744
rect 14464 7701 14473 7735
rect 14473 7701 14507 7735
rect 14507 7701 14516 7735
rect 14464 7692 14516 7701
rect 14648 7735 14700 7744
rect 14648 7701 14657 7735
rect 14657 7701 14691 7735
rect 14691 7701 14700 7735
rect 14648 7692 14700 7701
rect 16764 7735 16816 7744
rect 16764 7701 16773 7735
rect 16773 7701 16807 7735
rect 16807 7701 16816 7735
rect 17960 7871 18012 7880
rect 17960 7837 17967 7871
rect 17967 7837 18012 7871
rect 17960 7828 18012 7837
rect 22100 8032 22152 8084
rect 22192 8032 22244 8084
rect 23480 8032 23532 8084
rect 25228 8075 25280 8084
rect 25228 8041 25237 8075
rect 25237 8041 25271 8075
rect 25271 8041 25280 8075
rect 25228 8032 25280 8041
rect 20904 7896 20956 7948
rect 20076 7871 20128 7880
rect 20076 7837 20085 7871
rect 20085 7837 20119 7871
rect 20119 7837 20128 7871
rect 20076 7828 20128 7837
rect 22284 7871 22336 7880
rect 20812 7760 20864 7812
rect 22284 7837 22293 7871
rect 22293 7837 22327 7871
rect 22327 7837 22336 7871
rect 22284 7828 22336 7837
rect 22468 7896 22520 7948
rect 22560 7871 22612 7880
rect 22560 7837 22569 7871
rect 22569 7837 22603 7871
rect 22603 7837 22612 7871
rect 22560 7828 22612 7837
rect 22836 7828 22888 7880
rect 23020 7830 23072 7882
rect 23112 7871 23164 7880
rect 23112 7837 23127 7871
rect 23127 7837 23161 7871
rect 23161 7837 23164 7871
rect 23112 7828 23164 7837
rect 23296 7871 23348 7880
rect 23296 7837 23305 7871
rect 23305 7837 23339 7871
rect 23339 7837 23348 7871
rect 23296 7828 23348 7837
rect 22652 7803 22704 7812
rect 22652 7769 22661 7803
rect 22661 7769 22695 7803
rect 22695 7769 22704 7803
rect 22652 7760 22704 7769
rect 16764 7692 16816 7701
rect 18328 7692 18380 7744
rect 22100 7692 22152 7744
rect 22468 7692 22520 7744
rect 23388 7803 23440 7812
rect 23388 7769 23397 7803
rect 23397 7769 23431 7803
rect 23431 7769 23440 7803
rect 23388 7760 23440 7769
rect 23572 7964 23624 8016
rect 24032 7964 24084 8016
rect 26148 8032 26200 8084
rect 27344 8032 27396 8084
rect 28080 8032 28132 8084
rect 23572 7828 23624 7880
rect 23664 7871 23716 7880
rect 23664 7837 23673 7871
rect 23673 7837 23707 7871
rect 23707 7837 23716 7871
rect 23664 7828 23716 7837
rect 23756 7871 23808 7880
rect 23756 7837 23765 7871
rect 23765 7837 23799 7871
rect 23799 7837 23808 7871
rect 23756 7828 23808 7837
rect 23940 7896 23992 7948
rect 24124 7828 24176 7880
rect 24584 7871 24636 7880
rect 24584 7837 24593 7871
rect 24593 7837 24627 7871
rect 24627 7837 24636 7871
rect 24584 7828 24636 7837
rect 24676 7828 24728 7880
rect 26148 7896 26200 7948
rect 27528 7939 27580 7948
rect 27528 7905 27537 7939
rect 27537 7905 27571 7939
rect 27571 7905 27580 7939
rect 27528 7896 27580 7905
rect 24308 7760 24360 7812
rect 24032 7692 24084 7744
rect 25596 7735 25648 7744
rect 25596 7701 25605 7735
rect 25605 7701 25639 7735
rect 25639 7701 25648 7735
rect 25596 7692 25648 7701
rect 25872 7803 25924 7812
rect 25872 7769 25881 7803
rect 25881 7769 25915 7803
rect 25915 7769 25924 7803
rect 25872 7760 25924 7769
rect 26240 7760 26292 7812
rect 26608 7828 26660 7880
rect 26424 7692 26476 7744
rect 8032 7590 8084 7642
rect 8096 7590 8148 7642
rect 8160 7590 8212 7642
rect 8224 7590 8276 7642
rect 8288 7590 8340 7642
rect 15115 7590 15167 7642
rect 15179 7590 15231 7642
rect 15243 7590 15295 7642
rect 15307 7590 15359 7642
rect 15371 7590 15423 7642
rect 22198 7590 22250 7642
rect 22262 7590 22314 7642
rect 22326 7590 22378 7642
rect 22390 7590 22442 7642
rect 22454 7590 22506 7642
rect 29281 7590 29333 7642
rect 29345 7590 29397 7642
rect 29409 7590 29461 7642
rect 29473 7590 29525 7642
rect 29537 7590 29589 7642
rect 5264 7488 5316 7540
rect 5816 7488 5868 7540
rect 6552 7488 6604 7540
rect 12808 7488 12860 7540
rect 5724 7284 5776 7336
rect 10508 7352 10560 7404
rect 11336 7352 11388 7404
rect 12716 7420 12768 7472
rect 12072 7352 12124 7404
rect 14648 7488 14700 7540
rect 16764 7488 16816 7540
rect 16856 7488 16908 7540
rect 14280 7420 14332 7472
rect 13360 7395 13412 7404
rect 13360 7361 13369 7395
rect 13369 7361 13403 7395
rect 13403 7361 13412 7395
rect 13360 7352 13412 7361
rect 13544 7395 13596 7404
rect 13544 7361 13553 7395
rect 13553 7361 13587 7395
rect 13587 7361 13596 7395
rect 13544 7352 13596 7361
rect 4988 7216 5040 7268
rect 6000 7216 6052 7268
rect 11152 7284 11204 7336
rect 11428 7148 11480 7200
rect 11980 7191 12032 7200
rect 11980 7157 11989 7191
rect 11989 7157 12023 7191
rect 12023 7157 12032 7191
rect 11980 7148 12032 7157
rect 14004 7148 14056 7200
rect 15016 7284 15068 7336
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 17960 7488 18012 7540
rect 22652 7488 22704 7540
rect 22928 7531 22980 7540
rect 22928 7497 22937 7531
rect 22937 7497 22971 7531
rect 22971 7497 22980 7531
rect 22928 7488 22980 7497
rect 23020 7488 23072 7540
rect 23388 7488 23440 7540
rect 17408 7395 17460 7404
rect 17408 7361 17417 7395
rect 17417 7361 17451 7395
rect 17451 7361 17460 7395
rect 17408 7352 17460 7361
rect 17500 7395 17552 7404
rect 17500 7361 17509 7395
rect 17509 7361 17543 7395
rect 17543 7361 17552 7395
rect 17500 7352 17552 7361
rect 17684 7352 17736 7404
rect 17868 7395 17920 7404
rect 17868 7361 17877 7395
rect 17877 7361 17911 7395
rect 17911 7361 17920 7395
rect 17868 7352 17920 7361
rect 18052 7395 18104 7404
rect 18052 7361 18061 7395
rect 18061 7361 18095 7395
rect 18095 7361 18104 7395
rect 18052 7352 18104 7361
rect 23480 7420 23532 7472
rect 24584 7420 24636 7472
rect 17040 7216 17092 7268
rect 17776 7216 17828 7268
rect 22100 7352 22152 7404
rect 22284 7284 22336 7336
rect 23112 7284 23164 7336
rect 24032 7395 24084 7404
rect 24032 7361 24041 7395
rect 24041 7361 24075 7395
rect 24075 7361 24084 7395
rect 24032 7352 24084 7361
rect 24308 7352 24360 7404
rect 25596 7488 25648 7540
rect 25872 7488 25924 7540
rect 27528 7488 27580 7540
rect 26516 7420 26568 7472
rect 27068 7420 27120 7472
rect 24952 7395 25004 7404
rect 24952 7361 24961 7395
rect 24961 7361 24995 7395
rect 24995 7361 25004 7395
rect 24952 7352 25004 7361
rect 26240 7352 26292 7404
rect 26608 7352 26660 7404
rect 27344 7352 27396 7404
rect 16764 7191 16816 7200
rect 16764 7157 16773 7191
rect 16773 7157 16807 7191
rect 16807 7157 16816 7191
rect 16764 7148 16816 7157
rect 17408 7148 17460 7200
rect 17868 7191 17920 7200
rect 17868 7157 17877 7191
rect 17877 7157 17911 7191
rect 17911 7157 17920 7191
rect 17868 7148 17920 7157
rect 18328 7148 18380 7200
rect 27804 7352 27856 7404
rect 28724 7395 28776 7404
rect 28724 7361 28733 7395
rect 28733 7361 28767 7395
rect 28767 7361 28776 7395
rect 28724 7352 28776 7361
rect 24124 7148 24176 7200
rect 24400 7191 24452 7200
rect 24400 7157 24409 7191
rect 24409 7157 24443 7191
rect 24443 7157 24452 7191
rect 24400 7148 24452 7157
rect 29000 7191 29052 7200
rect 29000 7157 29009 7191
rect 29009 7157 29043 7191
rect 29043 7157 29052 7191
rect 29000 7148 29052 7157
rect 4491 7046 4543 7098
rect 4555 7046 4607 7098
rect 4619 7046 4671 7098
rect 4683 7046 4735 7098
rect 4747 7046 4799 7098
rect 11574 7046 11626 7098
rect 11638 7046 11690 7098
rect 11702 7046 11754 7098
rect 11766 7046 11818 7098
rect 11830 7046 11882 7098
rect 18657 7046 18709 7098
rect 18721 7046 18773 7098
rect 18785 7046 18837 7098
rect 18849 7046 18901 7098
rect 18913 7046 18965 7098
rect 25740 7046 25792 7098
rect 25804 7046 25856 7098
rect 25868 7046 25920 7098
rect 25932 7046 25984 7098
rect 25996 7046 26048 7098
rect 4988 6944 5040 6996
rect 4620 6740 4672 6792
rect 5908 6808 5960 6860
rect 4988 6740 5040 6792
rect 5080 6740 5132 6792
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 6184 6783 6236 6792
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 6828 6783 6880 6792
rect 6828 6749 6837 6783
rect 6837 6749 6871 6783
rect 6871 6749 6880 6783
rect 6828 6740 6880 6749
rect 7564 6876 7616 6928
rect 7288 6808 7340 6860
rect 10508 6944 10560 6996
rect 10600 6944 10652 6996
rect 11244 6944 11296 6996
rect 11336 6987 11388 6996
rect 11336 6953 11345 6987
rect 11345 6953 11379 6987
rect 11379 6953 11388 6987
rect 11336 6944 11388 6953
rect 11520 6944 11572 6996
rect 12072 6944 12124 6996
rect 13636 6944 13688 6996
rect 7380 6740 7432 6792
rect 7472 6783 7524 6792
rect 7472 6749 7481 6783
rect 7481 6749 7515 6783
rect 7515 6749 7524 6783
rect 7472 6740 7524 6749
rect 7564 6740 7616 6792
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 11428 6808 11480 6860
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 10968 6740 11020 6792
rect 11704 6808 11756 6860
rect 11796 6808 11848 6860
rect 12072 6783 12124 6792
rect 12072 6749 12081 6783
rect 12081 6749 12115 6783
rect 12115 6749 12124 6783
rect 12072 6740 12124 6749
rect 5080 6647 5132 6656
rect 5080 6613 5089 6647
rect 5089 6613 5123 6647
rect 5123 6613 5132 6647
rect 5080 6604 5132 6613
rect 6276 6715 6328 6724
rect 6276 6681 6285 6715
rect 6285 6681 6319 6715
rect 6319 6681 6328 6715
rect 6276 6672 6328 6681
rect 7748 6715 7800 6724
rect 7748 6681 7757 6715
rect 7757 6681 7791 6715
rect 7791 6681 7800 6715
rect 7748 6672 7800 6681
rect 10416 6672 10468 6724
rect 11336 6672 11388 6724
rect 11520 6672 11572 6724
rect 13912 6876 13964 6928
rect 14464 6987 14516 6996
rect 14464 6953 14473 6987
rect 14473 6953 14507 6987
rect 14507 6953 14516 6987
rect 14464 6944 14516 6953
rect 16764 6944 16816 6996
rect 14096 6808 14148 6860
rect 13912 6783 13964 6792
rect 13912 6749 13921 6783
rect 13921 6749 13955 6783
rect 13955 6749 13964 6783
rect 13912 6740 13964 6749
rect 15476 6808 15528 6860
rect 17592 6944 17644 6996
rect 22008 6944 22060 6996
rect 22284 6987 22336 6996
rect 22284 6953 22293 6987
rect 22293 6953 22327 6987
rect 22327 6953 22336 6987
rect 22284 6944 22336 6953
rect 24400 6944 24452 6996
rect 16856 6876 16908 6928
rect 16948 6876 17000 6928
rect 17500 6876 17552 6928
rect 14740 6672 14792 6724
rect 17224 6740 17276 6792
rect 17408 6783 17460 6792
rect 17408 6749 17417 6783
rect 17417 6749 17451 6783
rect 17451 6749 17460 6783
rect 17408 6740 17460 6749
rect 24032 6876 24084 6928
rect 24124 6876 24176 6928
rect 20076 6808 20128 6860
rect 22744 6808 22796 6860
rect 22836 6808 22888 6860
rect 24308 6740 24360 6792
rect 24768 6740 24820 6792
rect 17592 6715 17644 6724
rect 17592 6681 17601 6715
rect 17601 6681 17635 6715
rect 17635 6681 17644 6715
rect 17592 6672 17644 6681
rect 6552 6647 6604 6656
rect 6552 6613 6561 6647
rect 6561 6613 6595 6647
rect 6595 6613 6604 6647
rect 6552 6604 6604 6613
rect 6920 6604 6972 6656
rect 7564 6604 7616 6656
rect 10784 6604 10836 6656
rect 11152 6647 11204 6656
rect 11152 6613 11161 6647
rect 11161 6613 11195 6647
rect 11195 6613 11204 6647
rect 11152 6604 11204 6613
rect 12164 6604 12216 6656
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 17132 6604 17184 6656
rect 20812 6672 20864 6724
rect 17776 6647 17828 6656
rect 17776 6613 17785 6647
rect 17785 6613 17819 6647
rect 17819 6613 17828 6647
rect 17776 6604 17828 6613
rect 17960 6647 18012 6656
rect 17960 6613 17969 6647
rect 17969 6613 18003 6647
rect 18003 6613 18012 6647
rect 17960 6604 18012 6613
rect 18052 6604 18104 6656
rect 26516 6604 26568 6656
rect 8032 6502 8084 6554
rect 8096 6502 8148 6554
rect 8160 6502 8212 6554
rect 8224 6502 8276 6554
rect 8288 6502 8340 6554
rect 15115 6502 15167 6554
rect 15179 6502 15231 6554
rect 15243 6502 15295 6554
rect 15307 6502 15359 6554
rect 15371 6502 15423 6554
rect 22198 6502 22250 6554
rect 22262 6502 22314 6554
rect 22326 6502 22378 6554
rect 22390 6502 22442 6554
rect 22454 6502 22506 6554
rect 29281 6502 29333 6554
rect 29345 6502 29397 6554
rect 29409 6502 29461 6554
rect 29473 6502 29525 6554
rect 29537 6502 29589 6554
rect 5080 6400 5132 6452
rect 5908 6400 5960 6452
rect 6276 6400 6328 6452
rect 7472 6400 7524 6452
rect 10232 6400 10284 6452
rect 11428 6400 11480 6452
rect 11704 6400 11756 6452
rect 11796 6400 11848 6452
rect 6828 6332 6880 6384
rect 10508 6375 10560 6384
rect 10508 6341 10517 6375
rect 10517 6341 10551 6375
rect 10551 6341 10560 6375
rect 10508 6332 10560 6341
rect 2688 6264 2740 6316
rect 3792 6196 3844 6248
rect 6184 6264 6236 6316
rect 5356 6196 5408 6248
rect 5724 6196 5776 6248
rect 7196 6264 7248 6316
rect 7932 6264 7984 6316
rect 9956 6307 10008 6316
rect 9956 6273 9965 6307
rect 9965 6273 9999 6307
rect 9999 6273 10008 6307
rect 9956 6264 10008 6273
rect 10140 6264 10192 6316
rect 10416 6196 10468 6248
rect 7380 6128 7432 6180
rect 7840 6128 7892 6180
rect 10600 6307 10652 6316
rect 10600 6273 10609 6307
rect 10609 6273 10643 6307
rect 10643 6273 10652 6307
rect 10600 6264 10652 6273
rect 10968 6307 11020 6316
rect 10968 6273 10977 6307
rect 10977 6273 11011 6307
rect 11011 6273 11020 6307
rect 10968 6264 11020 6273
rect 11152 6307 11204 6316
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 14096 6400 14148 6452
rect 16580 6400 16632 6452
rect 17776 6400 17828 6452
rect 17960 6400 18012 6452
rect 20076 6443 20128 6452
rect 20076 6409 20085 6443
rect 20085 6409 20119 6443
rect 20119 6409 20128 6443
rect 20076 6400 20128 6409
rect 20536 6400 20588 6452
rect 28724 6400 28776 6452
rect 14188 6332 14240 6384
rect 15476 6375 15528 6384
rect 15476 6341 15485 6375
rect 15485 6341 15519 6375
rect 15519 6341 15528 6375
rect 15476 6332 15528 6341
rect 16856 6332 16908 6384
rect 17868 6332 17920 6384
rect 20260 6307 20312 6316
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 4620 6060 4672 6112
rect 7564 6060 7616 6112
rect 11152 6128 11204 6180
rect 12440 6196 12492 6248
rect 13452 6239 13504 6248
rect 13452 6205 13461 6239
rect 13461 6205 13495 6239
rect 13495 6205 13504 6239
rect 13452 6196 13504 6205
rect 20536 6128 20588 6180
rect 17592 6060 17644 6112
rect 20444 6060 20496 6112
rect 4491 5958 4543 6010
rect 4555 5958 4607 6010
rect 4619 5958 4671 6010
rect 4683 5958 4735 6010
rect 4747 5958 4799 6010
rect 11574 5958 11626 6010
rect 11638 5958 11690 6010
rect 11702 5958 11754 6010
rect 11766 5958 11818 6010
rect 11830 5958 11882 6010
rect 18657 5958 18709 6010
rect 18721 5958 18773 6010
rect 18785 5958 18837 6010
rect 18849 5958 18901 6010
rect 18913 5958 18965 6010
rect 25740 5958 25792 6010
rect 25804 5958 25856 6010
rect 25868 5958 25920 6010
rect 25932 5958 25984 6010
rect 25996 5958 26048 6010
rect 6552 5856 6604 5908
rect 7196 5856 7248 5908
rect 9634 5856 9686 5908
rect 10048 5856 10100 5908
rect 11060 5899 11112 5908
rect 11060 5865 11069 5899
rect 11069 5865 11103 5899
rect 11103 5865 11112 5899
rect 11060 5856 11112 5865
rect 11152 5856 11204 5908
rect 11336 5856 11388 5908
rect 16948 5856 17000 5908
rect 5724 5831 5776 5840
rect 5724 5797 5733 5831
rect 5733 5797 5767 5831
rect 5767 5797 5776 5831
rect 5724 5788 5776 5797
rect 7564 5788 7616 5840
rect 14004 5788 14056 5840
rect 17224 5788 17276 5840
rect 2688 5720 2740 5772
rect 6276 5763 6328 5772
rect 6276 5729 6285 5763
rect 6285 5729 6319 5763
rect 6319 5729 6328 5763
rect 6276 5720 6328 5729
rect 6920 5720 6972 5772
rect 5356 5652 5408 5704
rect 9496 5652 9548 5704
rect 11428 5720 11480 5772
rect 7012 5584 7064 5636
rect 9312 5516 9364 5568
rect 9772 5559 9824 5568
rect 9772 5525 9781 5559
rect 9781 5525 9815 5559
rect 9815 5525 9824 5559
rect 9772 5516 9824 5525
rect 9864 5516 9916 5568
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 11152 5695 11204 5704
rect 11152 5661 11161 5695
rect 11161 5661 11195 5695
rect 11195 5661 11204 5695
rect 11152 5652 11204 5661
rect 11244 5695 11296 5704
rect 11244 5661 11253 5695
rect 11253 5661 11287 5695
rect 11287 5661 11296 5695
rect 11244 5652 11296 5661
rect 17040 5720 17092 5772
rect 17408 5720 17460 5772
rect 10324 5584 10376 5636
rect 10876 5584 10928 5636
rect 11336 5584 11388 5636
rect 11428 5627 11480 5636
rect 11428 5593 11437 5627
rect 11437 5593 11471 5627
rect 11471 5593 11480 5627
rect 11428 5584 11480 5593
rect 17500 5584 17552 5636
rect 11796 5559 11848 5568
rect 11796 5525 11805 5559
rect 11805 5525 11839 5559
rect 11839 5525 11848 5559
rect 11796 5516 11848 5525
rect 16304 5516 16356 5568
rect 17776 5516 17828 5568
rect 18328 5652 18380 5704
rect 17960 5516 18012 5568
rect 18236 5516 18288 5568
rect 18512 5516 18564 5568
rect 8032 5414 8084 5466
rect 8096 5414 8148 5466
rect 8160 5414 8212 5466
rect 8224 5414 8276 5466
rect 8288 5414 8340 5466
rect 15115 5414 15167 5466
rect 15179 5414 15231 5466
rect 15243 5414 15295 5466
rect 15307 5414 15359 5466
rect 15371 5414 15423 5466
rect 22198 5414 22250 5466
rect 22262 5414 22314 5466
rect 22326 5414 22378 5466
rect 22390 5414 22442 5466
rect 22454 5414 22506 5466
rect 29281 5414 29333 5466
rect 29345 5414 29397 5466
rect 29409 5414 29461 5466
rect 29473 5414 29525 5466
rect 29537 5414 29589 5466
rect 7288 5312 7340 5364
rect 7932 5312 7984 5364
rect 7104 5244 7156 5296
rect 6276 5176 6328 5228
rect 8944 5312 8996 5364
rect 9772 5176 9824 5228
rect 9956 5176 10008 5228
rect 10140 5176 10192 5228
rect 10876 5176 10928 5228
rect 12348 5312 12400 5364
rect 12440 5312 12492 5364
rect 14556 5312 14608 5364
rect 17224 5312 17276 5364
rect 17316 5355 17368 5364
rect 17316 5321 17325 5355
rect 17325 5321 17359 5355
rect 17359 5321 17368 5355
rect 17316 5312 17368 5321
rect 11796 5176 11848 5228
rect 10048 5108 10100 5160
rect 11336 5108 11388 5160
rect 12072 5108 12124 5160
rect 12440 5108 12492 5160
rect 10324 4972 10376 5024
rect 14188 5176 14240 5228
rect 16764 5244 16816 5296
rect 17040 5176 17092 5228
rect 16396 5108 16448 5160
rect 17408 5176 17460 5228
rect 17684 5244 17736 5296
rect 17868 5176 17920 5228
rect 18236 5219 18288 5228
rect 18236 5185 18245 5219
rect 18245 5185 18279 5219
rect 18279 5185 18288 5219
rect 18236 5176 18288 5185
rect 18328 5176 18380 5228
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 20260 5312 20312 5364
rect 28264 5355 28316 5364
rect 28264 5321 28273 5355
rect 28273 5321 28307 5355
rect 28307 5321 28316 5355
rect 28264 5312 28316 5321
rect 16856 5015 16908 5024
rect 16856 4981 16865 5015
rect 16865 4981 16899 5015
rect 16899 4981 16908 5015
rect 16856 4972 16908 4981
rect 17040 5015 17092 5024
rect 17040 4981 17049 5015
rect 17049 4981 17083 5015
rect 17083 4981 17092 5015
rect 17040 4972 17092 4981
rect 17132 4972 17184 5024
rect 18052 5040 18104 5092
rect 18144 5040 18196 5092
rect 28080 5219 28132 5228
rect 28080 5185 28089 5219
rect 28089 5185 28123 5219
rect 28123 5185 28132 5219
rect 28080 5176 28132 5185
rect 17868 5015 17920 5024
rect 17868 4981 17877 5015
rect 17877 4981 17911 5015
rect 17911 4981 17920 5015
rect 17868 4972 17920 4981
rect 17960 4972 18012 5024
rect 19524 4972 19576 5024
rect 20720 4972 20772 5024
rect 4491 4870 4543 4922
rect 4555 4870 4607 4922
rect 4619 4870 4671 4922
rect 4683 4870 4735 4922
rect 4747 4870 4799 4922
rect 11574 4870 11626 4922
rect 11638 4870 11690 4922
rect 11702 4870 11754 4922
rect 11766 4870 11818 4922
rect 11830 4870 11882 4922
rect 18657 4870 18709 4922
rect 18721 4870 18773 4922
rect 18785 4870 18837 4922
rect 18849 4870 18901 4922
rect 18913 4870 18965 4922
rect 25740 4870 25792 4922
rect 25804 4870 25856 4922
rect 25868 4870 25920 4922
rect 25932 4870 25984 4922
rect 25996 4870 26048 4922
rect 10140 4768 10192 4820
rect 11060 4768 11112 4820
rect 11428 4768 11480 4820
rect 8944 4675 8996 4684
rect 8944 4641 8953 4675
rect 8953 4641 8987 4675
rect 8987 4641 8996 4675
rect 8944 4632 8996 4641
rect 9312 4675 9364 4684
rect 9312 4641 9321 4675
rect 9321 4641 9355 4675
rect 9355 4641 9364 4675
rect 9312 4632 9364 4641
rect 10324 4632 10376 4684
rect 11336 4564 11388 4616
rect 12992 4564 13044 4616
rect 13268 4607 13320 4616
rect 13268 4573 13277 4607
rect 13277 4573 13311 4607
rect 13311 4573 13320 4607
rect 13268 4564 13320 4573
rect 16304 4768 16356 4820
rect 16488 4768 16540 4820
rect 16948 4811 17000 4820
rect 16948 4777 16957 4811
rect 16957 4777 16991 4811
rect 16991 4777 17000 4811
rect 16948 4768 17000 4777
rect 17592 4811 17644 4820
rect 17592 4777 17601 4811
rect 17601 4777 17635 4811
rect 17635 4777 17644 4811
rect 17592 4768 17644 4777
rect 17868 4768 17920 4820
rect 19800 4768 19852 4820
rect 28080 4768 28132 4820
rect 16028 4675 16080 4684
rect 16028 4641 16037 4675
rect 16037 4641 16071 4675
rect 16071 4641 16080 4675
rect 16028 4632 16080 4641
rect 16396 4564 16448 4616
rect 16488 4607 16540 4616
rect 16488 4573 16497 4607
rect 16497 4573 16531 4607
rect 16531 4573 16540 4607
rect 16488 4564 16540 4573
rect 16580 4607 16632 4616
rect 16580 4573 16589 4607
rect 16589 4573 16623 4607
rect 16623 4573 16632 4607
rect 16580 4564 16632 4573
rect 17040 4632 17092 4684
rect 19340 4700 19392 4752
rect 20536 4700 20588 4752
rect 14004 4496 14056 4548
rect 16212 4539 16264 4548
rect 16212 4505 16221 4539
rect 16221 4505 16255 4539
rect 16255 4505 16264 4539
rect 16212 4496 16264 4505
rect 16304 4496 16356 4548
rect 17408 4607 17460 4616
rect 17408 4573 17417 4607
rect 17417 4573 17451 4607
rect 17451 4573 17460 4607
rect 17408 4564 17460 4573
rect 17868 4564 17920 4616
rect 18052 4564 18104 4616
rect 6460 4428 6512 4480
rect 16856 4428 16908 4480
rect 17592 4496 17644 4548
rect 19524 4675 19576 4684
rect 19524 4641 19533 4675
rect 19533 4641 19567 4675
rect 19567 4641 19576 4675
rect 19524 4632 19576 4641
rect 19248 4564 19300 4616
rect 19432 4607 19484 4616
rect 19432 4573 19441 4607
rect 19441 4573 19475 4607
rect 19475 4573 19484 4607
rect 19432 4564 19484 4573
rect 19800 4564 19852 4616
rect 20168 4607 20220 4616
rect 20168 4573 20177 4607
rect 20177 4573 20211 4607
rect 20211 4573 20220 4607
rect 20168 4564 20220 4573
rect 20444 4564 20496 4616
rect 20720 4607 20772 4616
rect 20720 4573 20729 4607
rect 20729 4573 20763 4607
rect 20763 4573 20772 4607
rect 20720 4564 20772 4573
rect 17224 4471 17276 4480
rect 17224 4437 17233 4471
rect 17233 4437 17267 4471
rect 17267 4437 17276 4471
rect 17224 4428 17276 4437
rect 17684 4428 17736 4480
rect 17868 4428 17920 4480
rect 18236 4428 18288 4480
rect 18328 4428 18380 4480
rect 8032 4326 8084 4378
rect 8096 4326 8148 4378
rect 8160 4326 8212 4378
rect 8224 4326 8276 4378
rect 8288 4326 8340 4378
rect 15115 4326 15167 4378
rect 15179 4326 15231 4378
rect 15243 4326 15295 4378
rect 15307 4326 15359 4378
rect 15371 4326 15423 4378
rect 22198 4326 22250 4378
rect 22262 4326 22314 4378
rect 22326 4326 22378 4378
rect 22390 4326 22442 4378
rect 22454 4326 22506 4378
rect 29281 4326 29333 4378
rect 29345 4326 29397 4378
rect 29409 4326 29461 4378
rect 29473 4326 29525 4378
rect 29537 4326 29589 4378
rect 2412 4224 2464 4276
rect 13176 4267 13228 4276
rect 13176 4233 13185 4267
rect 13185 4233 13219 4267
rect 13219 4233 13228 4267
rect 13176 4224 13228 4233
rect 14188 4224 14240 4276
rect 15568 4224 15620 4276
rect 15844 4224 15896 4276
rect 16028 4224 16080 4276
rect 16856 4224 16908 4276
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 12992 4088 13044 4140
rect 14280 4156 14332 4208
rect 3608 3952 3660 4004
rect 13360 3952 13412 4004
rect 14096 4020 14148 4072
rect 2228 3927 2280 3936
rect 2228 3893 2237 3927
rect 2237 3893 2271 3927
rect 2271 3893 2280 3927
rect 2228 3884 2280 3893
rect 13084 3884 13136 3936
rect 13452 3884 13504 3936
rect 13912 3884 13964 3936
rect 14464 4020 14516 4072
rect 16028 4131 16080 4140
rect 16028 4097 16037 4131
rect 16037 4097 16071 4131
rect 16071 4097 16080 4131
rect 16028 4088 16080 4097
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 16580 4088 16632 4140
rect 16948 4088 17000 4140
rect 17224 4088 17276 4140
rect 17776 4224 17828 4276
rect 19524 4224 19576 4276
rect 20444 4224 20496 4276
rect 20536 4224 20588 4276
rect 19248 4131 19300 4140
rect 19248 4097 19257 4131
rect 19257 4097 19291 4131
rect 19291 4097 19300 4131
rect 19248 4088 19300 4097
rect 19432 4088 19484 4140
rect 19800 4131 19852 4140
rect 19800 4097 19809 4131
rect 19809 4097 19843 4131
rect 19843 4097 19852 4131
rect 19800 4088 19852 4097
rect 24308 4156 24360 4208
rect 24492 4088 24544 4140
rect 17408 4063 17460 4072
rect 17408 4029 17417 4063
rect 17417 4029 17451 4063
rect 17451 4029 17460 4063
rect 17408 4020 17460 4029
rect 19524 4063 19576 4072
rect 19524 4029 19533 4063
rect 19533 4029 19567 4063
rect 19567 4029 19576 4063
rect 19524 4020 19576 4029
rect 19616 4020 19668 4072
rect 15568 3952 15620 4004
rect 22100 3952 22152 4004
rect 14556 3884 14608 3936
rect 16028 3884 16080 3936
rect 17040 3884 17092 3936
rect 17132 3884 17184 3936
rect 18512 3884 18564 3936
rect 20168 3927 20220 3936
rect 20168 3893 20177 3927
rect 20177 3893 20211 3927
rect 20211 3893 20220 3927
rect 20168 3884 20220 3893
rect 24400 3927 24452 3936
rect 24400 3893 24409 3927
rect 24409 3893 24443 3927
rect 24443 3893 24452 3927
rect 24400 3884 24452 3893
rect 24952 3927 25004 3936
rect 24952 3893 24961 3927
rect 24961 3893 24995 3927
rect 24995 3893 25004 3927
rect 24952 3884 25004 3893
rect 4491 3782 4543 3834
rect 4555 3782 4607 3834
rect 4619 3782 4671 3834
rect 4683 3782 4735 3834
rect 4747 3782 4799 3834
rect 11574 3782 11626 3834
rect 11638 3782 11690 3834
rect 11702 3782 11754 3834
rect 11766 3782 11818 3834
rect 11830 3782 11882 3834
rect 18657 3782 18709 3834
rect 18721 3782 18773 3834
rect 18785 3782 18837 3834
rect 18849 3782 18901 3834
rect 18913 3782 18965 3834
rect 25740 3782 25792 3834
rect 25804 3782 25856 3834
rect 25868 3782 25920 3834
rect 25932 3782 25984 3834
rect 25996 3782 26048 3834
rect 2228 3680 2280 3732
rect 13176 3680 13228 3732
rect 14280 3723 14332 3732
rect 14280 3689 14289 3723
rect 14289 3689 14323 3723
rect 14323 3689 14332 3723
rect 14280 3680 14332 3689
rect 12900 3476 12952 3528
rect 13544 3612 13596 3664
rect 14004 3612 14056 3664
rect 15568 3680 15620 3732
rect 15660 3680 15712 3732
rect 19524 3680 19576 3732
rect 14556 3612 14608 3664
rect 15200 3612 15252 3664
rect 24400 3680 24452 3732
rect 24952 3680 25004 3732
rect 13360 3476 13412 3528
rect 13452 3519 13504 3528
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 14096 3544 14148 3596
rect 13820 3476 13872 3528
rect 14188 3476 14240 3528
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 15844 3544 15896 3596
rect 13176 3408 13228 3460
rect 940 3340 992 3392
rect 2228 3383 2280 3392
rect 2228 3349 2237 3383
rect 2237 3349 2271 3383
rect 2271 3349 2280 3383
rect 2228 3340 2280 3349
rect 12808 3383 12860 3392
rect 12808 3349 12817 3383
rect 12817 3349 12851 3383
rect 12851 3349 12860 3383
rect 12808 3340 12860 3349
rect 12900 3340 12952 3392
rect 13728 3340 13780 3392
rect 13912 3408 13964 3460
rect 14280 3340 14332 3392
rect 14372 3340 14424 3392
rect 14648 3340 14700 3392
rect 14924 3340 14976 3392
rect 16580 3476 16632 3528
rect 17040 3519 17092 3528
rect 17040 3485 17049 3519
rect 17049 3485 17083 3519
rect 17083 3485 17092 3519
rect 17040 3476 17092 3485
rect 17592 3544 17644 3596
rect 20168 3544 20220 3596
rect 17776 3408 17828 3460
rect 18512 3476 18564 3528
rect 17500 3383 17552 3392
rect 17500 3349 17509 3383
rect 17509 3349 17543 3383
rect 17543 3349 17552 3383
rect 17500 3340 17552 3349
rect 17592 3340 17644 3392
rect 18788 3383 18840 3392
rect 18788 3349 18797 3383
rect 18797 3349 18831 3383
rect 18831 3349 18840 3383
rect 18788 3340 18840 3349
rect 25228 3383 25280 3392
rect 25228 3349 25237 3383
rect 25237 3349 25271 3383
rect 25271 3349 25280 3383
rect 25228 3340 25280 3349
rect 8032 3238 8084 3290
rect 8096 3238 8148 3290
rect 8160 3238 8212 3290
rect 8224 3238 8276 3290
rect 8288 3238 8340 3290
rect 15115 3238 15167 3290
rect 15179 3238 15231 3290
rect 15243 3238 15295 3290
rect 15307 3238 15359 3290
rect 15371 3238 15423 3290
rect 22198 3238 22250 3290
rect 22262 3238 22314 3290
rect 22326 3238 22378 3290
rect 22390 3238 22442 3290
rect 22454 3238 22506 3290
rect 29281 3238 29333 3290
rect 29345 3238 29397 3290
rect 29409 3238 29461 3290
rect 29473 3238 29525 3290
rect 29537 3238 29589 3290
rect 12992 3179 13044 3188
rect 12992 3145 13001 3179
rect 13001 3145 13035 3179
rect 13035 3145 13044 3179
rect 12992 3136 13044 3145
rect 13084 3136 13136 3188
rect 14556 3179 14608 3188
rect 14556 3145 14565 3179
rect 14565 3145 14599 3179
rect 14599 3145 14608 3179
rect 14556 3136 14608 3145
rect 15660 3136 15712 3188
rect 17500 3136 17552 3188
rect 17592 3179 17644 3188
rect 17592 3145 17601 3179
rect 17601 3145 17635 3179
rect 17635 3145 17644 3179
rect 17592 3136 17644 3145
rect 17776 3136 17828 3188
rect 18788 3136 18840 3188
rect 14096 3068 14148 3120
rect 13544 3000 13596 3052
rect 13360 2864 13412 2916
rect 13912 3000 13964 3052
rect 14004 3043 14056 3052
rect 14004 3009 14013 3043
rect 14013 3009 14047 3043
rect 14047 3009 14056 3043
rect 14004 3000 14056 3009
rect 14924 3068 14976 3120
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 14648 3000 14700 3052
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 17500 2975 17552 2984
rect 17500 2941 17509 2975
rect 17509 2941 17543 2975
rect 17543 2941 17552 2975
rect 17500 2932 17552 2941
rect 18144 3000 18196 3052
rect 18236 3043 18288 3052
rect 18236 3009 18245 3043
rect 18245 3009 18279 3043
rect 18279 3009 18288 3043
rect 18236 3000 18288 3009
rect 17960 2975 18012 2984
rect 17960 2941 17969 2975
rect 17969 2941 18003 2975
rect 18003 2941 18012 2975
rect 17960 2932 18012 2941
rect 13176 2839 13228 2848
rect 13176 2805 13185 2839
rect 13185 2805 13219 2839
rect 13219 2805 13228 2839
rect 13176 2796 13228 2805
rect 13728 2796 13780 2848
rect 14464 2796 14516 2848
rect 17132 2796 17184 2848
rect 19800 2796 19852 2848
rect 29000 2839 29052 2848
rect 29000 2805 29009 2839
rect 29009 2805 29043 2839
rect 29043 2805 29052 2839
rect 29000 2796 29052 2805
rect 4491 2694 4543 2746
rect 4555 2694 4607 2746
rect 4619 2694 4671 2746
rect 4683 2694 4735 2746
rect 4747 2694 4799 2746
rect 11574 2694 11626 2746
rect 11638 2694 11690 2746
rect 11702 2694 11754 2746
rect 11766 2694 11818 2746
rect 11830 2694 11882 2746
rect 18657 2694 18709 2746
rect 18721 2694 18773 2746
rect 18785 2694 18837 2746
rect 18849 2694 18901 2746
rect 18913 2694 18965 2746
rect 25740 2694 25792 2746
rect 25804 2694 25856 2746
rect 25868 2694 25920 2746
rect 25932 2694 25984 2746
rect 25996 2694 26048 2746
rect 2228 2388 2280 2440
rect 12808 2592 12860 2644
rect 13268 2592 13320 2644
rect 13176 2388 13228 2440
rect 13544 2388 13596 2440
rect 13728 2388 13780 2440
rect 27068 2524 27120 2576
rect 19340 2431 19392 2440
rect 19340 2397 19349 2431
rect 19349 2397 19383 2431
rect 19383 2397 19392 2431
rect 19340 2388 19392 2397
rect 22100 2431 22152 2440
rect 22100 2397 22109 2431
rect 22109 2397 22143 2431
rect 22143 2397 22152 2431
rect 22100 2388 22152 2397
rect 25228 2388 25280 2440
rect 28540 2388 28592 2440
rect 17500 2320 17552 2372
rect 29644 2320 29696 2372
rect 20 2252 72 2304
rect 3424 2252 3476 2304
rect 7104 2252 7156 2304
rect 11152 2252 11204 2304
rect 14924 2252 14976 2304
rect 19064 2252 19116 2304
rect 22008 2252 22060 2304
rect 26148 2252 26200 2304
rect 8032 2150 8084 2202
rect 8096 2150 8148 2202
rect 8160 2150 8212 2202
rect 8224 2150 8276 2202
rect 8288 2150 8340 2202
rect 15115 2150 15167 2202
rect 15179 2150 15231 2202
rect 15243 2150 15295 2202
rect 15307 2150 15359 2202
rect 15371 2150 15423 2202
rect 22198 2150 22250 2202
rect 22262 2150 22314 2202
rect 22326 2150 22378 2202
rect 22390 2150 22442 2202
rect 22454 2150 22506 2202
rect 29281 2150 29333 2202
rect 29345 2150 29397 2202
rect 29409 2150 29461 2202
rect 29473 2150 29525 2202
rect 29537 2150 29589 2202
<< metal2 >>
rect 2594 32042 2650 32725
rect 6458 32042 6514 32725
rect 2594 32014 2728 32042
rect 2594 31925 2650 32014
rect 1582 30968 1638 30977
rect 1582 30903 1638 30912
rect 1596 30258 1624 30903
rect 2700 30274 2728 32014
rect 6458 32014 6776 32042
rect 6458 31925 6514 32014
rect 6748 30394 6776 32014
rect 9678 31925 9734 32725
rect 13542 32042 13598 32725
rect 13542 32014 13768 32042
rect 13542 31925 13598 32014
rect 8032 30492 8340 30501
rect 8032 30490 8038 30492
rect 8094 30490 8118 30492
rect 8174 30490 8198 30492
rect 8254 30490 8278 30492
rect 8334 30490 8340 30492
rect 8094 30438 8096 30490
rect 8276 30438 8278 30490
rect 8032 30436 8038 30438
rect 8094 30436 8118 30438
rect 8174 30436 8198 30438
rect 8254 30436 8278 30438
rect 8334 30436 8340 30438
rect 8032 30427 8340 30436
rect 6736 30388 6788 30394
rect 6736 30330 6788 30336
rect 9692 30326 9720 31925
rect 9680 30320 9732 30326
rect 1584 30252 1636 30258
rect 2700 30246 2820 30274
rect 9680 30262 9732 30268
rect 13740 30274 13768 32014
rect 17406 31925 17462 32725
rect 21270 31925 21326 32725
rect 25134 32042 25190 32725
rect 25134 32014 25452 32042
rect 25134 31925 25190 32014
rect 15115 30492 15423 30501
rect 15115 30490 15121 30492
rect 15177 30490 15201 30492
rect 15257 30490 15281 30492
rect 15337 30490 15361 30492
rect 15417 30490 15423 30492
rect 15177 30438 15179 30490
rect 15359 30438 15361 30490
rect 15115 30436 15121 30438
rect 15177 30436 15201 30438
rect 15257 30436 15281 30438
rect 15337 30436 15361 30438
rect 15417 30436 15423 30438
rect 15115 30427 15423 30436
rect 1584 30194 1636 30200
rect 2792 30122 2820 30246
rect 3424 30252 3476 30258
rect 3424 30194 3476 30200
rect 6092 30252 6144 30258
rect 6092 30194 6144 30200
rect 9864 30252 9916 30258
rect 13740 30246 13860 30274
rect 9864 30194 9916 30200
rect 2780 30116 2832 30122
rect 2780 30058 2832 30064
rect 1584 30048 1636 30054
rect 1584 29990 1636 29996
rect 1596 29238 1624 29990
rect 3240 29300 3292 29306
rect 3240 29242 3292 29248
rect 1584 29232 1636 29238
rect 1584 29174 1636 29180
rect 3252 29170 3280 29242
rect 3240 29164 3292 29170
rect 3240 29106 3292 29112
rect 3148 29028 3200 29034
rect 3148 28970 3200 28976
rect 3160 27538 3188 28970
rect 3148 27532 3200 27538
rect 3148 27474 3200 27480
rect 1492 27396 1544 27402
rect 1492 27338 1544 27344
rect 940 27328 992 27334
rect 938 27296 940 27305
rect 992 27296 994 27305
rect 938 27231 994 27240
rect 1504 26586 1532 27338
rect 2780 27328 2832 27334
rect 2780 27270 2832 27276
rect 1492 26580 1544 26586
rect 1492 26522 1544 26528
rect 2412 26376 2464 26382
rect 2412 26318 2464 26324
rect 1492 23724 1544 23730
rect 1492 23666 1544 23672
rect 1504 23089 1532 23666
rect 1584 23520 1636 23526
rect 1582 23488 1584 23497
rect 1636 23488 1638 23497
rect 1582 23423 1638 23432
rect 1490 23080 1546 23089
rect 1490 23015 1546 23024
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1872 19854 1900 20878
rect 1860 19848 1912 19854
rect 1860 19790 1912 19796
rect 1582 19544 1638 19553
rect 1582 19479 1584 19488
rect 1636 19479 1638 19488
rect 1584 19450 1636 19456
rect 1492 19372 1544 19378
rect 1492 19314 1544 19320
rect 1400 16584 1452 16590
rect 1400 16526 1452 16532
rect 940 16108 992 16114
rect 940 16050 992 16056
rect 952 15745 980 16050
rect 1412 16046 1440 16526
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 938 15736 994 15745
rect 938 15671 994 15680
rect 1412 15570 1440 15982
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1412 14958 1440 15506
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1412 13938 1440 14894
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 12850 1440 13874
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 952 11665 980 11698
rect 938 11656 994 11665
rect 938 11591 994 11600
rect 1504 6361 1532 19314
rect 1872 18426 1900 19790
rect 1860 18420 1912 18426
rect 1860 18362 1912 18368
rect 2424 16574 2452 26318
rect 2792 25158 2820 27270
rect 3436 26234 3464 30194
rect 4491 29948 4799 29957
rect 4491 29946 4497 29948
rect 4553 29946 4577 29948
rect 4633 29946 4657 29948
rect 4713 29946 4737 29948
rect 4793 29946 4799 29948
rect 4553 29894 4555 29946
rect 4735 29894 4737 29946
rect 4491 29892 4497 29894
rect 4553 29892 4577 29894
rect 4633 29892 4657 29894
rect 4713 29892 4737 29894
rect 4793 29892 4799 29894
rect 4491 29883 4799 29892
rect 5080 29776 5132 29782
rect 5080 29718 5132 29724
rect 5448 29776 5500 29782
rect 5448 29718 5500 29724
rect 4896 29504 4948 29510
rect 4896 29446 4948 29452
rect 3976 29232 4028 29238
rect 4028 29180 4384 29186
rect 3976 29174 4384 29180
rect 3988 29158 4384 29174
rect 3516 29096 3568 29102
rect 3516 29038 3568 29044
rect 3528 28218 3556 29038
rect 4160 28960 4212 28966
rect 4160 28902 4212 28908
rect 4172 28558 4200 28902
rect 4252 28620 4304 28626
rect 4252 28562 4304 28568
rect 4160 28552 4212 28558
rect 4160 28494 4212 28500
rect 3608 28416 3660 28422
rect 3608 28358 3660 28364
rect 4160 28416 4212 28422
rect 4160 28358 4212 28364
rect 3620 28218 3648 28358
rect 3516 28212 3568 28218
rect 3516 28154 3568 28160
rect 3608 28212 3660 28218
rect 3608 28154 3660 28160
rect 3608 28076 3660 28082
rect 3608 28018 3660 28024
rect 3620 27674 3648 28018
rect 3608 27668 3660 27674
rect 3608 27610 3660 27616
rect 4172 27402 4200 28358
rect 4264 27538 4292 28562
rect 4356 28506 4384 29158
rect 4491 28860 4799 28869
rect 4491 28858 4497 28860
rect 4553 28858 4577 28860
rect 4633 28858 4657 28860
rect 4713 28858 4737 28860
rect 4793 28858 4799 28860
rect 4553 28806 4555 28858
rect 4735 28806 4737 28858
rect 4491 28804 4497 28806
rect 4553 28804 4577 28806
rect 4633 28804 4657 28806
rect 4713 28804 4737 28806
rect 4793 28804 4799 28806
rect 4491 28795 4799 28804
rect 4356 28478 4476 28506
rect 4908 28490 4936 29446
rect 5092 28966 5120 29718
rect 5356 29640 5408 29646
rect 5356 29582 5408 29588
rect 5172 29028 5224 29034
rect 5172 28970 5224 28976
rect 5080 28960 5132 28966
rect 5080 28902 5132 28908
rect 4988 28620 5040 28626
rect 4988 28562 5040 28568
rect 4344 28416 4396 28422
rect 4344 28358 4396 28364
rect 4252 27532 4304 27538
rect 4252 27474 4304 27480
rect 4356 27470 4384 28358
rect 4448 28150 4476 28478
rect 4896 28484 4948 28490
rect 4896 28426 4948 28432
rect 4436 28144 4488 28150
rect 4436 28086 4488 28092
rect 5000 28014 5028 28562
rect 4988 28008 5040 28014
rect 4988 27950 5040 27956
rect 4491 27772 4799 27781
rect 4491 27770 4497 27772
rect 4553 27770 4577 27772
rect 4633 27770 4657 27772
rect 4713 27770 4737 27772
rect 4793 27770 4799 27772
rect 4553 27718 4555 27770
rect 4735 27718 4737 27770
rect 4491 27716 4497 27718
rect 4553 27716 4577 27718
rect 4633 27716 4657 27718
rect 4713 27716 4737 27718
rect 4793 27716 4799 27718
rect 4491 27707 4799 27716
rect 4344 27464 4396 27470
rect 4344 27406 4396 27412
rect 4160 27396 4212 27402
rect 4160 27338 4212 27344
rect 4491 26684 4799 26693
rect 4491 26682 4497 26684
rect 4553 26682 4577 26684
rect 4633 26682 4657 26684
rect 4713 26682 4737 26684
rect 4793 26682 4799 26684
rect 4553 26630 4555 26682
rect 4735 26630 4737 26682
rect 4491 26628 4497 26630
rect 4553 26628 4577 26630
rect 4633 26628 4657 26630
rect 4713 26628 4737 26630
rect 4793 26628 4799 26630
rect 4491 26619 4799 26628
rect 3436 26206 3648 26234
rect 3516 25220 3568 25226
rect 3516 25162 3568 25168
rect 2780 25152 2832 25158
rect 2780 25094 2832 25100
rect 3528 24886 3556 25162
rect 3516 24880 3568 24886
rect 3516 24822 3568 24828
rect 3424 24744 3476 24750
rect 3424 24686 3476 24692
rect 3436 24410 3464 24686
rect 3528 24614 3556 24822
rect 3516 24608 3568 24614
rect 3516 24550 3568 24556
rect 3424 24404 3476 24410
rect 3424 24346 3476 24352
rect 3332 21888 3384 21894
rect 3332 21830 3384 21836
rect 3344 21622 3372 21830
rect 3332 21616 3384 21622
rect 3332 21558 3384 21564
rect 3424 21548 3476 21554
rect 3424 21490 3476 21496
rect 3436 20534 3464 21490
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 3424 20528 3476 20534
rect 3424 20470 3476 20476
rect 3528 20346 3556 20742
rect 3436 20318 3556 20346
rect 3436 19786 3464 20318
rect 3424 19780 3476 19786
rect 3424 19722 3476 19728
rect 3436 19334 3464 19722
rect 3252 19306 3464 19334
rect 3252 18290 3280 19306
rect 3516 18760 3568 18766
rect 3516 18702 3568 18708
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 3252 17882 3280 18226
rect 3528 18222 3556 18702
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3240 17876 3292 17882
rect 3240 17818 3292 17824
rect 3436 17610 3464 18158
rect 3424 17604 3476 17610
rect 3424 17546 3476 17552
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 2332 16546 2452 16574
rect 1676 16516 1728 16522
rect 1676 16458 1728 16464
rect 1688 16250 1716 16458
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 1872 13530 1900 13806
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 2056 12442 2084 12718
rect 2044 12436 2096 12442
rect 2044 12378 2096 12384
rect 2226 11792 2282 11801
rect 2226 11727 2228 11736
rect 2280 11727 2282 11736
rect 2228 11698 2280 11704
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2240 11218 2268 11494
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2240 9654 2268 11154
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2240 9042 2268 9590
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2240 8634 2268 8978
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1688 7886 1716 8434
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 2332 6914 2360 16546
rect 3344 15570 3372 16934
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3252 14006 3280 15438
rect 3528 14006 3556 17070
rect 3240 14000 3292 14006
rect 3160 13960 3240 13988
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 3068 12345 3096 13262
rect 3160 12850 3188 13960
rect 3240 13942 3292 13948
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 3528 13394 3556 13942
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3054 12336 3110 12345
rect 3054 12271 3110 12280
rect 3068 12238 3096 12271
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 3160 11830 3188 12786
rect 3252 12238 3280 13126
rect 3528 12918 3556 13330
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 3528 12306 3556 12854
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3148 11824 3200 11830
rect 3148 11766 3200 11772
rect 3160 11150 3188 11766
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3160 9674 3188 11086
rect 3160 9646 3372 9674
rect 3344 9586 3372 9646
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 2332 6886 2452 6914
rect 1490 6352 1546 6361
rect 1490 6287 1546 6296
rect 2424 4282 2452 6886
rect 2700 6322 2728 8502
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2700 5778 2728 6258
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2424 4049 2452 4082
rect 2410 4040 2466 4049
rect 3620 4010 3648 26206
rect 4344 25696 4396 25702
rect 4344 25638 4396 25644
rect 4356 25294 4384 25638
rect 4491 25596 4799 25605
rect 4491 25594 4497 25596
rect 4553 25594 4577 25596
rect 4633 25594 4657 25596
rect 4713 25594 4737 25596
rect 4793 25594 4799 25596
rect 4553 25542 4555 25594
rect 4735 25542 4737 25594
rect 4491 25540 4497 25542
rect 4553 25540 4577 25542
rect 4633 25540 4657 25542
rect 4713 25540 4737 25542
rect 4793 25540 4799 25542
rect 4491 25531 4799 25540
rect 5000 25362 5028 27950
rect 5092 27878 5120 28902
rect 5184 28762 5212 28970
rect 5264 28960 5316 28966
rect 5264 28902 5316 28908
rect 5172 28756 5224 28762
rect 5172 28698 5224 28704
rect 5276 28490 5304 28902
rect 5264 28484 5316 28490
rect 5264 28426 5316 28432
rect 5276 28218 5304 28426
rect 5368 28422 5396 29582
rect 5460 29102 5488 29718
rect 5724 29640 5776 29646
rect 5724 29582 5776 29588
rect 5448 29096 5500 29102
rect 5448 29038 5500 29044
rect 5356 28416 5408 28422
rect 5356 28358 5408 28364
rect 5460 28218 5488 29038
rect 5736 28762 5764 29582
rect 6000 29572 6052 29578
rect 6000 29514 6052 29520
rect 5816 29504 5868 29510
rect 5816 29446 5868 29452
rect 5724 28756 5776 28762
rect 5724 28698 5776 28704
rect 5264 28212 5316 28218
rect 5448 28212 5500 28218
rect 5316 28172 5396 28200
rect 5264 28154 5316 28160
rect 5368 28098 5396 28172
rect 5448 28154 5500 28160
rect 5368 28070 5764 28098
rect 5080 27872 5132 27878
rect 5080 27814 5132 27820
rect 5448 27872 5500 27878
rect 5448 27814 5500 27820
rect 5460 27470 5488 27814
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 5172 27396 5224 27402
rect 5172 27338 5224 27344
rect 5184 25906 5212 27338
rect 5172 25900 5224 25906
rect 5172 25842 5224 25848
rect 5356 25900 5408 25906
rect 5356 25842 5408 25848
rect 5080 25696 5132 25702
rect 5080 25638 5132 25644
rect 5092 25498 5120 25638
rect 5080 25492 5132 25498
rect 5080 25434 5132 25440
rect 4988 25356 5040 25362
rect 4988 25298 5040 25304
rect 4344 25288 4396 25294
rect 4344 25230 4396 25236
rect 4620 25288 4672 25294
rect 4620 25230 4672 25236
rect 4632 24750 4660 25230
rect 4896 25152 4948 25158
rect 4896 25094 4948 25100
rect 4908 24886 4936 25094
rect 5000 24886 5028 25298
rect 5080 25152 5132 25158
rect 5080 25094 5132 25100
rect 4896 24880 4948 24886
rect 4896 24822 4948 24828
rect 4988 24880 5040 24886
rect 4988 24822 5040 24828
rect 4620 24744 4672 24750
rect 4620 24686 4672 24692
rect 4491 24508 4799 24517
rect 4491 24506 4497 24508
rect 4553 24506 4577 24508
rect 4633 24506 4657 24508
rect 4713 24506 4737 24508
rect 4793 24506 4799 24508
rect 4553 24454 4555 24506
rect 4735 24454 4737 24506
rect 4491 24452 4497 24454
rect 4553 24452 4577 24454
rect 4633 24452 4657 24454
rect 4713 24452 4737 24454
rect 4793 24452 4799 24454
rect 4491 24443 4799 24452
rect 5000 24274 5028 24822
rect 5092 24614 5120 25094
rect 5080 24608 5132 24614
rect 5080 24550 5132 24556
rect 4988 24268 5040 24274
rect 4988 24210 5040 24216
rect 4491 23420 4799 23429
rect 4491 23418 4497 23420
rect 4553 23418 4577 23420
rect 4633 23418 4657 23420
rect 4713 23418 4737 23420
rect 4793 23418 4799 23420
rect 4553 23366 4555 23418
rect 4735 23366 4737 23418
rect 4491 23364 4497 23366
rect 4553 23364 4577 23366
rect 4633 23364 4657 23366
rect 4713 23364 4737 23366
rect 4793 23364 4799 23366
rect 4491 23355 4799 23364
rect 5092 23066 5120 24550
rect 5184 23866 5212 25842
rect 5368 25362 5396 25842
rect 5540 25832 5592 25838
rect 5540 25774 5592 25780
rect 5736 25786 5764 28070
rect 5828 27946 5856 29446
rect 6012 28218 6040 29514
rect 6000 28212 6052 28218
rect 6000 28154 6052 28160
rect 5816 27940 5868 27946
rect 5816 27882 5868 27888
rect 5816 26240 5868 26246
rect 5816 26182 5868 26188
rect 5828 25974 5856 26182
rect 5816 25968 5868 25974
rect 5816 25910 5868 25916
rect 5552 25498 5580 25774
rect 5736 25758 5856 25786
rect 5632 25696 5684 25702
rect 5632 25638 5684 25644
rect 5724 25696 5776 25702
rect 5724 25638 5776 25644
rect 5540 25492 5592 25498
rect 5540 25434 5592 25440
rect 5356 25356 5408 25362
rect 5356 25298 5408 25304
rect 5264 25220 5316 25226
rect 5264 25162 5316 25168
rect 5276 24954 5304 25162
rect 5264 24948 5316 24954
rect 5264 24890 5316 24896
rect 5368 24834 5396 25298
rect 5448 24948 5500 24954
rect 5448 24890 5500 24896
rect 5276 24806 5396 24834
rect 5276 24682 5304 24806
rect 5264 24676 5316 24682
rect 5264 24618 5316 24624
rect 5356 24404 5408 24410
rect 5460 24392 5488 24890
rect 5644 24818 5672 25638
rect 5736 25158 5764 25638
rect 5724 25152 5776 25158
rect 5724 25094 5776 25100
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 5736 24750 5764 25094
rect 5724 24744 5776 24750
rect 5724 24686 5776 24692
rect 5828 24664 5856 25758
rect 6000 24676 6052 24682
rect 5828 24636 6000 24664
rect 6000 24618 6052 24624
rect 5408 24364 5488 24392
rect 5356 24346 5408 24352
rect 6012 24138 6040 24618
rect 6000 24132 6052 24138
rect 6000 24074 6052 24080
rect 5172 23860 5224 23866
rect 5172 23802 5224 23808
rect 5724 23792 5776 23798
rect 5724 23734 5776 23740
rect 5092 23038 5212 23066
rect 5080 22976 5132 22982
rect 5080 22918 5132 22924
rect 4160 22432 4212 22438
rect 4160 22374 4212 22380
rect 4068 21888 4120 21894
rect 4068 21830 4120 21836
rect 4080 21570 4108 21830
rect 4172 21690 4200 22374
rect 4491 22332 4799 22341
rect 4491 22330 4497 22332
rect 4553 22330 4577 22332
rect 4633 22330 4657 22332
rect 4713 22330 4737 22332
rect 4793 22330 4799 22332
rect 4553 22278 4555 22330
rect 4735 22278 4737 22330
rect 4491 22276 4497 22278
rect 4553 22276 4577 22278
rect 4633 22276 4657 22278
rect 4713 22276 4737 22278
rect 4793 22276 4799 22278
rect 4491 22267 4799 22276
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 4160 21684 4212 21690
rect 4160 21626 4212 21632
rect 4158 21584 4214 21593
rect 4080 21542 4158 21570
rect 4158 21519 4214 21528
rect 3700 21344 3752 21350
rect 3700 21286 3752 21292
rect 3792 21344 3844 21350
rect 3792 21286 3844 21292
rect 4068 21344 4120 21350
rect 4068 21286 4120 21292
rect 3712 21146 3740 21286
rect 3700 21140 3752 21146
rect 3700 21082 3752 21088
rect 3804 21010 3832 21286
rect 3792 21004 3844 21010
rect 3792 20946 3844 20952
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3896 20058 3924 20198
rect 3988 20058 4016 20538
rect 4080 20534 4108 21286
rect 4068 20528 4120 20534
rect 4068 20470 4120 20476
rect 3884 20052 3936 20058
rect 3884 19994 3936 20000
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 3976 18624 4028 18630
rect 3976 18566 4028 18572
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 3712 18290 3740 18362
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 3712 17746 3740 18226
rect 3700 17740 3752 17746
rect 3700 17682 3752 17688
rect 3700 17332 3752 17338
rect 3752 17292 3924 17320
rect 3700 17274 3752 17280
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3804 12209 3832 17138
rect 3896 17082 3924 17292
rect 3988 17202 4016 18566
rect 4172 17626 4200 21519
rect 4264 20534 4292 21966
rect 4436 21956 4488 21962
rect 4436 21898 4488 21904
rect 4448 21690 4476 21898
rect 4528 21888 4580 21894
rect 4528 21830 4580 21836
rect 4436 21684 4488 21690
rect 4436 21626 4488 21632
rect 4540 21622 4568 21830
rect 4528 21616 4580 21622
rect 4356 21564 4528 21570
rect 4356 21558 4580 21564
rect 4356 21542 4568 21558
rect 4356 20806 4384 21542
rect 5092 21486 5120 22918
rect 5184 21894 5212 23038
rect 5264 22976 5316 22982
rect 5264 22918 5316 22924
rect 5276 22710 5304 22918
rect 5264 22704 5316 22710
rect 5264 22646 5316 22652
rect 5632 22568 5684 22574
rect 5632 22510 5684 22516
rect 5356 22024 5408 22030
rect 5448 22024 5500 22030
rect 5356 21966 5408 21972
rect 5446 21992 5448 22001
rect 5500 21992 5502 22001
rect 5172 21888 5224 21894
rect 5172 21830 5224 21836
rect 5368 21690 5396 21966
rect 5446 21927 5502 21936
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 5080 21480 5132 21486
rect 5080 21422 5132 21428
rect 4491 21244 4799 21253
rect 4491 21242 4497 21244
rect 4553 21242 4577 21244
rect 4633 21242 4657 21244
rect 4713 21242 4737 21244
rect 4793 21242 4799 21244
rect 4553 21190 4555 21242
rect 4735 21190 4737 21242
rect 4491 21188 4497 21190
rect 4553 21188 4577 21190
rect 4633 21188 4657 21190
rect 4713 21188 4737 21190
rect 4793 21188 4799 21190
rect 4491 21179 4799 21188
rect 5368 20942 5396 21626
rect 5644 21146 5672 22510
rect 5736 21486 5764 23734
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 6012 22098 6040 22510
rect 6000 22092 6052 22098
rect 6000 22034 6052 22040
rect 5908 22024 5960 22030
rect 5908 21966 5960 21972
rect 5920 21690 5948 21966
rect 5908 21684 5960 21690
rect 5908 21626 5960 21632
rect 5816 21548 5868 21554
rect 6000 21548 6052 21554
rect 5816 21490 5868 21496
rect 5920 21508 6000 21536
rect 5724 21480 5776 21486
rect 5828 21457 5856 21490
rect 5724 21422 5776 21428
rect 5814 21448 5870 21457
rect 5814 21383 5870 21392
rect 5920 21321 5948 21508
rect 6000 21490 6052 21496
rect 5906 21312 5962 21321
rect 5906 21247 5962 21256
rect 5632 21140 5684 21146
rect 5632 21082 5684 21088
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 5644 20806 5672 21082
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 4344 20800 4396 20806
rect 4344 20742 4396 20748
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 5356 20460 5408 20466
rect 5356 20402 5408 20408
rect 4896 20392 4948 20398
rect 4894 20360 4896 20369
rect 4948 20360 4950 20369
rect 4894 20295 4950 20304
rect 4491 20156 4799 20165
rect 4491 20154 4497 20156
rect 4553 20154 4577 20156
rect 4633 20154 4657 20156
rect 4713 20154 4737 20156
rect 4793 20154 4799 20156
rect 4553 20102 4555 20154
rect 4735 20102 4737 20154
rect 4491 20100 4497 20102
rect 4553 20100 4577 20102
rect 4633 20100 4657 20102
rect 4713 20100 4737 20102
rect 4793 20100 4799 20102
rect 4491 20091 4799 20100
rect 4491 19068 4799 19077
rect 4491 19066 4497 19068
rect 4553 19066 4577 19068
rect 4633 19066 4657 19068
rect 4713 19066 4737 19068
rect 4793 19066 4799 19068
rect 4553 19014 4555 19066
rect 4735 19014 4737 19066
rect 4491 19012 4497 19014
rect 4553 19012 4577 19014
rect 4633 19012 4657 19014
rect 4713 19012 4737 19014
rect 4793 19012 4799 19014
rect 4491 19003 4799 19012
rect 4491 17980 4799 17989
rect 4491 17978 4497 17980
rect 4553 17978 4577 17980
rect 4633 17978 4657 17980
rect 4713 17978 4737 17980
rect 4793 17978 4799 17980
rect 4553 17926 4555 17978
rect 4735 17926 4737 17978
rect 4491 17924 4497 17926
rect 4553 17924 4577 17926
rect 4633 17924 4657 17926
rect 4713 17924 4737 17926
rect 4793 17924 4799 17926
rect 4491 17915 4799 17924
rect 4080 17598 4200 17626
rect 4528 17604 4580 17610
rect 4080 17202 4108 17598
rect 4528 17546 4580 17552
rect 4804 17604 4856 17610
rect 4804 17546 4856 17552
rect 4540 17338 4568 17546
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4528 17332 4580 17338
rect 4528 17274 4580 17280
rect 4356 17202 4384 17274
rect 4816 17270 4844 17546
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 4908 17218 4936 20295
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5276 18358 5304 18566
rect 5264 18352 5316 18358
rect 5264 18294 5316 18300
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 5080 18148 5132 18154
rect 5080 18090 5132 18096
rect 5092 17338 5120 18090
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5184 17678 5212 18022
rect 5276 17882 5304 18158
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5172 17536 5224 17542
rect 5172 17478 5224 17484
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4528 17196 4580 17202
rect 4908 17190 5120 17218
rect 4528 17138 4580 17144
rect 4080 17082 4108 17138
rect 3896 17054 4108 17082
rect 3884 16516 3936 16522
rect 3884 16458 3936 16464
rect 3896 16114 3924 16458
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 3896 15502 3924 16050
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 3988 13818 4016 17054
rect 4264 16658 4292 17138
rect 4540 17082 4568 17138
rect 4804 17128 4856 17134
rect 4618 17096 4674 17105
rect 4540 17054 4618 17082
rect 4856 17088 4936 17116
rect 4804 17070 4856 17076
rect 4618 17031 4674 17040
rect 4491 16892 4799 16901
rect 4491 16890 4497 16892
rect 4553 16890 4577 16892
rect 4633 16890 4657 16892
rect 4713 16890 4737 16892
rect 4793 16890 4799 16892
rect 4553 16838 4555 16890
rect 4735 16838 4737 16890
rect 4491 16836 4497 16838
rect 4553 16836 4577 16838
rect 4633 16836 4657 16838
rect 4713 16836 4737 16838
rect 4793 16836 4799 16838
rect 4491 16827 4799 16836
rect 4908 16658 4936 17088
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 4448 16250 4476 16390
rect 5000 16250 5028 16934
rect 5092 16726 5120 17190
rect 5184 17066 5212 17478
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5276 17105 5304 17138
rect 5262 17096 5318 17105
rect 5172 17060 5224 17066
rect 5262 17031 5264 17040
rect 5172 17002 5224 17008
rect 5316 17031 5318 17040
rect 5264 17002 5316 17008
rect 5080 16720 5132 16726
rect 5080 16662 5132 16668
rect 5092 16590 5120 16662
rect 5368 16590 5396 20402
rect 5828 18714 5856 20878
rect 5920 19334 5948 21247
rect 5920 19306 6040 19334
rect 5736 18686 5856 18714
rect 5736 18290 5764 18686
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5828 17610 5856 18566
rect 5816 17604 5868 17610
rect 5816 17546 5868 17552
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5460 17270 5488 17478
rect 5448 17264 5500 17270
rect 5448 17206 5500 17212
rect 6012 17202 6040 19306
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 5552 16794 5580 17138
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5080 16584 5132 16590
rect 5356 16584 5408 16590
rect 5080 16526 5132 16532
rect 5276 16544 5356 16572
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 4344 15972 4396 15978
rect 4344 15914 4396 15920
rect 4356 15706 4384 15914
rect 4491 15804 4799 15813
rect 4491 15802 4497 15804
rect 4553 15802 4577 15804
rect 4633 15802 4657 15804
rect 4713 15802 4737 15804
rect 4793 15802 4799 15804
rect 4553 15750 4555 15802
rect 4735 15750 4737 15802
rect 4491 15748 4497 15750
rect 4553 15748 4577 15750
rect 4633 15748 4657 15750
rect 4713 15748 4737 15750
rect 4793 15748 4799 15750
rect 4491 15739 4799 15748
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4068 15496 4120 15502
rect 4066 15464 4068 15473
rect 4120 15464 4122 15473
rect 4066 15399 4122 15408
rect 4080 14958 4108 15399
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4491 14716 4799 14725
rect 4491 14714 4497 14716
rect 4553 14714 4577 14716
rect 4633 14714 4657 14716
rect 4713 14714 4737 14716
rect 4793 14714 4799 14716
rect 4553 14662 4555 14714
rect 4735 14662 4737 14714
rect 4491 14660 4497 14662
rect 4553 14660 4577 14662
rect 4633 14660 4657 14662
rect 4713 14660 4737 14662
rect 4793 14660 4799 14662
rect 4491 14651 4799 14660
rect 3988 13790 4108 13818
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3790 12200 3846 12209
rect 3790 12135 3846 12144
rect 3896 12102 3924 12582
rect 4080 12434 4108 13790
rect 4491 13628 4799 13637
rect 4491 13626 4497 13628
rect 4553 13626 4577 13628
rect 4633 13626 4657 13628
rect 4713 13626 4737 13628
rect 4793 13626 4799 13628
rect 4553 13574 4555 13626
rect 4735 13574 4737 13626
rect 4491 13572 4497 13574
rect 4553 13572 4577 13574
rect 4633 13572 4657 13574
rect 4713 13572 4737 13574
rect 4793 13572 4799 13574
rect 4491 13563 4799 13572
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 3988 12406 4108 12434
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3896 11082 3924 12038
rect 3988 11150 4016 12406
rect 4264 12374 4292 12582
rect 4491 12540 4799 12549
rect 4491 12538 4497 12540
rect 4553 12538 4577 12540
rect 4633 12538 4657 12540
rect 4713 12538 4737 12540
rect 4793 12538 4799 12540
rect 4553 12486 4555 12538
rect 4735 12486 4737 12538
rect 4491 12484 4497 12486
rect 4553 12484 4577 12486
rect 4633 12484 4657 12486
rect 4713 12484 4737 12486
rect 4793 12484 4799 12486
rect 4491 12475 4799 12484
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4448 11898 4476 12174
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4252 11552 4304 11558
rect 4080 11512 4252 11540
rect 4080 11218 4108 11512
rect 4252 11494 4304 11500
rect 4356 11354 4384 11630
rect 4632 11608 4660 12174
rect 4908 11830 4936 12786
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 5000 11898 5028 12242
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 4896 11824 4948 11830
rect 4896 11766 4948 11772
rect 4712 11620 4764 11626
rect 4632 11580 4712 11608
rect 4712 11562 4764 11568
rect 4491 11452 4799 11461
rect 4491 11450 4497 11452
rect 4553 11450 4577 11452
rect 4633 11450 4657 11452
rect 4713 11450 4737 11452
rect 4793 11450 4799 11452
rect 4553 11398 4555 11450
rect 4735 11398 4737 11450
rect 4491 11396 4497 11398
rect 4553 11396 4577 11398
rect 4633 11396 4657 11398
rect 4713 11396 4737 11398
rect 4793 11396 4799 11398
rect 4491 11387 4799 11396
rect 4908 11354 4936 11766
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 3976 11144 4028 11150
rect 4028 11092 4108 11098
rect 3976 11086 4108 11092
rect 3884 11076 3936 11082
rect 3988 11070 4108 11086
rect 3884 11018 3936 11024
rect 4080 10690 4108 11070
rect 4172 10810 4200 11290
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4804 11280 4856 11286
rect 4856 11228 4936 11234
rect 4804 11222 4936 11228
rect 4264 11082 4292 11222
rect 4816 11206 4936 11222
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4080 10662 4292 10690
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 3988 10198 4016 10542
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4080 10266 4108 10406
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4080 9654 4108 9998
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3804 8906 3832 9522
rect 4080 9489 4108 9590
rect 4172 9518 4200 10406
rect 4160 9512 4212 9518
rect 4066 9480 4122 9489
rect 4160 9454 4212 9460
rect 4066 9415 4122 9424
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 3804 8498 3832 8842
rect 4172 8634 4200 9046
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4264 8514 4292 10662
rect 4632 10538 4660 10950
rect 4724 10674 4752 10950
rect 4816 10742 4844 11086
rect 4804 10736 4856 10742
rect 4804 10678 4856 10684
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4491 10364 4799 10373
rect 4491 10362 4497 10364
rect 4553 10362 4577 10364
rect 4633 10362 4657 10364
rect 4713 10362 4737 10364
rect 4793 10362 4799 10364
rect 4553 10310 4555 10362
rect 4735 10310 4737 10362
rect 4491 10308 4497 10310
rect 4553 10308 4577 10310
rect 4633 10308 4657 10310
rect 4713 10308 4737 10310
rect 4793 10308 4799 10310
rect 4491 10299 4799 10308
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4356 9042 4384 9318
rect 4491 9276 4799 9285
rect 4491 9274 4497 9276
rect 4553 9274 4577 9276
rect 4633 9274 4657 9276
rect 4713 9274 4737 9276
rect 4793 9274 4799 9276
rect 4553 9222 4555 9274
rect 4735 9222 4737 9274
rect 4491 9220 4497 9222
rect 4553 9220 4577 9222
rect 4633 9220 4657 9222
rect 4713 9220 4737 9222
rect 4793 9220 4799 9222
rect 4491 9211 4799 9220
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4172 8498 4292 8514
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 4160 8492 4292 8498
rect 4212 8486 4292 8492
rect 4160 8434 4212 8440
rect 3804 7818 3832 8434
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 3792 7812 3844 7818
rect 3792 7754 3844 7760
rect 3804 6254 3832 7754
rect 4080 7585 4108 7958
rect 4264 7818 4292 8486
rect 4356 8362 4384 8774
rect 4908 8650 4936 11206
rect 5000 10538 5028 11834
rect 5092 11218 5120 16526
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5184 12306 5212 12922
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5170 12200 5226 12209
rect 5170 12135 5226 12144
rect 5184 11286 5212 12135
rect 5172 11280 5224 11286
rect 5172 11222 5224 11228
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 5000 9450 5028 10474
rect 5092 9674 5120 11154
rect 5276 10606 5304 16544
rect 5356 16526 5408 16532
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5460 16250 5488 16390
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5460 15026 5488 16050
rect 5448 15020 5500 15026
rect 5448 14962 5500 14968
rect 5552 14958 5580 16390
rect 5736 16114 5764 16526
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5644 15178 5672 16050
rect 5736 15706 5764 16050
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5828 15502 5856 16934
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5644 15162 5764 15178
rect 5644 15156 5776 15162
rect 5644 15150 5724 15156
rect 5724 15098 5776 15104
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5736 13938 5764 15098
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5920 13734 5948 17138
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 6012 13462 6040 17138
rect 6000 13456 6052 13462
rect 6000 13398 6052 13404
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 5356 12164 5408 12170
rect 5356 12106 5408 12112
rect 5368 10742 5396 12106
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5460 11218 5488 11630
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5552 10742 5580 12038
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5920 10810 5948 10950
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 5356 10736 5408 10742
rect 5356 10678 5408 10684
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5264 10600 5316 10606
rect 5316 10560 5488 10588
rect 5264 10542 5316 10548
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 5092 9646 5212 9674
rect 5184 9586 5212 9646
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 5000 9110 5028 9386
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 4816 8622 5028 8650
rect 4816 8498 4844 8622
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4491 8188 4799 8197
rect 4491 8186 4497 8188
rect 4553 8186 4577 8188
rect 4633 8186 4657 8188
rect 4713 8186 4737 8188
rect 4793 8186 4799 8188
rect 4553 8134 4555 8186
rect 4735 8134 4737 8186
rect 4491 8132 4497 8134
rect 4553 8132 4577 8134
rect 4633 8132 4657 8134
rect 4713 8132 4737 8134
rect 4793 8132 4799 8134
rect 4491 8123 4799 8132
rect 5000 7886 5028 8622
rect 5092 8430 5120 9318
rect 5080 8424 5132 8430
rect 5276 8378 5304 10134
rect 5460 9625 5488 10560
rect 6012 9674 6040 12650
rect 6104 9738 6132 30194
rect 9036 29640 9088 29646
rect 9036 29582 9088 29588
rect 7380 29572 7432 29578
rect 7380 29514 7432 29520
rect 7564 29572 7616 29578
rect 7564 29514 7616 29520
rect 7024 29430 7328 29458
rect 7024 29186 7052 29430
rect 7104 29300 7156 29306
rect 7104 29242 7156 29248
rect 6840 29170 7052 29186
rect 6828 29164 7052 29170
rect 6880 29158 7052 29164
rect 6828 29106 6880 29112
rect 7116 28994 7144 29242
rect 6932 28966 7144 28994
rect 6920 28960 6972 28966
rect 6920 28902 6972 28908
rect 7196 28960 7248 28966
rect 7196 28902 7248 28908
rect 7208 28642 7236 28902
rect 6368 28620 6420 28626
rect 6368 28562 6420 28568
rect 7116 28614 7236 28642
rect 6184 28484 6236 28490
rect 6184 28426 6236 28432
rect 6196 28150 6224 28426
rect 6184 28144 6236 28150
rect 6184 28086 6236 28092
rect 6380 27878 6408 28562
rect 6460 28552 6512 28558
rect 6460 28494 6512 28500
rect 6472 28014 6500 28494
rect 7116 28422 7144 28614
rect 7300 28558 7328 29430
rect 7392 28966 7420 29514
rect 7472 29232 7524 29238
rect 7472 29174 7524 29180
rect 7380 28960 7432 28966
rect 7380 28902 7432 28908
rect 7288 28552 7340 28558
rect 7288 28494 7340 28500
rect 7196 28484 7248 28490
rect 7196 28426 7248 28432
rect 7012 28416 7064 28422
rect 7012 28358 7064 28364
rect 7104 28416 7156 28422
rect 7104 28358 7156 28364
rect 7024 28218 7052 28358
rect 7012 28212 7064 28218
rect 7012 28154 7064 28160
rect 7116 28082 7144 28358
rect 7104 28076 7156 28082
rect 7104 28018 7156 28024
rect 6460 28008 6512 28014
rect 6460 27950 6512 27956
rect 7116 27946 7144 28018
rect 7104 27940 7156 27946
rect 7104 27882 7156 27888
rect 6368 27872 6420 27878
rect 6368 27814 6420 27820
rect 6552 27872 6604 27878
rect 6552 27814 6604 27820
rect 6276 26376 6328 26382
rect 6276 26318 6328 26324
rect 6288 26234 6316 26318
rect 6288 26206 6500 26234
rect 6472 25974 6500 26206
rect 6460 25968 6512 25974
rect 6460 25910 6512 25916
rect 6472 25498 6500 25910
rect 6564 25906 6592 27814
rect 7208 27606 7236 28426
rect 7288 28416 7340 28422
rect 7288 28358 7340 28364
rect 7300 28218 7328 28358
rect 7288 28212 7340 28218
rect 7288 28154 7340 28160
rect 7484 28014 7512 29174
rect 7576 29102 7604 29514
rect 7748 29504 7800 29510
rect 7748 29446 7800 29452
rect 7564 29096 7616 29102
rect 7564 29038 7616 29044
rect 7576 28558 7604 29038
rect 7760 28762 7788 29446
rect 8032 29404 8340 29413
rect 8032 29402 8038 29404
rect 8094 29402 8118 29404
rect 8174 29402 8198 29404
rect 8254 29402 8278 29404
rect 8334 29402 8340 29404
rect 8094 29350 8096 29402
rect 8276 29350 8278 29402
rect 8032 29348 8038 29350
rect 8094 29348 8118 29350
rect 8174 29348 8198 29350
rect 8254 29348 8278 29350
rect 8334 29348 8340 29350
rect 8032 29339 8340 29348
rect 8484 29232 8536 29238
rect 8484 29174 8536 29180
rect 7840 28960 7892 28966
rect 7840 28902 7892 28908
rect 7748 28756 7800 28762
rect 7748 28698 7800 28704
rect 7564 28552 7616 28558
rect 7564 28494 7616 28500
rect 7576 28082 7604 28494
rect 7852 28490 7880 28902
rect 7840 28484 7892 28490
rect 7840 28426 7892 28432
rect 8032 28316 8340 28325
rect 8032 28314 8038 28316
rect 8094 28314 8118 28316
rect 8174 28314 8198 28316
rect 8254 28314 8278 28316
rect 8334 28314 8340 28316
rect 8094 28262 8096 28314
rect 8276 28262 8278 28314
rect 8032 28260 8038 28262
rect 8094 28260 8118 28262
rect 8174 28260 8198 28262
rect 8254 28260 8278 28262
rect 8334 28260 8340 28262
rect 8032 28251 8340 28260
rect 7564 28076 7616 28082
rect 7564 28018 7616 28024
rect 7472 28008 7524 28014
rect 7472 27950 7524 27956
rect 7656 28008 7708 28014
rect 7656 27950 7708 27956
rect 7196 27600 7248 27606
rect 7196 27542 7248 27548
rect 7668 26926 7696 27950
rect 7932 27396 7984 27402
rect 7932 27338 7984 27344
rect 7656 26920 7708 26926
rect 7656 26862 7708 26868
rect 7012 26444 7064 26450
rect 7012 26386 7064 26392
rect 6552 25900 6604 25906
rect 6552 25842 6604 25848
rect 6920 25900 6972 25906
rect 6920 25842 6972 25848
rect 6736 25832 6788 25838
rect 6736 25774 6788 25780
rect 6748 25498 6776 25774
rect 6460 25492 6512 25498
rect 6460 25434 6512 25440
rect 6736 25492 6788 25498
rect 6736 25434 6788 25440
rect 6472 24954 6500 25434
rect 6460 24948 6512 24954
rect 6460 24890 6512 24896
rect 6748 24886 6776 25434
rect 6736 24880 6788 24886
rect 6736 24822 6788 24828
rect 6552 24812 6604 24818
rect 6552 24754 6604 24760
rect 6564 24342 6592 24754
rect 6828 24744 6880 24750
rect 6828 24686 6880 24692
rect 6552 24336 6604 24342
rect 6552 24278 6604 24284
rect 6840 24274 6868 24686
rect 6932 24682 6960 25842
rect 7024 25498 7052 26386
rect 7288 25900 7340 25906
rect 7288 25842 7340 25848
rect 7196 25696 7248 25702
rect 7196 25638 7248 25644
rect 7012 25492 7064 25498
rect 7012 25434 7064 25440
rect 6920 24676 6972 24682
rect 6920 24618 6972 24624
rect 6828 24268 6880 24274
rect 6828 24210 6880 24216
rect 6840 23186 6868 24210
rect 7024 24206 7052 25434
rect 7208 24206 7236 25638
rect 7300 25226 7328 25842
rect 7288 25220 7340 25226
rect 7288 25162 7340 25168
rect 7300 24682 7328 25162
rect 7472 25152 7524 25158
rect 7472 25094 7524 25100
rect 7484 24954 7512 25094
rect 7472 24948 7524 24954
rect 7472 24890 7524 24896
rect 7288 24676 7340 24682
rect 7288 24618 7340 24624
rect 7484 24342 7512 24890
rect 7668 24818 7696 26862
rect 7944 26042 7972 27338
rect 8032 27228 8340 27237
rect 8032 27226 8038 27228
rect 8094 27226 8118 27228
rect 8174 27226 8198 27228
rect 8254 27226 8278 27228
rect 8334 27226 8340 27228
rect 8094 27174 8096 27226
rect 8276 27174 8278 27226
rect 8032 27172 8038 27174
rect 8094 27172 8118 27174
rect 8174 27172 8198 27174
rect 8254 27172 8278 27174
rect 8334 27172 8340 27174
rect 8032 27163 8340 27172
rect 8496 26234 8524 29174
rect 8760 28960 8812 28966
rect 8760 28902 8812 28908
rect 8772 28626 8800 28902
rect 8760 28620 8812 28626
rect 8760 28562 8812 28568
rect 8576 28416 8628 28422
rect 8576 28358 8628 28364
rect 8588 28218 8616 28358
rect 8576 28212 8628 28218
rect 8576 28154 8628 28160
rect 9048 28082 9076 29582
rect 9404 29572 9456 29578
rect 9404 29514 9456 29520
rect 9416 29306 9444 29514
rect 9404 29300 9456 29306
rect 9404 29242 9456 29248
rect 9772 29232 9824 29238
rect 9772 29174 9824 29180
rect 9784 28762 9812 29174
rect 9772 28756 9824 28762
rect 9772 28698 9824 28704
rect 9404 28620 9456 28626
rect 9404 28562 9456 28568
rect 9416 28218 9444 28562
rect 9404 28212 9456 28218
rect 9404 28154 9456 28160
rect 9036 28076 9088 28082
rect 9036 28018 9088 28024
rect 9312 28076 9364 28082
rect 9312 28018 9364 28024
rect 9324 27674 9352 28018
rect 9772 28008 9824 28014
rect 9772 27950 9824 27956
rect 9312 27668 9364 27674
rect 9312 27610 9364 27616
rect 9784 27470 9812 27950
rect 9772 27464 9824 27470
rect 9772 27406 9824 27412
rect 8576 27328 8628 27334
rect 8576 27270 8628 27276
rect 8944 27328 8996 27334
rect 8944 27270 8996 27276
rect 8588 26926 8616 27270
rect 8956 27130 8984 27270
rect 9784 27130 9812 27406
rect 8944 27124 8996 27130
rect 8944 27066 8996 27072
rect 9772 27124 9824 27130
rect 9772 27066 9824 27072
rect 9220 26988 9272 26994
rect 9220 26930 9272 26936
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 8404 26206 8524 26234
rect 8032 26140 8340 26149
rect 8032 26138 8038 26140
rect 8094 26138 8118 26140
rect 8174 26138 8198 26140
rect 8254 26138 8278 26140
rect 8334 26138 8340 26140
rect 8094 26086 8096 26138
rect 8276 26086 8278 26138
rect 8032 26084 8038 26086
rect 8094 26084 8118 26086
rect 8174 26084 8198 26086
rect 8254 26084 8278 26086
rect 8334 26084 8340 26086
rect 8032 26075 8340 26084
rect 7932 26036 7984 26042
rect 7932 25978 7984 25984
rect 7748 25764 7800 25770
rect 7748 25706 7800 25712
rect 7760 25498 7788 25706
rect 7748 25492 7800 25498
rect 7748 25434 7800 25440
rect 8404 25294 8432 26206
rect 8588 25974 8616 26862
rect 9232 26382 9260 26930
rect 9220 26376 9272 26382
rect 9220 26318 9272 26324
rect 8576 25968 8628 25974
rect 8576 25910 8628 25916
rect 8760 25696 8812 25702
rect 8760 25638 8812 25644
rect 8772 25498 8800 25638
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 8392 25288 8444 25294
rect 8392 25230 8444 25236
rect 8032 25052 8340 25061
rect 8032 25050 8038 25052
rect 8094 25050 8118 25052
rect 8174 25050 8198 25052
rect 8254 25050 8278 25052
rect 8334 25050 8340 25052
rect 8094 24998 8096 25050
rect 8276 24998 8278 25050
rect 8032 24996 8038 24998
rect 8094 24996 8118 24998
rect 8174 24996 8198 24998
rect 8254 24996 8278 24998
rect 8334 24996 8340 24998
rect 8032 24987 8340 24996
rect 9232 24818 9260 26318
rect 9312 25288 9364 25294
rect 9312 25230 9364 25236
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 9220 24812 9272 24818
rect 9220 24754 9272 24760
rect 7656 24608 7708 24614
rect 7656 24550 7708 24556
rect 7472 24336 7524 24342
rect 7472 24278 7524 24284
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 7196 24200 7248 24206
rect 7196 24142 7248 24148
rect 7668 23866 7696 24550
rect 8032 23964 8340 23973
rect 8032 23962 8038 23964
rect 8094 23962 8118 23964
rect 8174 23962 8198 23964
rect 8254 23962 8278 23964
rect 8334 23962 8340 23964
rect 8094 23910 8096 23962
rect 8276 23910 8278 23962
rect 8032 23908 8038 23910
rect 8094 23908 8118 23910
rect 8174 23908 8198 23910
rect 8254 23908 8278 23910
rect 8334 23908 8340 23910
rect 8032 23899 8340 23908
rect 7656 23860 7708 23866
rect 7656 23802 7708 23808
rect 9324 23526 9352 25230
rect 9588 24812 9640 24818
rect 9588 24754 9640 24760
rect 9680 24812 9732 24818
rect 9680 24754 9732 24760
rect 9496 24064 9548 24070
rect 9496 24006 9548 24012
rect 9508 23798 9536 24006
rect 9496 23792 9548 23798
rect 9496 23734 9548 23740
rect 9312 23520 9364 23526
rect 9312 23462 9364 23468
rect 9324 23186 9352 23462
rect 6828 23180 6880 23186
rect 6828 23122 6880 23128
rect 9312 23180 9364 23186
rect 9312 23122 9364 23128
rect 6184 23112 6236 23118
rect 6184 23054 6236 23060
rect 6196 21690 6224 23054
rect 9220 23044 9272 23050
rect 9220 22986 9272 22992
rect 8032 22876 8340 22885
rect 8032 22874 8038 22876
rect 8094 22874 8118 22876
rect 8174 22874 8198 22876
rect 8254 22874 8278 22876
rect 8334 22874 8340 22876
rect 8094 22822 8096 22874
rect 8276 22822 8278 22874
rect 8032 22820 8038 22822
rect 8094 22820 8118 22822
rect 8174 22820 8198 22822
rect 8254 22820 8278 22822
rect 8334 22820 8340 22822
rect 8032 22811 8340 22820
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6932 22438 6960 22714
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8852 22636 8904 22642
rect 8852 22578 8904 22584
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 7288 22432 7340 22438
rect 7288 22374 7340 22380
rect 6368 22092 6420 22098
rect 6368 22034 6420 22040
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6380 21146 6408 22034
rect 6932 21593 6960 22374
rect 7300 22234 7328 22374
rect 7668 22234 7696 22510
rect 7748 22432 7800 22438
rect 7748 22374 7800 22380
rect 7288 22228 7340 22234
rect 7288 22170 7340 22176
rect 7656 22228 7708 22234
rect 7656 22170 7708 22176
rect 7288 22092 7340 22098
rect 7288 22034 7340 22040
rect 7300 22001 7328 22034
rect 7286 21992 7342 22001
rect 7286 21927 7342 21936
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 7116 21622 7144 21830
rect 7104 21616 7156 21622
rect 6918 21584 6974 21593
rect 7104 21558 7156 21564
rect 6918 21519 6974 21528
rect 6460 21344 6512 21350
rect 6460 21286 6512 21292
rect 6368 21140 6420 21146
rect 6368 21082 6420 21088
rect 6184 20936 6236 20942
rect 6184 20878 6236 20884
rect 6196 20602 6224 20878
rect 6184 20596 6236 20602
rect 6184 20538 6236 20544
rect 6196 16114 6224 20538
rect 6380 20398 6408 21082
rect 6368 20392 6420 20398
rect 6368 20334 6420 20340
rect 6380 18834 6408 20334
rect 6472 19854 6500 21286
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 6644 20392 6696 20398
rect 6644 20334 6696 20340
rect 6656 20058 6684 20334
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 6460 19848 6512 19854
rect 6460 19790 6512 19796
rect 6552 19780 6604 19786
rect 6552 19722 6604 19728
rect 6564 19378 6592 19722
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 6460 19236 6512 19242
rect 6460 19178 6512 19184
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6472 18766 6500 19178
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6276 18692 6328 18698
rect 6276 18634 6328 18640
rect 6288 18426 6316 18634
rect 6276 18420 6328 18426
rect 6276 18362 6328 18368
rect 6276 18284 6328 18290
rect 6276 18226 6328 18232
rect 6288 16250 6316 18226
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 6184 16108 6236 16114
rect 6184 16050 6236 16056
rect 6196 13870 6224 16050
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6288 12714 6316 16186
rect 6380 14074 6408 17478
rect 6472 16590 6500 18702
rect 6748 18290 6776 20878
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6932 19854 6960 20742
rect 7024 20602 7052 20878
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 7116 20534 7144 21558
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 7392 20942 7420 21286
rect 7668 20942 7696 22170
rect 7760 21418 7788 22374
rect 8128 22273 8156 22578
rect 8114 22264 8170 22273
rect 8680 22234 8708 22578
rect 8114 22199 8170 22208
rect 8668 22228 8720 22234
rect 8128 22166 8156 22199
rect 8668 22170 8720 22176
rect 8116 22160 8168 22166
rect 8116 22102 8168 22108
rect 8864 21962 8892 22578
rect 9232 22506 9260 22986
rect 9324 22642 9352 23122
rect 9312 22636 9364 22642
rect 9312 22578 9364 22584
rect 9600 22556 9628 24754
rect 9692 24410 9720 24754
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9680 24064 9732 24070
rect 9680 24006 9732 24012
rect 9692 22710 9720 24006
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 9600 22528 9812 22556
rect 9220 22500 9272 22506
rect 9220 22442 9272 22448
rect 9404 22432 9456 22438
rect 9456 22380 9536 22386
rect 9404 22374 9536 22380
rect 9416 22358 9536 22374
rect 9508 22094 9536 22358
rect 9416 22066 9536 22094
rect 9416 22030 9444 22066
rect 9404 22024 9456 22030
rect 9404 21966 9456 21972
rect 8392 21956 8444 21962
rect 8392 21898 8444 21904
rect 8852 21956 8904 21962
rect 8852 21898 8904 21904
rect 7840 21888 7892 21894
rect 7840 21830 7892 21836
rect 7748 21412 7800 21418
rect 7748 21354 7800 21360
rect 7380 20936 7432 20942
rect 7380 20878 7432 20884
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 7104 20256 7156 20262
rect 7104 20198 7156 20204
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 6840 18748 6868 19790
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 6920 18760 6972 18766
rect 6840 18720 6920 18748
rect 6920 18702 6972 18708
rect 6932 18290 6960 18702
rect 7024 18698 7052 19314
rect 7012 18692 7064 18698
rect 7012 18634 7064 18640
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 7024 18222 7052 18634
rect 6552 18216 6604 18222
rect 6552 18158 6604 18164
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 6564 16182 6592 18158
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 6932 16182 6960 16662
rect 6552 16176 6604 16182
rect 6552 16118 6604 16124
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 6564 15586 6592 16118
rect 6564 15558 6776 15586
rect 6644 15496 6696 15502
rect 6642 15464 6644 15473
rect 6696 15464 6698 15473
rect 6642 15399 6698 15408
rect 6656 15162 6684 15399
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 6276 12708 6328 12714
rect 6276 12650 6328 12656
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6196 12306 6224 12582
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6380 12102 6408 13738
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6460 13456 6512 13462
rect 6460 13398 6512 13404
rect 6472 12850 6500 13398
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6564 12782 6592 13670
rect 6656 13530 6684 13806
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6748 12918 6776 15558
rect 6932 15366 6960 16118
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6840 14618 6868 14894
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 7024 14482 7052 18158
rect 7116 18154 7144 20198
rect 7208 19854 7236 20198
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7300 18698 7328 19722
rect 7760 19446 7788 21354
rect 7852 21350 7880 21830
rect 8032 21788 8340 21797
rect 8032 21786 8038 21788
rect 8094 21786 8118 21788
rect 8174 21786 8198 21788
rect 8254 21786 8278 21788
rect 8334 21786 8340 21788
rect 8094 21734 8096 21786
rect 8276 21734 8278 21786
rect 8032 21732 8038 21734
rect 8094 21732 8118 21734
rect 8174 21732 8198 21734
rect 8254 21732 8278 21734
rect 8334 21732 8340 21734
rect 8032 21723 8340 21732
rect 7932 21684 7984 21690
rect 7932 21626 7984 21632
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 7748 19440 7800 19446
rect 7748 19382 7800 19388
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7288 18692 7340 18698
rect 7288 18634 7340 18640
rect 7104 18148 7156 18154
rect 7104 18090 7156 18096
rect 7116 18034 7144 18090
rect 7116 18006 7236 18034
rect 7102 17640 7158 17649
rect 7102 17575 7104 17584
rect 7156 17575 7158 17584
rect 7104 17546 7156 17552
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 7208 13326 7236 18006
rect 7300 17678 7328 18634
rect 7668 18290 7696 19314
rect 7852 19310 7880 19790
rect 7944 19378 7972 21626
rect 8404 21622 8432 21898
rect 9416 21894 9444 21966
rect 9496 21956 9548 21962
rect 9496 21898 9548 21904
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8576 21888 8628 21894
rect 8576 21830 8628 21836
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 8496 21622 8524 21830
rect 8392 21616 8444 21622
rect 8392 21558 8444 21564
rect 8484 21616 8536 21622
rect 8484 21558 8536 21564
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8220 21418 8248 21490
rect 8404 21457 8432 21558
rect 8588 21554 8616 21830
rect 8576 21548 8628 21554
rect 8576 21490 8628 21496
rect 8390 21448 8446 21457
rect 8208 21412 8260 21418
rect 8390 21383 8446 21392
rect 8208 21354 8260 21360
rect 8220 20890 8248 21354
rect 8588 21321 8616 21490
rect 8574 21312 8630 21321
rect 8574 21247 8630 21256
rect 8484 20936 8536 20942
rect 8220 20862 8432 20890
rect 8484 20878 8536 20884
rect 8032 20700 8340 20709
rect 8032 20698 8038 20700
rect 8094 20698 8118 20700
rect 8174 20698 8198 20700
rect 8254 20698 8278 20700
rect 8334 20698 8340 20700
rect 8094 20646 8096 20698
rect 8276 20646 8278 20698
rect 8032 20644 8038 20646
rect 8094 20644 8118 20646
rect 8174 20644 8198 20646
rect 8254 20644 8278 20646
rect 8334 20644 8340 20646
rect 8032 20635 8340 20644
rect 8404 20602 8432 20862
rect 8392 20596 8444 20602
rect 8392 20538 8444 20544
rect 8496 20534 8524 20878
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8484 20528 8536 20534
rect 8484 20470 8536 20476
rect 8484 20324 8536 20330
rect 8484 20266 8536 20272
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8220 20058 8248 20198
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 8032 19612 8340 19621
rect 8032 19610 8038 19612
rect 8094 19610 8118 19612
rect 8174 19610 8198 19612
rect 8254 19610 8278 19612
rect 8334 19610 8340 19612
rect 8094 19558 8096 19610
rect 8276 19558 8278 19610
rect 8032 19556 8038 19558
rect 8094 19556 8118 19558
rect 8174 19556 8198 19558
rect 8254 19556 8278 19558
rect 8334 19556 8340 19558
rect 8032 19547 8340 19556
rect 8496 19446 8524 20266
rect 8484 19440 8536 19446
rect 8484 19382 8536 19388
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 7840 19304 7892 19310
rect 7840 19246 7892 19252
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7852 18834 7880 19110
rect 7840 18828 7892 18834
rect 7840 18770 7892 18776
rect 8588 18766 8616 20742
rect 9404 19984 9456 19990
rect 9404 19926 9456 19932
rect 8852 19848 8904 19854
rect 8852 19790 8904 19796
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8864 19310 8892 19790
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 8956 18970 8984 19790
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 9232 18834 9260 19246
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9416 18766 9444 19926
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 7748 18692 7800 18698
rect 7748 18634 7800 18640
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 7576 17814 7604 18158
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7564 17808 7616 17814
rect 7564 17750 7616 17756
rect 7668 17678 7696 18022
rect 7760 17882 7788 18634
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 8032 18524 8340 18533
rect 8032 18522 8038 18524
rect 8094 18522 8118 18524
rect 8174 18522 8198 18524
rect 8254 18522 8278 18524
rect 8334 18522 8340 18524
rect 8094 18470 8096 18522
rect 8276 18470 8278 18522
rect 8032 18468 8038 18470
rect 8094 18468 8118 18470
rect 8174 18468 8198 18470
rect 8254 18468 8278 18470
rect 8334 18468 8340 18470
rect 8032 18459 8340 18468
rect 9324 18426 9352 18566
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7300 15314 7328 17614
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7472 16516 7524 16522
rect 7472 16458 7524 16464
rect 7484 16114 7512 16458
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7576 15570 7604 16186
rect 7760 16182 7788 16934
rect 7748 16176 7800 16182
rect 7748 16118 7800 16124
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7300 15286 7512 15314
rect 7484 15162 7512 15286
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6932 12442 6960 13262
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7116 12986 7144 13126
rect 7208 12986 7236 13126
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7300 12850 7328 13330
rect 7288 12844 7340 12850
rect 7208 12804 7288 12832
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 7208 12374 7236 12804
rect 7288 12786 7340 12792
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7208 12238 7236 12310
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 6368 12096 6420 12102
rect 6368 12038 6420 12044
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 6380 11830 6408 12038
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6472 10810 6500 11562
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6104 9710 6408 9738
rect 6012 9646 6224 9674
rect 5446 9616 5502 9625
rect 5502 9586 5580 9602
rect 5502 9580 5592 9586
rect 5502 9574 5540 9580
rect 5446 9551 5502 9560
rect 5540 9522 5592 9528
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5644 9178 5672 9318
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5460 8634 5488 9046
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5816 8560 5868 8566
rect 5446 8528 5502 8537
rect 5816 8502 5868 8508
rect 5446 8463 5448 8472
rect 5500 8463 5502 8472
rect 5448 8434 5500 8440
rect 5080 8366 5132 8372
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4066 7576 4122 7585
rect 4066 7511 4122 7520
rect 4491 7100 4799 7109
rect 4491 7098 4497 7100
rect 4553 7098 4577 7100
rect 4633 7098 4657 7100
rect 4713 7098 4737 7100
rect 4793 7098 4799 7100
rect 4553 7046 4555 7098
rect 4735 7046 4737 7098
rect 4491 7044 4497 7046
rect 4553 7044 4577 7046
rect 4633 7044 4657 7046
rect 4713 7044 4737 7046
rect 4793 7044 4799 7046
rect 4491 7035 4799 7044
rect 4620 6792 4672 6798
rect 4908 6780 4936 7754
rect 5000 7274 5028 7822
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 5000 6798 5028 6938
rect 5092 6798 5120 8366
rect 5184 8350 5304 8378
rect 5184 7818 5212 8350
rect 5264 8288 5316 8294
rect 5540 8288 5592 8294
rect 5264 8230 5316 8236
rect 5460 8236 5540 8242
rect 5460 8230 5592 8236
rect 5172 7812 5224 7818
rect 5172 7754 5224 7760
rect 5276 7546 5304 8230
rect 5460 8214 5580 8230
rect 5460 7954 5488 8214
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5828 7886 5856 8502
rect 5920 8430 5948 9386
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 6012 8566 6040 8910
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 6104 8634 6132 8774
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6000 8560 6052 8566
rect 6196 8514 6224 9646
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6288 8906 6316 9590
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 6000 8502 6052 8508
rect 6012 8430 6040 8502
rect 6104 8486 6224 8514
rect 6288 8498 6316 8842
rect 6380 8514 6408 9710
rect 6472 9704 6500 10746
rect 7024 10606 7052 12038
rect 7208 11898 7236 12174
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6552 9716 6604 9722
rect 6472 9676 6552 9704
rect 6472 8974 6500 9676
rect 6552 9658 6604 9664
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6932 9489 6960 9522
rect 6918 9480 6974 9489
rect 6552 9444 6604 9450
rect 6918 9415 6974 9424
rect 6552 9386 6604 9392
rect 6564 8974 6592 9386
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6472 8634 6500 8910
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6276 8492 6328 8498
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 5920 7970 5948 8366
rect 5920 7954 6040 7970
rect 5920 7948 6052 7954
rect 5920 7942 6000 7948
rect 6000 7890 6052 7896
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5828 7546 5856 7822
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 4672 6752 4936 6780
rect 4988 6792 5040 6798
rect 4620 6734 4672 6740
rect 4988 6734 5040 6740
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 3792 6248 3844 6254
rect 3792 6190 3844 6196
rect 4632 6118 4660 6734
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5092 6458 5120 6598
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5736 6254 5764 7278
rect 5920 6866 5948 7822
rect 6012 7274 6040 7890
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5920 6458 5948 6802
rect 6000 6792 6052 6798
rect 5998 6760 6000 6769
rect 6104 6780 6132 8486
rect 6380 8486 6500 8514
rect 6276 8434 6328 8440
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6196 7818 6224 8230
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6184 6792 6236 6798
rect 6052 6760 6054 6769
rect 6104 6752 6184 6780
rect 6184 6734 6236 6740
rect 5998 6695 6054 6704
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 6196 6322 6224 6734
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 6288 6458 6316 6666
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4491 6012 4799 6021
rect 4491 6010 4497 6012
rect 4553 6010 4577 6012
rect 4633 6010 4657 6012
rect 4713 6010 4737 6012
rect 4793 6010 4799 6012
rect 4553 5958 4555 6010
rect 4735 5958 4737 6010
rect 4491 5956 4497 5958
rect 4553 5956 4577 5958
rect 4633 5956 4657 5958
rect 4713 5956 4737 5958
rect 4793 5956 4799 5958
rect 4491 5947 4799 5956
rect 5368 5710 5396 6190
rect 5736 5846 5764 6190
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 6288 5234 6316 5714
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 4491 4924 4799 4933
rect 4491 4922 4497 4924
rect 4553 4922 4577 4924
rect 4633 4922 4657 4924
rect 4713 4922 4737 4924
rect 4793 4922 4799 4924
rect 4553 4870 4555 4922
rect 4735 4870 4737 4922
rect 4491 4868 4497 4870
rect 4553 4868 4577 4870
rect 4633 4868 4657 4870
rect 4713 4868 4737 4870
rect 4793 4868 4799 4870
rect 4491 4859 4799 4868
rect 6472 4486 6500 8486
rect 6656 8430 6684 9318
rect 7116 8906 7144 11018
rect 7208 10674 7236 11494
rect 7300 11286 7328 11698
rect 7392 11642 7420 14418
rect 7760 14346 7788 16118
rect 7852 14414 7880 18226
rect 8032 17436 8340 17445
rect 8032 17434 8038 17436
rect 8094 17434 8118 17436
rect 8174 17434 8198 17436
rect 8254 17434 8278 17436
rect 8334 17434 8340 17436
rect 8094 17382 8096 17434
rect 8276 17382 8278 17434
rect 8032 17380 8038 17382
rect 8094 17380 8118 17382
rect 8174 17380 8198 17382
rect 8254 17380 8278 17382
rect 8334 17380 8340 17382
rect 8032 17371 8340 17380
rect 8032 16348 8340 16357
rect 8032 16346 8038 16348
rect 8094 16346 8118 16348
rect 8174 16346 8198 16348
rect 8254 16346 8278 16348
rect 8334 16346 8340 16348
rect 8094 16294 8096 16346
rect 8276 16294 8278 16346
rect 8032 16292 8038 16294
rect 8094 16292 8118 16294
rect 8174 16292 8198 16294
rect 8254 16292 8278 16294
rect 8334 16292 8340 16294
rect 8032 16283 8340 16292
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 7944 15706 7972 16050
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 8220 15502 8248 15982
rect 8392 15972 8444 15978
rect 8392 15914 8444 15920
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 7944 15026 7972 15438
rect 8032 15260 8340 15269
rect 8032 15258 8038 15260
rect 8094 15258 8118 15260
rect 8174 15258 8198 15260
rect 8254 15258 8278 15260
rect 8334 15258 8340 15260
rect 8094 15206 8096 15258
rect 8276 15206 8278 15258
rect 8032 15204 8038 15206
rect 8094 15204 8118 15206
rect 8174 15204 8198 15206
rect 8254 15204 8278 15206
rect 8334 15204 8340 15206
rect 8032 15195 8340 15204
rect 8404 15026 8432 15914
rect 8680 15706 8708 15982
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8680 15162 8708 15642
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8128 14482 8156 14758
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 7840 14408 7892 14414
rect 7840 14350 7892 14356
rect 7748 14340 7800 14346
rect 7748 14282 7800 14288
rect 7852 14074 7880 14350
rect 8032 14172 8340 14181
rect 8032 14170 8038 14172
rect 8094 14170 8118 14172
rect 8174 14170 8198 14172
rect 8254 14170 8278 14172
rect 8334 14170 8340 14172
rect 8094 14118 8096 14170
rect 8276 14118 8278 14170
rect 8032 14116 8038 14118
rect 8094 14116 8118 14118
rect 8174 14116 8198 14118
rect 8254 14116 8278 14118
rect 8334 14116 8340 14118
rect 8032 14107 8340 14116
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7484 13190 7512 13806
rect 7564 13796 7616 13802
rect 7564 13738 7616 13744
rect 7576 13326 7604 13738
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7484 12306 7512 13126
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7576 12442 7604 12786
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7484 11898 7512 12242
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7392 11614 7512 11642
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7288 11280 7340 11286
rect 7288 11222 7340 11228
rect 7392 11150 7420 11494
rect 7484 11150 7512 11614
rect 7852 11150 7880 14010
rect 8588 13326 8616 14962
rect 9232 14958 9260 15438
rect 9416 15162 9444 18702
rect 9508 18154 9536 21898
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9692 20058 9720 20402
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 9600 19514 9628 19654
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9784 19446 9812 22528
rect 9876 21457 9904 30194
rect 13832 30122 13860 30246
rect 14188 30252 14240 30258
rect 14188 30194 14240 30200
rect 13820 30116 13872 30122
rect 13820 30058 13872 30064
rect 11574 29948 11882 29957
rect 11574 29946 11580 29948
rect 11636 29946 11660 29948
rect 11716 29946 11740 29948
rect 11796 29946 11820 29948
rect 11876 29946 11882 29948
rect 11636 29894 11638 29946
rect 11818 29894 11820 29946
rect 11574 29892 11580 29894
rect 11636 29892 11660 29894
rect 11716 29892 11740 29894
rect 11796 29892 11820 29894
rect 11876 29892 11882 29894
rect 11574 29883 11882 29892
rect 14096 29708 14148 29714
rect 14096 29650 14148 29656
rect 11336 29640 11388 29646
rect 11336 29582 11388 29588
rect 13268 29640 13320 29646
rect 13268 29582 13320 29588
rect 11060 29504 11112 29510
rect 11060 29446 11112 29452
rect 11244 29504 11296 29510
rect 11244 29446 11296 29452
rect 10416 28552 10468 28558
rect 10416 28494 10468 28500
rect 11072 28506 11100 29446
rect 11256 29306 11284 29446
rect 11244 29300 11296 29306
rect 11244 29242 11296 29248
rect 11244 29096 11296 29102
rect 11244 29038 11296 29044
rect 11152 28960 11204 28966
rect 11152 28902 11204 28908
rect 11164 28626 11192 28902
rect 11256 28626 11284 29038
rect 11152 28620 11204 28626
rect 11152 28562 11204 28568
rect 11244 28620 11296 28626
rect 11244 28562 11296 28568
rect 9956 28484 10008 28490
rect 9956 28426 10008 28432
rect 9968 28218 9996 28426
rect 9956 28212 10008 28218
rect 9956 28154 10008 28160
rect 9968 27470 9996 28154
rect 9956 27464 10008 27470
rect 9956 27406 10008 27412
rect 10428 26450 10456 28494
rect 11072 28490 11192 28506
rect 11072 28484 11204 28490
rect 11072 28478 11152 28484
rect 11152 28426 11204 28432
rect 11058 28112 11114 28121
rect 11058 28047 11114 28056
rect 11072 27674 11100 28047
rect 11060 27668 11112 27674
rect 11060 27610 11112 27616
rect 10784 27328 10836 27334
rect 10784 27270 10836 27276
rect 10796 27130 10824 27270
rect 10784 27124 10836 27130
rect 10784 27066 10836 27072
rect 11164 27062 11192 28426
rect 11256 28218 11284 28562
rect 11244 28212 11296 28218
rect 11244 28154 11296 28160
rect 11348 28082 11376 29582
rect 12256 29572 12308 29578
rect 12256 29514 12308 29520
rect 12268 29238 12296 29514
rect 13280 29306 13308 29582
rect 12624 29300 12676 29306
rect 12624 29242 12676 29248
rect 13268 29300 13320 29306
rect 13268 29242 13320 29248
rect 12256 29232 12308 29238
rect 12256 29174 12308 29180
rect 11574 28860 11882 28869
rect 11574 28858 11580 28860
rect 11636 28858 11660 28860
rect 11716 28858 11740 28860
rect 11796 28858 11820 28860
rect 11876 28858 11882 28860
rect 11636 28806 11638 28858
rect 11818 28806 11820 28858
rect 11574 28804 11580 28806
rect 11636 28804 11660 28806
rect 11716 28804 11740 28806
rect 11796 28804 11820 28806
rect 11876 28804 11882 28806
rect 11574 28795 11882 28804
rect 12636 28762 12664 29242
rect 13452 29096 13504 29102
rect 13452 29038 13504 29044
rect 13728 29096 13780 29102
rect 13728 29038 13780 29044
rect 12624 28756 12676 28762
rect 12624 28698 12676 28704
rect 12900 28756 12952 28762
rect 12900 28698 12952 28704
rect 12164 28416 12216 28422
rect 12164 28358 12216 28364
rect 12348 28416 12400 28422
rect 12348 28358 12400 28364
rect 12176 28218 12204 28358
rect 12164 28212 12216 28218
rect 12164 28154 12216 28160
rect 12360 28121 12388 28358
rect 12912 28218 12940 28698
rect 13360 28552 13412 28558
rect 13360 28494 13412 28500
rect 12900 28212 12952 28218
rect 12900 28154 12952 28160
rect 13084 28144 13136 28150
rect 12346 28112 12402 28121
rect 11336 28076 11388 28082
rect 11336 28018 11388 28024
rect 11980 28076 12032 28082
rect 13084 28086 13136 28092
rect 12346 28047 12402 28056
rect 11980 28018 12032 28024
rect 11348 27946 11376 28018
rect 11428 28008 11480 28014
rect 11428 27950 11480 27956
rect 11336 27940 11388 27946
rect 11336 27882 11388 27888
rect 11348 27674 11376 27882
rect 11336 27668 11388 27674
rect 11336 27610 11388 27616
rect 11440 27470 11468 27950
rect 11574 27772 11882 27781
rect 11574 27770 11580 27772
rect 11636 27770 11660 27772
rect 11716 27770 11740 27772
rect 11796 27770 11820 27772
rect 11876 27770 11882 27772
rect 11636 27718 11638 27770
rect 11818 27718 11820 27770
rect 11574 27716 11580 27718
rect 11636 27716 11660 27718
rect 11716 27716 11740 27718
rect 11796 27716 11820 27718
rect 11876 27716 11882 27718
rect 11574 27707 11882 27716
rect 11428 27464 11480 27470
rect 11428 27406 11480 27412
rect 11888 27464 11940 27470
rect 11992 27452 12020 28018
rect 12072 27872 12124 27878
rect 12072 27814 12124 27820
rect 12440 27872 12492 27878
rect 12440 27814 12492 27820
rect 12084 27470 12112 27814
rect 12452 27538 12480 27814
rect 13096 27538 13124 28086
rect 13372 27985 13400 28494
rect 13464 28082 13492 29038
rect 13740 28762 13768 29038
rect 13728 28756 13780 28762
rect 13728 28698 13780 28704
rect 13634 28656 13690 28665
rect 13634 28591 13636 28600
rect 13688 28591 13690 28600
rect 13636 28562 13688 28568
rect 14004 28552 14056 28558
rect 13634 28520 13690 28529
rect 14004 28494 14056 28500
rect 13634 28455 13636 28464
rect 13688 28455 13690 28464
rect 13636 28426 13688 28432
rect 13912 28416 13964 28422
rect 13832 28376 13912 28404
rect 13452 28076 13504 28082
rect 13452 28018 13504 28024
rect 13358 27976 13414 27985
rect 13358 27911 13414 27920
rect 13372 27674 13400 27911
rect 13360 27668 13412 27674
rect 13360 27610 13412 27616
rect 12440 27532 12492 27538
rect 12440 27474 12492 27480
rect 13084 27532 13136 27538
rect 13084 27474 13136 27480
rect 11940 27424 12020 27452
rect 11888 27406 11940 27412
rect 11520 27396 11572 27402
rect 11520 27338 11572 27344
rect 11152 27056 11204 27062
rect 11152 26998 11204 27004
rect 10416 26444 10468 26450
rect 10416 26386 10468 26392
rect 11164 26314 11192 26998
rect 11532 26926 11560 27338
rect 11992 27334 12020 27424
rect 12072 27464 12124 27470
rect 12072 27406 12124 27412
rect 11888 27328 11940 27334
rect 11888 27270 11940 27276
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 11900 26926 11928 27270
rect 12256 26988 12308 26994
rect 12256 26930 12308 26936
rect 11520 26920 11572 26926
rect 11520 26862 11572 26868
rect 11888 26920 11940 26926
rect 11888 26862 11940 26868
rect 11244 26784 11296 26790
rect 11244 26726 11296 26732
rect 11256 26586 11284 26726
rect 11574 26684 11882 26693
rect 11574 26682 11580 26684
rect 11636 26682 11660 26684
rect 11716 26682 11740 26684
rect 11796 26682 11820 26684
rect 11876 26682 11882 26684
rect 11636 26630 11638 26682
rect 11818 26630 11820 26682
rect 11574 26628 11580 26630
rect 11636 26628 11660 26630
rect 11716 26628 11740 26630
rect 11796 26628 11820 26630
rect 11876 26628 11882 26630
rect 11574 26619 11882 26628
rect 11244 26580 11296 26586
rect 11244 26522 11296 26528
rect 12268 26450 12296 26930
rect 12452 26926 12480 27474
rect 12808 27464 12860 27470
rect 12808 27406 12860 27412
rect 12532 27328 12584 27334
rect 12532 27270 12584 27276
rect 12440 26920 12492 26926
rect 12440 26862 12492 26868
rect 12544 26586 12572 27270
rect 12820 27062 12848 27406
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 12808 27056 12860 27062
rect 12808 26998 12860 27004
rect 12728 26874 12756 26998
rect 12728 26846 12848 26874
rect 12820 26790 12848 26846
rect 12808 26784 12860 26790
rect 12808 26726 12860 26732
rect 12532 26580 12584 26586
rect 12532 26522 12584 26528
rect 11428 26444 11480 26450
rect 11428 26386 11480 26392
rect 12256 26444 12308 26450
rect 12256 26386 12308 26392
rect 11152 26308 11204 26314
rect 11152 26250 11204 26256
rect 11440 24818 11468 26386
rect 11574 25596 11882 25605
rect 11574 25594 11580 25596
rect 11636 25594 11660 25596
rect 11716 25594 11740 25596
rect 11796 25594 11820 25596
rect 11876 25594 11882 25596
rect 11636 25542 11638 25594
rect 11818 25542 11820 25594
rect 11574 25540 11580 25542
rect 11636 25540 11660 25542
rect 11716 25540 11740 25542
rect 11796 25540 11820 25542
rect 11876 25540 11882 25542
rect 11574 25531 11882 25540
rect 13464 25294 13492 28018
rect 13636 27124 13688 27130
rect 13636 27066 13688 27072
rect 13648 27010 13676 27066
rect 13832 27010 13860 28376
rect 13912 28358 13964 28364
rect 14016 27674 14044 28494
rect 14004 27668 14056 27674
rect 14004 27610 14056 27616
rect 14004 27532 14056 27538
rect 14004 27474 14056 27480
rect 14016 27334 14044 27474
rect 14004 27328 14056 27334
rect 14004 27270 14056 27276
rect 13648 26982 13860 27010
rect 13912 26988 13964 26994
rect 13912 26930 13964 26936
rect 13924 26858 13952 26930
rect 13912 26852 13964 26858
rect 13912 26794 13964 26800
rect 12992 25288 13044 25294
rect 12992 25230 13044 25236
rect 13452 25288 13504 25294
rect 13452 25230 13504 25236
rect 11888 25152 11940 25158
rect 11888 25094 11940 25100
rect 11900 24886 11928 25094
rect 11888 24880 11940 24886
rect 11888 24822 11940 24828
rect 11428 24812 11480 24818
rect 11428 24754 11480 24760
rect 11336 24744 11388 24750
rect 11336 24686 11388 24692
rect 10416 24608 10468 24614
rect 10416 24550 10468 24556
rect 10048 24200 10100 24206
rect 10048 24142 10100 24148
rect 10060 23322 10088 24142
rect 10048 23316 10100 23322
rect 10048 23258 10100 23264
rect 10232 22772 10284 22778
rect 10232 22714 10284 22720
rect 9956 22568 10008 22574
rect 10244 22522 10272 22714
rect 9956 22510 10008 22516
rect 9968 22098 9996 22510
rect 10152 22494 10272 22522
rect 9956 22092 10008 22098
rect 9956 22034 10008 22040
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 9862 21448 9918 21457
rect 9862 21383 9918 21392
rect 9968 20874 9996 21626
rect 10048 20936 10100 20942
rect 10048 20878 10100 20884
rect 10152 20890 10180 22494
rect 10232 22432 10284 22438
rect 10232 22374 10284 22380
rect 10244 21962 10272 22374
rect 10232 21956 10284 21962
rect 10232 21898 10284 21904
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 9956 20868 10008 20874
rect 9956 20810 10008 20816
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 9876 20369 9904 20402
rect 9862 20360 9918 20369
rect 9862 20295 9918 20304
rect 9772 19440 9824 19446
rect 9772 19382 9824 19388
rect 9876 19378 9904 20295
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9588 19236 9640 19242
rect 9588 19178 9640 19184
rect 9600 18970 9628 19178
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9968 18834 9996 20810
rect 10060 19854 10088 20878
rect 10152 20862 10272 20890
rect 10140 20800 10192 20806
rect 10140 20742 10192 20748
rect 10152 20466 10180 20742
rect 10244 20534 10272 20862
rect 10232 20528 10284 20534
rect 10232 20470 10284 20476
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 10152 19417 10180 19654
rect 10138 19408 10194 19417
rect 10138 19343 10194 19352
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9692 18290 9720 18362
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9496 18148 9548 18154
rect 9496 18090 9548 18096
rect 9784 17762 9812 18226
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9692 17734 9812 17762
rect 9692 16590 9720 17734
rect 9876 17134 9904 18022
rect 9968 17746 9996 18770
rect 10244 18290 10272 20470
rect 10336 20330 10364 21422
rect 10428 20618 10456 24550
rect 11348 23798 11376 24686
rect 10784 23792 10836 23798
rect 10704 23752 10784 23780
rect 10508 23316 10560 23322
rect 10508 23258 10560 23264
rect 10520 22030 10548 23258
rect 10704 23118 10732 23752
rect 10784 23734 10836 23740
rect 11336 23792 11388 23798
rect 11336 23734 11388 23740
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10598 22264 10654 22273
rect 10598 22199 10600 22208
rect 10652 22199 10654 22208
rect 10600 22170 10652 22176
rect 10796 22030 10824 23462
rect 11440 23186 11468 24754
rect 11574 24508 11882 24517
rect 11574 24506 11580 24508
rect 11636 24506 11660 24508
rect 11716 24506 11740 24508
rect 11796 24506 11820 24508
rect 11876 24506 11882 24508
rect 11636 24454 11638 24506
rect 11818 24454 11820 24506
rect 11574 24452 11580 24454
rect 11636 24452 11660 24454
rect 11716 24452 11740 24454
rect 11796 24452 11820 24454
rect 11876 24452 11882 24454
rect 11574 24443 11882 24452
rect 11888 24132 11940 24138
rect 11888 24074 11940 24080
rect 11900 23866 11928 24074
rect 13004 23866 13032 25230
rect 13544 24744 13596 24750
rect 13544 24686 13596 24692
rect 13452 24132 13504 24138
rect 13452 24074 13504 24080
rect 11888 23860 11940 23866
rect 11888 23802 11940 23808
rect 12992 23860 13044 23866
rect 12992 23802 13044 23808
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 11574 23420 11882 23429
rect 11574 23418 11580 23420
rect 11636 23418 11660 23420
rect 11716 23418 11740 23420
rect 11796 23418 11820 23420
rect 11876 23418 11882 23420
rect 11636 23366 11638 23418
rect 11818 23366 11820 23418
rect 11574 23364 11580 23366
rect 11636 23364 11660 23366
rect 11716 23364 11740 23366
rect 11796 23364 11820 23366
rect 11876 23364 11882 23366
rect 11574 23355 11882 23364
rect 11428 23180 11480 23186
rect 11428 23122 11480 23128
rect 10876 23112 10928 23118
rect 10876 23054 10928 23060
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10784 22024 10836 22030
rect 10784 21966 10836 21972
rect 10600 21956 10652 21962
rect 10600 21898 10652 21904
rect 10692 21956 10744 21962
rect 10692 21898 10744 21904
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 10520 21078 10548 21830
rect 10508 21072 10560 21078
rect 10508 21014 10560 21020
rect 10428 20590 10548 20618
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 10324 20324 10376 20330
rect 10324 20266 10376 20272
rect 10428 20210 10456 20402
rect 10336 20182 10456 20210
rect 10232 18284 10284 18290
rect 10232 18226 10284 18232
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9968 17338 9996 17682
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 9232 14414 9260 14894
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8032 13084 8340 13093
rect 8032 13082 8038 13084
rect 8094 13082 8118 13084
rect 8174 13082 8198 13084
rect 8254 13082 8278 13084
rect 8334 13082 8340 13084
rect 8094 13030 8096 13082
rect 8276 13030 8278 13082
rect 8032 13028 8038 13030
rect 8094 13028 8118 13030
rect 8174 13028 8198 13030
rect 8254 13028 8278 13030
rect 8334 13028 8340 13030
rect 8032 13019 8340 13028
rect 9232 12782 9260 14350
rect 9416 13190 9444 15098
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9232 12306 9260 12718
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9600 12102 9628 15370
rect 9692 13462 9720 16526
rect 9876 15978 9904 16526
rect 10060 16522 10088 18022
rect 10152 17610 10180 18022
rect 10140 17604 10192 17610
rect 10140 17546 10192 17552
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9968 16096 9996 16390
rect 10060 16266 10088 16458
rect 10244 16454 10272 18226
rect 10336 18222 10364 20182
rect 10414 19952 10470 19961
rect 10414 19887 10470 19896
rect 10428 19786 10456 19887
rect 10416 19780 10468 19786
rect 10416 19722 10468 19728
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10060 16238 10272 16266
rect 10048 16108 10100 16114
rect 9968 16068 10048 16096
rect 10048 16050 10100 16056
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 9864 15972 9916 15978
rect 9864 15914 9916 15920
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9968 15706 9996 15846
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9956 15428 10008 15434
rect 9956 15370 10008 15376
rect 9968 15094 9996 15370
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 9968 13870 9996 15030
rect 10060 13938 10088 16050
rect 10152 15978 10180 16050
rect 10140 15972 10192 15978
rect 10140 15914 10192 15920
rect 10152 15570 10180 15914
rect 10140 15564 10192 15570
rect 10140 15506 10192 15512
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 10152 13977 10180 14486
rect 10138 13968 10194 13977
rect 10048 13932 10100 13938
rect 10138 13903 10194 13912
rect 10048 13874 10100 13880
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9680 13456 9732 13462
rect 9678 13424 9680 13433
rect 9772 13456 9824 13462
rect 9732 13424 9734 13433
rect 9772 13398 9824 13404
rect 9968 13410 9996 13806
rect 10244 13734 10272 16238
rect 10336 16114 10364 18158
rect 10520 16454 10548 20590
rect 10612 20534 10640 21898
rect 10704 21146 10732 21898
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10692 21140 10744 21146
rect 10692 21082 10744 21088
rect 10796 21010 10824 21286
rect 10784 21004 10836 21010
rect 10784 20946 10836 20952
rect 10796 20806 10824 20946
rect 10888 20942 10916 23054
rect 12176 22642 12204 23462
rect 12820 22778 12848 23666
rect 12808 22772 12860 22778
rect 12808 22714 12860 22720
rect 12532 22704 12584 22710
rect 12532 22646 12584 22652
rect 10968 22636 11020 22642
rect 10968 22578 11020 22584
rect 12164 22636 12216 22642
rect 12164 22578 12216 22584
rect 10980 21894 11008 22578
rect 11428 22568 11480 22574
rect 11428 22510 11480 22516
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 10968 21888 11020 21894
rect 10968 21830 11020 21836
rect 10980 21622 11008 21830
rect 10968 21616 11020 21622
rect 10968 21558 11020 21564
rect 11164 21468 11192 22170
rect 10980 21440 11192 21468
rect 10876 20936 10928 20942
rect 10876 20878 10928 20884
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 10600 20528 10652 20534
rect 10600 20470 10652 20476
rect 10980 20466 11008 21440
rect 11440 21128 11468 22510
rect 11574 22332 11882 22341
rect 11574 22330 11580 22332
rect 11636 22330 11660 22332
rect 11716 22330 11740 22332
rect 11796 22330 11820 22332
rect 11876 22330 11882 22332
rect 11636 22278 11638 22330
rect 11818 22278 11820 22330
rect 11574 22276 11580 22278
rect 11636 22276 11660 22278
rect 11716 22276 11740 22278
rect 11796 22276 11820 22278
rect 11876 22276 11882 22278
rect 11574 22267 11882 22276
rect 12544 22166 12572 22646
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 12636 22234 12664 22578
rect 12624 22228 12676 22234
rect 12624 22170 12676 22176
rect 12532 22160 12584 22166
rect 12532 22102 12584 22108
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 11574 21244 11882 21253
rect 11574 21242 11580 21244
rect 11636 21242 11660 21244
rect 11716 21242 11740 21244
rect 11796 21242 11820 21244
rect 11876 21242 11882 21244
rect 11636 21190 11638 21242
rect 11818 21190 11820 21242
rect 11574 21188 11580 21190
rect 11636 21188 11660 21190
rect 11716 21188 11740 21190
rect 11796 21188 11820 21190
rect 11876 21188 11882 21190
rect 11574 21179 11882 21188
rect 11440 21100 11560 21128
rect 11532 20942 11560 21100
rect 11796 21004 11848 21010
rect 11796 20946 11848 20952
rect 11428 20936 11480 20942
rect 11428 20878 11480 20884
rect 11520 20936 11572 20942
rect 11520 20878 11572 20884
rect 11152 20868 11204 20874
rect 11152 20810 11204 20816
rect 11164 20466 11192 20810
rect 11242 20632 11298 20641
rect 11242 20567 11244 20576
rect 11296 20567 11298 20576
rect 11244 20538 11296 20544
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 10876 19780 10928 19786
rect 10876 19722 10928 19728
rect 10888 19446 10916 19722
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11072 19514 11100 19654
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 10876 19440 10928 19446
rect 10876 19382 10928 19388
rect 11164 18834 11192 19654
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 10704 18086 10732 18566
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 11072 17882 11100 18566
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 11336 18216 11388 18222
rect 11336 18158 11388 18164
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11072 17134 11100 17818
rect 11256 17678 11284 18158
rect 11348 17882 11376 18158
rect 11336 17876 11388 17882
rect 11336 17818 11388 17824
rect 11440 17678 11468 20878
rect 11808 20466 11836 20946
rect 11992 20806 12020 21966
rect 12072 21888 12124 21894
rect 12072 21830 12124 21836
rect 12084 21554 12112 21830
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 11980 20800 12032 20806
rect 11980 20742 12032 20748
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11574 20156 11882 20165
rect 11574 20154 11580 20156
rect 11636 20154 11660 20156
rect 11716 20154 11740 20156
rect 11796 20154 11820 20156
rect 11876 20154 11882 20156
rect 11636 20102 11638 20154
rect 11818 20102 11820 20154
rect 11574 20100 11580 20102
rect 11636 20100 11660 20102
rect 11716 20100 11740 20102
rect 11796 20100 11820 20102
rect 11876 20100 11882 20102
rect 11574 20091 11882 20100
rect 11574 19068 11882 19077
rect 11574 19066 11580 19068
rect 11636 19066 11660 19068
rect 11716 19066 11740 19068
rect 11796 19066 11820 19068
rect 11876 19066 11882 19068
rect 11636 19014 11638 19066
rect 11818 19014 11820 19066
rect 11574 19012 11580 19014
rect 11636 19012 11660 19014
rect 11716 19012 11740 19014
rect 11796 19012 11820 19014
rect 11876 19012 11882 19014
rect 11574 19003 11882 19012
rect 11574 17980 11882 17989
rect 11574 17978 11580 17980
rect 11636 17978 11660 17980
rect 11716 17978 11740 17980
rect 11796 17978 11820 17980
rect 11876 17978 11882 17980
rect 11636 17926 11638 17978
rect 11818 17926 11820 17978
rect 11574 17924 11580 17926
rect 11636 17924 11660 17926
rect 11716 17924 11740 17926
rect 11796 17924 11820 17926
rect 11876 17924 11882 17926
rect 11574 17915 11882 17924
rect 11992 17678 12020 20742
rect 12072 20392 12124 20398
rect 12072 20334 12124 20340
rect 12084 20058 12112 20334
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 12072 19848 12124 19854
rect 12070 19816 12072 19825
rect 12124 19816 12126 19825
rect 12070 19751 12126 19760
rect 12176 19310 12204 21490
rect 12544 21026 12572 22102
rect 13464 22094 13492 24074
rect 13556 23662 13584 24686
rect 13924 24206 13952 26794
rect 14108 24886 14136 29650
rect 14096 24880 14148 24886
rect 14096 24822 14148 24828
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 13556 23118 13584 23598
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 14004 23112 14056 23118
rect 14004 23054 14056 23060
rect 13912 23044 13964 23050
rect 13912 22986 13964 22992
rect 13924 22506 13952 22986
rect 13912 22500 13964 22506
rect 13912 22442 13964 22448
rect 13464 22066 13768 22094
rect 13740 21978 13768 22066
rect 12624 21956 12676 21962
rect 12624 21898 12676 21904
rect 13360 21956 13412 21962
rect 13360 21898 13412 21904
rect 13648 21950 13768 21978
rect 12636 21554 12664 21898
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12624 21344 12676 21350
rect 12624 21286 12676 21292
rect 12636 21146 12664 21286
rect 12624 21140 12676 21146
rect 12624 21082 12676 21088
rect 12544 20998 12664 21026
rect 12636 20913 12664 20998
rect 12622 20904 12678 20913
rect 12622 20839 12678 20848
rect 12348 20528 12400 20534
rect 12400 20488 12480 20516
rect 12348 20470 12400 20476
rect 12360 19854 12388 20470
rect 12452 20398 12480 20488
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12268 19514 12296 19654
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 12452 19334 12480 19926
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12544 19514 12572 19790
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12360 19306 12480 19334
rect 12176 18970 12204 19246
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12360 18698 12388 19306
rect 12544 18834 12572 19450
rect 12636 19446 12664 20839
rect 12624 19440 12676 19446
rect 12624 19382 12676 19388
rect 12728 19174 12756 21422
rect 12912 20874 12940 21830
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 12992 21344 13044 21350
rect 12992 21286 13044 21292
rect 12900 20868 12952 20874
rect 12900 20810 12952 20816
rect 12808 20528 12860 20534
rect 12912 20516 12940 20810
rect 12860 20488 12940 20516
rect 12808 20470 12860 20476
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12636 18902 12664 19110
rect 12820 18970 12848 20470
rect 13004 19854 13032 21286
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 13188 19854 13216 20198
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12912 19378 12940 19654
rect 13188 19378 13216 19790
rect 13280 19514 13308 21422
rect 13372 21026 13400 21898
rect 13648 21894 13676 21950
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 13648 21622 13676 21830
rect 13636 21616 13688 21622
rect 13636 21558 13688 21564
rect 13452 21072 13504 21078
rect 13372 21020 13452 21026
rect 13372 21014 13504 21020
rect 13372 20998 13492 21014
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12624 18896 12676 18902
rect 12624 18838 12676 18844
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12348 18692 12400 18698
rect 12268 18652 12348 18680
rect 12268 18578 12296 18652
rect 12348 18634 12400 18640
rect 12176 18550 12296 18578
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11428 17672 11480 17678
rect 11980 17672 12032 17678
rect 11428 17614 11480 17620
rect 11900 17632 11980 17660
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10336 13938 10364 16050
rect 10428 15162 10456 16390
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10520 15609 10548 15982
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10506 15600 10562 15609
rect 10506 15535 10562 15544
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10508 14952 10560 14958
rect 10428 14912 10508 14940
rect 10428 14414 10456 14912
rect 10508 14894 10560 14900
rect 10796 14414 10824 15642
rect 10980 15162 11008 16594
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 11072 15706 11100 15982
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10428 13818 10456 14350
rect 10692 14340 10744 14346
rect 10692 14282 10744 14288
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10336 13790 10456 13818
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 9678 13359 9734 13368
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 8032 11996 8340 12005
rect 8032 11994 8038 11996
rect 8094 11994 8118 11996
rect 8174 11994 8198 11996
rect 8254 11994 8278 11996
rect 8334 11994 8340 11996
rect 8094 11942 8096 11994
rect 8276 11942 8278 11994
rect 8032 11940 8038 11942
rect 8094 11940 8118 11942
rect 8174 11940 8198 11942
rect 8254 11940 8278 11942
rect 8334 11940 8340 11942
rect 8032 11931 8340 11940
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7484 9674 7512 11086
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7668 10742 7696 10950
rect 7656 10736 7708 10742
rect 7656 10678 7708 10684
rect 7484 9646 7604 9674
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6748 8430 6776 8570
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6748 8022 6776 8366
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6840 7818 6868 8434
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6564 7546 6592 7686
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6564 5914 6592 6598
rect 6840 6390 6868 6734
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6932 5778 6960 6598
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 7012 5636 7064 5642
rect 7116 5624 7144 8842
rect 7208 7954 7236 9318
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7208 6322 7236 7686
rect 7576 6934 7604 9646
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7208 5914 7236 6258
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7064 5596 7144 5624
rect 7012 5578 7064 5584
rect 7116 5302 7144 5596
rect 7300 5370 7328 6802
rect 7576 6798 7604 6870
rect 7852 6798 7880 11086
rect 8956 11082 8984 11630
rect 9692 11286 9720 13262
rect 9784 12170 9812 13398
rect 9968 13382 10180 13410
rect 9968 12918 9996 13382
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 10060 12782 10088 13194
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10060 12434 10088 12718
rect 9968 12406 10088 12434
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 9876 11830 9904 12038
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8032 10908 8340 10917
rect 8032 10906 8038 10908
rect 8094 10906 8118 10908
rect 8174 10906 8198 10908
rect 8254 10906 8278 10908
rect 8334 10906 8340 10908
rect 8094 10854 8096 10906
rect 8276 10854 8278 10906
rect 8032 10852 8038 10854
rect 8094 10852 8118 10854
rect 8174 10852 8198 10854
rect 8254 10852 8278 10854
rect 8334 10852 8340 10854
rect 8032 10843 8340 10852
rect 8032 9820 8340 9829
rect 8032 9818 8038 9820
rect 8094 9818 8118 9820
rect 8174 9818 8198 9820
rect 8254 9818 8278 9820
rect 8334 9818 8340 9820
rect 8094 9766 8096 9818
rect 8276 9766 8278 9818
rect 8032 9764 8038 9766
rect 8094 9764 8118 9766
rect 8174 9764 8198 9766
rect 8254 9764 8278 9766
rect 8334 9764 8340 9766
rect 8032 9755 8340 9764
rect 8852 9512 8904 9518
rect 8850 9480 8852 9489
rect 8904 9480 8906 9489
rect 8850 9415 8906 9424
rect 8956 8974 8984 11018
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9048 9586 9076 9862
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9140 9042 9168 9454
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8032 8732 8340 8741
rect 8032 8730 8038 8732
rect 8094 8730 8118 8732
rect 8174 8730 8198 8732
rect 8254 8730 8278 8732
rect 8334 8730 8340 8732
rect 8094 8678 8096 8730
rect 8276 8678 8278 8730
rect 8032 8676 8038 8678
rect 8094 8676 8118 8678
rect 8174 8676 8198 8678
rect 8254 8676 8278 8678
rect 8334 8676 8340 8678
rect 8032 8667 8340 8676
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7564 6792 7616 6798
rect 7840 6792 7892 6798
rect 7564 6734 7616 6740
rect 7746 6760 7802 6769
rect 7392 6186 7420 6734
rect 7484 6458 7512 6734
rect 7840 6734 7892 6740
rect 7746 6695 7748 6704
rect 7800 6695 7802 6704
rect 7748 6666 7800 6672
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7576 6118 7604 6598
rect 7852 6186 7880 6734
rect 7944 6322 7972 8366
rect 8032 7644 8340 7653
rect 8032 7642 8038 7644
rect 8094 7642 8118 7644
rect 8174 7642 8198 7644
rect 8254 7642 8278 7644
rect 8334 7642 8340 7644
rect 8094 7590 8096 7642
rect 8276 7590 8278 7642
rect 8032 7588 8038 7590
rect 8094 7588 8118 7590
rect 8174 7588 8198 7590
rect 8254 7588 8278 7590
rect 8334 7588 8340 7590
rect 8032 7579 8340 7588
rect 8032 6556 8340 6565
rect 8032 6554 8038 6556
rect 8094 6554 8118 6556
rect 8174 6554 8198 6556
rect 8254 6554 8278 6556
rect 8334 6554 8340 6556
rect 8094 6502 8096 6554
rect 8276 6502 8278 6554
rect 8032 6500 8038 6502
rect 8094 6500 8118 6502
rect 8174 6500 8198 6502
rect 8254 6500 8278 6502
rect 8334 6500 8340 6502
rect 8032 6491 8340 6500
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 7840 6180 7892 6186
rect 7840 6122 7892 6128
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7576 5846 7604 6054
rect 7564 5840 7616 5846
rect 7564 5782 7616 5788
rect 7944 5370 7972 6258
rect 8032 5468 8340 5477
rect 8032 5466 8038 5468
rect 8094 5466 8118 5468
rect 8174 5466 8198 5468
rect 8254 5466 8278 5468
rect 8334 5466 8340 5468
rect 8094 5414 8096 5466
rect 8276 5414 8278 5466
rect 8032 5412 8038 5414
rect 8094 5412 8118 5414
rect 8174 5412 8198 5414
rect 8254 5412 8278 5414
rect 8334 5412 8340 5414
rect 8032 5403 8340 5412
rect 8956 5370 8984 8910
rect 9036 8560 9088 8566
rect 9034 8528 9036 8537
rect 9088 8528 9090 8537
rect 9034 8463 9090 8472
rect 9600 8430 9628 10066
rect 9692 9518 9720 11222
rect 9784 10810 9812 11630
rect 9968 10962 9996 12406
rect 10152 12186 10180 13382
rect 10244 13190 10272 13670
rect 10336 13326 10364 13790
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 10428 12986 10456 13670
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10520 12782 10548 13262
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10244 12442 10272 12718
rect 10508 12640 10560 12646
rect 10336 12600 10508 12628
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 10060 12170 10180 12186
rect 10048 12164 10180 12170
rect 10100 12158 10180 12164
rect 10048 12106 10100 12112
rect 9876 10934 9996 10962
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9784 10266 9812 10610
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9876 10146 9904 10934
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9784 10130 9904 10146
rect 9772 10124 9904 10130
rect 9824 10118 9904 10124
rect 9772 10066 9824 10072
rect 9876 9926 9904 10118
rect 9968 10062 9996 10746
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9968 9722 9996 9998
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9692 8498 9720 9454
rect 9784 9353 9812 9454
rect 9770 9344 9826 9353
rect 9770 9279 9826 9288
rect 9876 9042 9904 9522
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 10060 8906 10088 12106
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10152 10266 10180 10610
rect 10244 10470 10272 11834
rect 10336 10674 10364 12600
rect 10508 12582 10560 12588
rect 10414 12200 10470 12209
rect 10612 12186 10640 13874
rect 10704 13258 10732 14282
rect 10980 14278 11008 15098
rect 11164 14346 11192 17546
rect 11256 17066 11284 17614
rect 11336 17264 11388 17270
rect 11336 17206 11388 17212
rect 11244 17060 11296 17066
rect 11244 17002 11296 17008
rect 11348 15042 11376 17206
rect 11256 15014 11376 15042
rect 11440 15026 11468 17614
rect 11900 17270 11928 17632
rect 11980 17614 12032 17620
rect 12084 17490 12112 18022
rect 11992 17462 12112 17490
rect 11888 17264 11940 17270
rect 11888 17206 11940 17212
rect 11574 16892 11882 16901
rect 11574 16890 11580 16892
rect 11636 16890 11660 16892
rect 11716 16890 11740 16892
rect 11796 16890 11820 16892
rect 11876 16890 11882 16892
rect 11636 16838 11638 16890
rect 11818 16838 11820 16890
rect 11574 16836 11580 16838
rect 11636 16836 11660 16838
rect 11716 16836 11740 16838
rect 11796 16836 11820 16838
rect 11876 16836 11882 16838
rect 11574 16827 11882 16836
rect 11574 15804 11882 15813
rect 11574 15802 11580 15804
rect 11636 15802 11660 15804
rect 11716 15802 11740 15804
rect 11796 15802 11820 15804
rect 11876 15802 11882 15804
rect 11636 15750 11638 15802
rect 11818 15750 11820 15802
rect 11574 15748 11580 15750
rect 11636 15748 11660 15750
rect 11716 15748 11740 15750
rect 11796 15748 11820 15750
rect 11876 15748 11882 15750
rect 11574 15739 11882 15748
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11716 15094 11744 15642
rect 11796 15428 11848 15434
rect 11796 15370 11848 15376
rect 11808 15094 11836 15370
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 11796 15088 11848 15094
rect 11848 15048 11928 15076
rect 11796 15030 11848 15036
rect 11428 15020 11480 15026
rect 11256 14414 11284 15014
rect 11428 14962 11480 14968
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11348 14482 11376 14894
rect 11428 14884 11480 14890
rect 11428 14826 11480 14832
rect 11440 14618 11468 14826
rect 11900 14804 11928 15048
rect 11992 14906 12020 17462
rect 12176 15706 12204 18550
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12164 15700 12216 15706
rect 12164 15642 12216 15648
rect 12268 15502 12296 16526
rect 12348 16448 12400 16454
rect 12348 16390 12400 16396
rect 12360 15978 12388 16390
rect 12348 15972 12400 15978
rect 12348 15914 12400 15920
rect 12256 15496 12308 15502
rect 12544 15450 12572 18770
rect 12716 18760 12768 18766
rect 12636 18708 12716 18714
rect 12636 18702 12768 18708
rect 12636 18686 12756 18702
rect 12636 18426 12664 18686
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12728 18426 12756 18566
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12636 17882 12664 18226
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12820 17338 12848 18566
rect 12912 18290 12940 19110
rect 13176 18964 13228 18970
rect 13176 18906 13228 18912
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12636 15570 12664 16050
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12256 15438 12308 15444
rect 11992 14878 12112 14906
rect 11900 14776 12020 14804
rect 11574 14716 11882 14725
rect 11574 14714 11580 14716
rect 11636 14714 11660 14716
rect 11716 14714 11740 14716
rect 11796 14714 11820 14716
rect 11876 14714 11882 14716
rect 11636 14662 11638 14714
rect 11818 14662 11820 14714
rect 11574 14660 11580 14662
rect 11636 14660 11660 14662
rect 11716 14660 11740 14662
rect 11796 14660 11820 14662
rect 11876 14660 11882 14662
rect 11574 14651 11882 14660
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11072 13938 11100 14214
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10796 13326 10824 13806
rect 11256 13326 11284 14350
rect 11992 14074 12020 14776
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 12084 13802 12112 14878
rect 11428 13796 11480 13802
rect 11428 13738 11480 13744
rect 12072 13796 12124 13802
rect 12072 13738 12124 13744
rect 11440 13326 11468 13738
rect 11574 13628 11882 13637
rect 11574 13626 11580 13628
rect 11636 13626 11660 13628
rect 11716 13626 11740 13628
rect 11796 13626 11820 13628
rect 11876 13626 11882 13628
rect 11636 13574 11638 13626
rect 11818 13574 11820 13626
rect 11574 13572 11580 13574
rect 11636 13572 11660 13574
rect 11716 13572 11740 13574
rect 11796 13572 11820 13574
rect 11876 13572 11882 13574
rect 11574 13563 11882 13572
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11428 13320 11480 13326
rect 11612 13320 11664 13326
rect 11428 13262 11480 13268
rect 11518 13288 11574 13297
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10796 12986 10824 13262
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 11256 12646 11284 13262
rect 11440 12918 11468 13262
rect 11574 13268 11612 13274
rect 11574 13262 11664 13268
rect 11574 13246 11652 13262
rect 11796 13252 11848 13258
rect 11518 13223 11574 13232
rect 11796 13194 11848 13200
rect 11808 12986 11836 13194
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11428 12912 11480 12918
rect 11428 12854 11480 12860
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11574 12540 11882 12549
rect 11574 12538 11580 12540
rect 11636 12538 11660 12540
rect 11716 12538 11740 12540
rect 11796 12538 11820 12540
rect 11876 12538 11882 12540
rect 11636 12486 11638 12538
rect 11818 12486 11820 12538
rect 11574 12484 11580 12486
rect 11636 12484 11660 12486
rect 11716 12484 11740 12486
rect 11796 12484 11820 12486
rect 11876 12484 11882 12486
rect 11574 12475 11882 12484
rect 12268 12442 12296 15438
rect 12360 15422 12572 15450
rect 12360 15094 12388 15422
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12452 15094 12480 15302
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12544 14498 12572 15422
rect 12636 14618 12664 15506
rect 12728 15502 12756 16390
rect 12912 16182 12940 18226
rect 13188 17610 13216 18906
rect 13372 18290 13400 20998
rect 13740 20874 13860 20890
rect 13740 20868 13872 20874
rect 13740 20862 13820 20868
rect 13740 19174 13768 20862
rect 13820 20810 13872 20816
rect 13924 20754 13952 22442
rect 13832 20726 13952 20754
rect 13832 19174 13860 20726
rect 13910 20632 13966 20641
rect 14016 20618 14044 23054
rect 13966 20590 14044 20618
rect 13910 20567 13966 20576
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13832 18970 13860 19110
rect 13924 18970 13952 20567
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13912 18352 13964 18358
rect 13912 18294 13964 18300
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 13176 17604 13228 17610
rect 13176 17546 13228 17552
rect 13188 17270 13216 17546
rect 13176 17264 13228 17270
rect 13176 17206 13228 17212
rect 12900 16176 12952 16182
rect 12900 16118 12952 16124
rect 13372 16114 13400 18226
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13832 17338 13860 18158
rect 13924 17882 13952 18294
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13924 17202 13952 17818
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 14016 16658 14044 19790
rect 14108 18306 14136 24822
rect 14200 22094 14228 30194
rect 17420 30122 17448 31925
rect 21284 30326 21312 31925
rect 22198 30492 22506 30501
rect 22198 30490 22204 30492
rect 22260 30490 22284 30492
rect 22340 30490 22364 30492
rect 22420 30490 22444 30492
rect 22500 30490 22506 30492
rect 22260 30438 22262 30490
rect 22442 30438 22444 30490
rect 22198 30436 22204 30438
rect 22260 30436 22284 30438
rect 22340 30436 22364 30438
rect 22420 30436 22444 30438
rect 22500 30436 22506 30438
rect 22198 30427 22506 30436
rect 25424 30326 25452 32014
rect 28998 31925 29054 32725
rect 28906 30696 28962 30705
rect 28906 30631 28962 30640
rect 21272 30320 21324 30326
rect 21272 30262 21324 30268
rect 25412 30320 25464 30326
rect 25412 30262 25464 30268
rect 17592 30252 17644 30258
rect 17592 30194 17644 30200
rect 21916 30252 21968 30258
rect 21916 30194 21968 30200
rect 25320 30252 25372 30258
rect 25320 30194 25372 30200
rect 28724 30252 28776 30258
rect 28724 30194 28776 30200
rect 17408 30116 17460 30122
rect 17408 30058 17460 30064
rect 16212 29708 16264 29714
rect 16212 29650 16264 29656
rect 14280 29572 14332 29578
rect 14280 29514 14332 29520
rect 14292 29238 14320 29514
rect 15115 29404 15423 29413
rect 15115 29402 15121 29404
rect 15177 29402 15201 29404
rect 15257 29402 15281 29404
rect 15337 29402 15361 29404
rect 15417 29402 15423 29404
rect 15177 29350 15179 29402
rect 15359 29350 15361 29402
rect 15115 29348 15121 29350
rect 15177 29348 15201 29350
rect 15257 29348 15281 29350
rect 15337 29348 15361 29350
rect 15417 29348 15423 29350
rect 15115 29339 15423 29348
rect 14280 29232 14332 29238
rect 14280 29174 14332 29180
rect 14292 28150 14320 29174
rect 16224 29170 16252 29650
rect 16488 29572 16540 29578
rect 16488 29514 16540 29520
rect 16500 29306 16528 29514
rect 17132 29504 17184 29510
rect 17132 29446 17184 29452
rect 17316 29504 17368 29510
rect 17316 29446 17368 29452
rect 16488 29300 16540 29306
rect 16488 29242 16540 29248
rect 16672 29232 16724 29238
rect 16672 29174 16724 29180
rect 16212 29164 16264 29170
rect 16212 29106 16264 29112
rect 15568 28960 15620 28966
rect 15568 28902 15620 28908
rect 15936 28960 15988 28966
rect 15936 28902 15988 28908
rect 15580 28558 15608 28902
rect 15948 28626 15976 28902
rect 16224 28762 16252 29106
rect 16580 29096 16632 29102
rect 16580 29038 16632 29044
rect 16212 28756 16264 28762
rect 16212 28698 16264 28704
rect 15936 28620 15988 28626
rect 15936 28562 15988 28568
rect 16592 28558 16620 29038
rect 16684 28762 16712 29174
rect 16672 28756 16724 28762
rect 16672 28698 16724 28704
rect 17144 28626 17172 29446
rect 17328 29306 17356 29446
rect 17316 29300 17368 29306
rect 17316 29242 17368 29248
rect 17132 28620 17184 28626
rect 17132 28562 17184 28568
rect 14464 28552 14516 28558
rect 14464 28494 14516 28500
rect 15568 28552 15620 28558
rect 15568 28494 15620 28500
rect 16488 28552 16540 28558
rect 16488 28494 16540 28500
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 14280 28144 14332 28150
rect 14280 28086 14332 28092
rect 14292 26858 14320 28086
rect 14476 27878 14504 28494
rect 14740 28416 14792 28422
rect 14740 28358 14792 28364
rect 15016 28416 15068 28422
rect 15016 28358 15068 28364
rect 14464 27872 14516 27878
rect 14464 27814 14516 27820
rect 14476 27674 14504 27814
rect 14464 27668 14516 27674
rect 14464 27610 14516 27616
rect 14464 27328 14516 27334
rect 14464 27270 14516 27276
rect 14476 27130 14504 27270
rect 14464 27124 14516 27130
rect 14464 27066 14516 27072
rect 14752 27062 14780 28358
rect 15028 28218 15056 28358
rect 15115 28316 15423 28325
rect 15115 28314 15121 28316
rect 15177 28314 15201 28316
rect 15257 28314 15281 28316
rect 15337 28314 15361 28316
rect 15417 28314 15423 28316
rect 15177 28262 15179 28314
rect 15359 28262 15361 28314
rect 15115 28260 15121 28262
rect 15177 28260 15201 28262
rect 15257 28260 15281 28262
rect 15337 28260 15361 28262
rect 15417 28260 15423 28262
rect 15115 28251 15423 28260
rect 15016 28212 15068 28218
rect 15016 28154 15068 28160
rect 15476 28008 15528 28014
rect 15476 27950 15528 27956
rect 15115 27228 15423 27237
rect 15115 27226 15121 27228
rect 15177 27226 15201 27228
rect 15257 27226 15281 27228
rect 15337 27226 15361 27228
rect 15417 27226 15423 27228
rect 15177 27174 15179 27226
rect 15359 27174 15361 27226
rect 15115 27172 15121 27174
rect 15177 27172 15201 27174
rect 15257 27172 15281 27174
rect 15337 27172 15361 27174
rect 15417 27172 15423 27174
rect 15115 27163 15423 27172
rect 14740 27056 14792 27062
rect 14740 26998 14792 27004
rect 15488 26926 15516 27950
rect 15580 27538 15608 28494
rect 16304 28484 16356 28490
rect 16304 28426 16356 28432
rect 16316 28218 16344 28426
rect 16304 28212 16356 28218
rect 16304 28154 16356 28160
rect 16500 28082 16528 28494
rect 16488 28076 16540 28082
rect 16488 28018 16540 28024
rect 15568 27532 15620 27538
rect 15568 27474 15620 27480
rect 16488 27532 16540 27538
rect 16592 27520 16620 28494
rect 17132 27872 17184 27878
rect 17132 27814 17184 27820
rect 17144 27538 17172 27814
rect 16540 27492 16620 27520
rect 17132 27532 17184 27538
rect 16488 27474 16540 27480
rect 17132 27474 17184 27480
rect 16396 27464 16448 27470
rect 16396 27406 16448 27412
rect 16408 27130 16436 27406
rect 16396 27124 16448 27130
rect 16396 27066 16448 27072
rect 15476 26920 15528 26926
rect 15476 26862 15528 26868
rect 14280 26852 14332 26858
rect 14280 26794 14332 26800
rect 15115 26140 15423 26149
rect 15115 26138 15121 26140
rect 15177 26138 15201 26140
rect 15257 26138 15281 26140
rect 15337 26138 15361 26140
rect 15417 26138 15423 26140
rect 15177 26086 15179 26138
rect 15359 26086 15361 26138
rect 15115 26084 15121 26086
rect 15177 26084 15201 26086
rect 15257 26084 15281 26086
rect 15337 26084 15361 26086
rect 15417 26084 15423 26086
rect 15115 26075 15423 26084
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 14924 25220 14976 25226
rect 14924 25162 14976 25168
rect 14936 24954 14964 25162
rect 14924 24948 14976 24954
rect 14924 24890 14976 24896
rect 14832 24880 14884 24886
rect 14832 24822 14884 24828
rect 14464 24744 14516 24750
rect 14464 24686 14516 24692
rect 14556 24744 14608 24750
rect 14556 24686 14608 24692
rect 14476 24342 14504 24686
rect 14464 24336 14516 24342
rect 14464 24278 14516 24284
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14384 23662 14412 24006
rect 14372 23656 14424 23662
rect 14372 23598 14424 23604
rect 14384 22982 14412 23598
rect 14568 23322 14596 24686
rect 14740 24676 14792 24682
rect 14740 24618 14792 24624
rect 14556 23316 14608 23322
rect 14556 23258 14608 23264
rect 14568 23186 14596 23258
rect 14556 23180 14608 23186
rect 14556 23122 14608 23128
rect 14752 23118 14780 24618
rect 14844 23866 14872 24822
rect 15028 24274 15056 25230
rect 16500 25106 16528 27474
rect 17144 27062 17172 27474
rect 17224 27396 17276 27402
rect 17224 27338 17276 27344
rect 17132 27056 17184 27062
rect 17132 26998 17184 27004
rect 17236 25362 17264 27338
rect 17604 26194 17632 30194
rect 18657 29948 18965 29957
rect 18657 29946 18663 29948
rect 18719 29946 18743 29948
rect 18799 29946 18823 29948
rect 18879 29946 18903 29948
rect 18959 29946 18965 29948
rect 18719 29894 18721 29946
rect 18901 29894 18903 29946
rect 18657 29892 18663 29894
rect 18719 29892 18743 29894
rect 18799 29892 18823 29894
rect 18879 29892 18903 29894
rect 18959 29892 18965 29894
rect 18657 29883 18965 29892
rect 21928 29850 21956 30194
rect 21916 29844 21968 29850
rect 21916 29786 21968 29792
rect 19156 29708 19208 29714
rect 19156 29650 19208 29656
rect 19168 29306 19196 29650
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 25228 29640 25280 29646
rect 25228 29582 25280 29588
rect 19248 29504 19300 29510
rect 19248 29446 19300 29452
rect 20444 29504 20496 29510
rect 20444 29446 20496 29452
rect 19260 29306 19288 29446
rect 19156 29300 19208 29306
rect 19156 29242 19208 29248
rect 19248 29300 19300 29306
rect 19248 29242 19300 29248
rect 20456 29238 20484 29446
rect 20444 29232 20496 29238
rect 20444 29174 20496 29180
rect 20720 29232 20772 29238
rect 20720 29174 20772 29180
rect 18052 29164 18104 29170
rect 18052 29106 18104 29112
rect 18064 28994 18092 29106
rect 18420 29096 18472 29102
rect 18420 29038 18472 29044
rect 20168 29096 20220 29102
rect 20168 29038 20220 29044
rect 18064 28966 18184 28994
rect 18156 28694 18184 28966
rect 18328 28960 18380 28966
rect 18328 28902 18380 28908
rect 18144 28688 18196 28694
rect 18144 28630 18196 28636
rect 17958 28520 18014 28529
rect 17958 28455 18014 28464
rect 17868 28212 17920 28218
rect 17696 28172 17868 28200
rect 17696 28082 17724 28172
rect 17868 28154 17920 28160
rect 17684 28076 17736 28082
rect 17684 28018 17736 28024
rect 17972 27878 18000 28455
rect 18052 28416 18104 28422
rect 18052 28358 18104 28364
rect 18064 28014 18092 28358
rect 18144 28076 18196 28082
rect 18144 28018 18196 28024
rect 18052 28008 18104 28014
rect 18052 27950 18104 27956
rect 17960 27872 18012 27878
rect 17960 27814 18012 27820
rect 18052 27872 18104 27878
rect 18052 27814 18104 27820
rect 18064 26858 18092 27814
rect 18156 27674 18184 28018
rect 18340 28014 18368 28902
rect 18432 28422 18460 29038
rect 18657 28860 18965 28869
rect 18657 28858 18663 28860
rect 18719 28858 18743 28860
rect 18799 28858 18823 28860
rect 18879 28858 18903 28860
rect 18959 28858 18965 28860
rect 18719 28806 18721 28858
rect 18901 28806 18903 28858
rect 18657 28804 18663 28806
rect 18719 28804 18743 28806
rect 18799 28804 18823 28806
rect 18879 28804 18903 28806
rect 18959 28804 18965 28806
rect 18657 28795 18965 28804
rect 19248 28688 19300 28694
rect 19248 28630 19300 28636
rect 19340 28688 19392 28694
rect 19340 28630 19392 28636
rect 18420 28416 18472 28422
rect 18420 28358 18472 28364
rect 18432 28150 18460 28358
rect 19260 28150 19288 28630
rect 18420 28144 18472 28150
rect 18420 28086 18472 28092
rect 19248 28144 19300 28150
rect 19352 28121 19380 28630
rect 20180 28626 20208 29038
rect 20732 28966 20760 29174
rect 20720 28960 20772 28966
rect 20720 28902 20772 28908
rect 20168 28620 20220 28626
rect 20168 28562 20220 28568
rect 19432 28552 19484 28558
rect 19484 28512 19564 28540
rect 19432 28494 19484 28500
rect 19432 28416 19484 28422
rect 19432 28358 19484 28364
rect 19248 28086 19300 28092
rect 19338 28112 19394 28121
rect 18328 28008 18380 28014
rect 18328 27950 18380 27956
rect 18657 27772 18965 27781
rect 18657 27770 18663 27772
rect 18719 27770 18743 27772
rect 18799 27770 18823 27772
rect 18879 27770 18903 27772
rect 18959 27770 18965 27772
rect 18719 27718 18721 27770
rect 18901 27718 18903 27770
rect 18657 27716 18663 27718
rect 18719 27716 18743 27718
rect 18799 27716 18823 27718
rect 18879 27716 18903 27718
rect 18959 27716 18965 27718
rect 18657 27707 18965 27716
rect 18144 27668 18196 27674
rect 18144 27610 18196 27616
rect 18052 26852 18104 26858
rect 18052 26794 18104 26800
rect 18657 26684 18965 26693
rect 18657 26682 18663 26684
rect 18719 26682 18743 26684
rect 18799 26682 18823 26684
rect 18879 26682 18903 26684
rect 18959 26682 18965 26684
rect 18719 26630 18721 26682
rect 18901 26630 18903 26682
rect 18657 26628 18663 26630
rect 18719 26628 18743 26630
rect 18799 26628 18823 26630
rect 18879 26628 18903 26630
rect 18959 26628 18965 26630
rect 18657 26619 18965 26628
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 17604 26166 17724 26194
rect 17224 25356 17276 25362
rect 17224 25298 17276 25304
rect 16580 25220 16632 25226
rect 16580 25162 16632 25168
rect 16592 25106 16620 25162
rect 16408 25078 16620 25106
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 15115 25052 15423 25061
rect 15115 25050 15121 25052
rect 15177 25050 15201 25052
rect 15257 25050 15281 25052
rect 15337 25050 15361 25052
rect 15417 25050 15423 25052
rect 15177 24998 15179 25050
rect 15359 24998 15361 25050
rect 15115 24996 15121 24998
rect 15177 24996 15201 24998
rect 15257 24996 15281 24998
rect 15337 24996 15361 24998
rect 15417 24996 15423 24998
rect 15115 24987 15423 24996
rect 15292 24812 15344 24818
rect 15292 24754 15344 24760
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 15304 24410 15332 24754
rect 15292 24404 15344 24410
rect 15292 24346 15344 24352
rect 15016 24268 15068 24274
rect 15016 24210 15068 24216
rect 15016 24132 15068 24138
rect 15016 24074 15068 24080
rect 14832 23860 14884 23866
rect 14832 23802 14884 23808
rect 15028 23322 15056 24074
rect 15115 23964 15423 23973
rect 15115 23962 15121 23964
rect 15177 23962 15201 23964
rect 15257 23962 15281 23964
rect 15337 23962 15361 23964
rect 15417 23962 15423 23964
rect 15177 23910 15179 23962
rect 15359 23910 15361 23962
rect 15115 23908 15121 23910
rect 15177 23908 15201 23910
rect 15257 23908 15281 23910
rect 15337 23908 15361 23910
rect 15417 23908 15423 23910
rect 15115 23899 15423 23908
rect 15488 23746 15516 24754
rect 15672 24188 15700 24754
rect 15752 24744 15804 24750
rect 16040 24698 16068 24754
rect 15804 24692 16068 24698
rect 15752 24686 16068 24692
rect 15764 24670 16068 24686
rect 16120 24676 16172 24682
rect 15672 24160 15792 24188
rect 15396 23730 15516 23746
rect 15660 23792 15712 23798
rect 15660 23734 15712 23740
rect 15384 23724 15516 23730
rect 15436 23718 15516 23724
rect 15568 23724 15620 23730
rect 15384 23666 15436 23672
rect 15568 23666 15620 23672
rect 15200 23656 15252 23662
rect 15120 23604 15200 23610
rect 15120 23598 15252 23604
rect 15120 23582 15240 23598
rect 15476 23588 15528 23594
rect 14924 23316 14976 23322
rect 14924 23258 14976 23264
rect 15016 23316 15068 23322
rect 15016 23258 15068 23264
rect 14740 23112 14792 23118
rect 14740 23054 14792 23060
rect 14936 22982 14964 23258
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14372 22976 14424 22982
rect 14372 22918 14424 22924
rect 14924 22976 14976 22982
rect 14924 22918 14976 22924
rect 14292 22216 14320 22918
rect 15028 22778 15056 23258
rect 15120 22982 15148 23582
rect 15396 23548 15476 23576
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 15212 23254 15240 23462
rect 15200 23248 15252 23254
rect 15200 23190 15252 23196
rect 15396 23118 15424 23548
rect 15476 23530 15528 23536
rect 15580 23254 15608 23666
rect 15568 23248 15620 23254
rect 15568 23190 15620 23196
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 15476 23044 15528 23050
rect 15476 22986 15528 22992
rect 15568 23044 15620 23050
rect 15568 22986 15620 22992
rect 15108 22976 15160 22982
rect 15108 22918 15160 22924
rect 15115 22876 15423 22885
rect 15115 22874 15121 22876
rect 15177 22874 15201 22876
rect 15257 22874 15281 22876
rect 15337 22874 15361 22876
rect 15417 22874 15423 22876
rect 15177 22822 15179 22874
rect 15359 22822 15361 22874
rect 15115 22820 15121 22822
rect 15177 22820 15201 22822
rect 15257 22820 15281 22822
rect 15337 22820 15361 22822
rect 15417 22820 15423 22822
rect 15115 22811 15423 22820
rect 15016 22772 15068 22778
rect 15016 22714 15068 22720
rect 14832 22432 14884 22438
rect 14832 22374 14884 22380
rect 14844 22234 14872 22374
rect 14832 22228 14884 22234
rect 14292 22188 14688 22216
rect 14200 22066 14412 22094
rect 14280 21004 14332 21010
rect 14280 20946 14332 20952
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14200 20466 14228 20878
rect 14292 20602 14320 20946
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14292 19825 14320 20198
rect 14278 19816 14334 19825
rect 14278 19751 14334 19760
rect 14384 19334 14412 22066
rect 14464 22092 14516 22098
rect 14464 22034 14516 22040
rect 14476 21690 14504 22034
rect 14464 21684 14516 21690
rect 14464 21626 14516 21632
rect 14660 20466 14688 22188
rect 14832 22170 14884 22176
rect 15488 22094 15516 22986
rect 15580 22438 15608 22986
rect 15672 22574 15700 23734
rect 15764 23594 15792 24160
rect 15752 23588 15804 23594
rect 15752 23530 15804 23536
rect 15660 22568 15712 22574
rect 15660 22510 15712 22516
rect 15856 22438 15884 24670
rect 16120 24618 16172 24624
rect 16132 24562 16160 24618
rect 15948 24534 16160 24562
rect 15948 24274 15976 24534
rect 16028 24404 16080 24410
rect 16028 24346 16080 24352
rect 15936 24268 15988 24274
rect 15936 24210 15988 24216
rect 16040 24138 16068 24346
rect 16408 24274 16436 25078
rect 17052 24886 17080 25094
rect 17132 24948 17184 24954
rect 17132 24890 17184 24896
rect 17040 24880 17092 24886
rect 17040 24822 17092 24828
rect 17040 24744 17092 24750
rect 17040 24686 17092 24692
rect 16120 24268 16172 24274
rect 16120 24210 16172 24216
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 15936 24132 15988 24138
rect 15936 24074 15988 24080
rect 16028 24132 16080 24138
rect 16028 24074 16080 24080
rect 15948 23866 15976 24074
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 16040 23798 16068 24074
rect 16028 23792 16080 23798
rect 16028 23734 16080 23740
rect 15936 23588 15988 23594
rect 15936 23530 15988 23536
rect 15948 23254 15976 23530
rect 15936 23248 15988 23254
rect 15936 23190 15988 23196
rect 15948 22506 15976 23190
rect 16040 23186 16068 23734
rect 16132 23730 16160 24210
rect 16304 24200 16356 24206
rect 16304 24142 16356 24148
rect 16212 24132 16264 24138
rect 16212 24074 16264 24080
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 16028 23180 16080 23186
rect 16028 23122 16080 23128
rect 16132 23066 16160 23666
rect 16224 23526 16252 24074
rect 16316 23798 16344 24142
rect 16304 23792 16356 23798
rect 16304 23734 16356 23740
rect 17052 23730 17080 24686
rect 17144 23730 17172 24890
rect 17236 24138 17264 25298
rect 17408 25220 17460 25226
rect 17408 25162 17460 25168
rect 17224 24132 17276 24138
rect 17224 24074 17276 24080
rect 17040 23724 17092 23730
rect 17040 23666 17092 23672
rect 17132 23724 17184 23730
rect 17132 23666 17184 23672
rect 17144 23594 17172 23666
rect 17132 23588 17184 23594
rect 17132 23530 17184 23536
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 16396 23316 16448 23322
rect 16396 23258 16448 23264
rect 16040 23038 16160 23066
rect 15936 22500 15988 22506
rect 15936 22442 15988 22448
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 15488 22066 15608 22094
rect 15115 21788 15423 21797
rect 15115 21786 15121 21788
rect 15177 21786 15201 21788
rect 15257 21786 15281 21788
rect 15337 21786 15361 21788
rect 15417 21786 15423 21788
rect 15177 21734 15179 21786
rect 15359 21734 15361 21786
rect 15115 21732 15121 21734
rect 15177 21732 15201 21734
rect 15257 21732 15281 21734
rect 15337 21732 15361 21734
rect 15417 21732 15423 21734
rect 15115 21723 15423 21732
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14752 21146 14780 21286
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15115 20700 15423 20709
rect 15115 20698 15121 20700
rect 15177 20698 15201 20700
rect 15257 20698 15281 20700
rect 15337 20698 15361 20700
rect 15417 20698 15423 20700
rect 15177 20646 15179 20698
rect 15359 20646 15361 20698
rect 15115 20644 15121 20646
rect 15177 20644 15201 20646
rect 15257 20644 15281 20646
rect 15337 20644 15361 20646
rect 15417 20644 15423 20646
rect 15115 20635 15423 20644
rect 15488 20466 15516 20742
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 14568 19514 14596 20402
rect 14660 20262 14688 20402
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14660 19718 14688 20198
rect 14752 19854 14780 20402
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14924 19780 14976 19786
rect 14924 19722 14976 19728
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14936 19417 14964 19722
rect 15115 19612 15423 19621
rect 15115 19610 15121 19612
rect 15177 19610 15201 19612
rect 15257 19610 15281 19612
rect 15337 19610 15361 19612
rect 15417 19610 15423 19612
rect 15177 19558 15179 19610
rect 15359 19558 15361 19610
rect 15115 19556 15121 19558
rect 15177 19556 15201 19558
rect 15257 19556 15281 19558
rect 15337 19556 15361 19558
rect 15417 19556 15423 19558
rect 15115 19547 15423 19556
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 14922 19408 14978 19417
rect 15212 19394 15240 19450
rect 15120 19378 15240 19394
rect 15580 19378 15608 22066
rect 16040 20942 16068 23038
rect 16212 22976 16264 22982
rect 16212 22918 16264 22924
rect 16028 20936 16080 20942
rect 15948 20913 16028 20924
rect 15934 20904 16028 20913
rect 15990 20896 16028 20904
rect 16028 20878 16080 20884
rect 15934 20839 15990 20848
rect 16120 20868 16172 20874
rect 16120 20810 16172 20816
rect 15844 19780 15896 19786
rect 15844 19722 15896 19728
rect 14922 19343 14978 19352
rect 15108 19372 15240 19378
rect 14384 19306 14504 19334
rect 14372 18692 14424 18698
rect 14372 18634 14424 18640
rect 14384 18426 14412 18634
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14108 18278 14320 18306
rect 14188 17604 14240 17610
rect 14188 17546 14240 17552
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14004 16652 14056 16658
rect 14004 16594 14056 16600
rect 14108 16590 14136 16934
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13188 15994 13216 16050
rect 13084 15972 13136 15978
rect 13188 15966 13308 15994
rect 13084 15914 13136 15920
rect 13096 15570 13124 15914
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13188 15162 13216 15302
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12544 14470 12664 14498
rect 12636 14006 12664 14470
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12624 14000 12676 14006
rect 12346 13968 12402 13977
rect 12624 13942 12676 13948
rect 12346 13903 12402 13912
rect 12360 12850 12388 13903
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 10470 12158 10640 12186
rect 10968 12164 11020 12170
rect 10414 12135 10470 12144
rect 10968 12106 11020 12112
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 10520 10742 10548 11222
rect 10980 11150 11008 12106
rect 12084 11762 12112 12242
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 11164 10742 11192 11494
rect 11574 11452 11882 11461
rect 11574 11450 11580 11452
rect 11636 11450 11660 11452
rect 11716 11450 11740 11452
rect 11796 11450 11820 11452
rect 11876 11450 11882 11452
rect 11636 11398 11638 11450
rect 11818 11398 11820 11450
rect 11574 11396 11580 11398
rect 11636 11396 11660 11398
rect 11716 11396 11740 11398
rect 11796 11396 11820 11398
rect 11876 11396 11882 11398
rect 11574 11387 11882 11396
rect 10508 10736 10560 10742
rect 10508 10678 10560 10684
rect 11152 10736 11204 10742
rect 11152 10678 11204 10684
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10244 9654 10272 10066
rect 10336 10062 10364 10610
rect 10520 10606 10548 10678
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10336 9761 10364 9998
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10322 9752 10378 9761
rect 10322 9687 10378 9696
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10232 9444 10284 9450
rect 10232 9386 10284 9392
rect 10244 9110 10272 9386
rect 10336 9353 10364 9687
rect 10428 9518 10456 9862
rect 10520 9722 10548 10406
rect 10612 9722 10640 10474
rect 10968 10192 11020 10198
rect 10968 10134 11020 10140
rect 10980 10062 11008 10134
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10704 9654 10732 9862
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10416 9512 10468 9518
rect 10692 9512 10744 9518
rect 10468 9460 10692 9466
rect 10416 9454 10744 9460
rect 10428 9438 10732 9454
rect 10508 9376 10560 9382
rect 10322 9344 10378 9353
rect 10508 9318 10560 9324
rect 10322 9279 10378 9288
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9968 8634 9996 8774
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 10152 6798 10180 8978
rect 10520 8498 10548 9318
rect 10796 9042 10824 9998
rect 10874 9752 10930 9761
rect 10930 9722 11008 9738
rect 10930 9716 11020 9722
rect 10930 9710 10968 9716
rect 10874 9687 10930 9696
rect 10968 9658 11020 9664
rect 11072 9518 11100 9998
rect 11164 9926 11192 10678
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11440 10062 11468 10542
rect 11574 10364 11882 10373
rect 11574 10362 11580 10364
rect 11636 10362 11660 10364
rect 11716 10362 11740 10364
rect 11796 10362 11820 10364
rect 11876 10362 11882 10364
rect 11636 10310 11638 10362
rect 11818 10310 11820 10362
rect 11574 10308 11580 10310
rect 11636 10308 11660 10310
rect 11716 10308 11740 10310
rect 11796 10308 11820 10310
rect 11876 10308 11882 10310
rect 11574 10299 11882 10308
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11150 9752 11206 9761
rect 11256 9738 11284 9998
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11206 9710 11284 9738
rect 11150 9687 11206 9696
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10506 8256 10562 8265
rect 10506 8191 10562 8200
rect 10520 7410 10548 8191
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10520 7002 10548 7346
rect 11164 7342 11192 8978
rect 11348 8906 11376 9590
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11336 8900 11388 8906
rect 11256 8860 11336 8888
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9634 5908 9686 5914
rect 9508 5868 9634 5896
rect 9508 5710 9536 5868
rect 9634 5850 9686 5856
rect 9968 5794 9996 6258
rect 10060 5914 10088 6734
rect 10152 6322 10180 6734
rect 10244 6458 10272 6734
rect 10416 6724 10468 6730
rect 10416 6666 10468 6672
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9968 5766 10088 5794
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 7104 5296 7156 5302
rect 7104 5238 7156 5244
rect 8956 4690 8984 5306
rect 9324 4690 9352 5510
rect 9784 5234 9812 5510
rect 9876 5250 9904 5510
rect 9876 5234 9996 5250
rect 9772 5228 9824 5234
rect 9876 5228 10008 5234
rect 9876 5222 9956 5228
rect 9772 5170 9824 5176
rect 9956 5170 10008 5176
rect 10060 5166 10088 5766
rect 10152 5710 10180 6258
rect 10428 6254 10456 6666
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10520 5760 10548 6326
rect 10612 6322 10640 6938
rect 11164 6882 11192 7278
rect 11256 7002 11284 8860
rect 11336 8842 11388 8848
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11348 7002 11376 7346
rect 11440 7206 11468 9318
rect 11574 9276 11882 9285
rect 11574 9274 11580 9276
rect 11636 9274 11660 9276
rect 11716 9274 11740 9276
rect 11796 9274 11820 9276
rect 11876 9274 11882 9276
rect 11636 9222 11638 9274
rect 11818 9222 11820 9274
rect 11574 9220 11580 9222
rect 11636 9220 11660 9222
rect 11716 9220 11740 9222
rect 11796 9220 11820 9222
rect 11876 9220 11882 9222
rect 11574 9211 11882 9220
rect 11992 9042 12020 9862
rect 12268 9625 12296 12378
rect 12544 12170 12572 13398
rect 12636 12850 12664 13942
rect 13004 13870 13032 14350
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12820 12434 12848 12582
rect 12728 12406 12848 12434
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12728 11898 12756 12406
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 13004 11694 13032 13806
rect 13280 13530 13308 15966
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13280 12986 13308 13466
rect 13372 13394 13400 16050
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13464 14482 13492 14962
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 13266 11112 13322 11121
rect 13648 11082 13676 15982
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13832 14006 13860 15846
rect 13924 15502 13952 16050
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13924 15162 13952 15438
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 14096 13796 14148 13802
rect 14096 13738 14148 13744
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13740 11762 13768 12106
rect 13832 11898 13860 12786
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13924 12238 13952 12582
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13266 11047 13322 11056
rect 13636 11076 13688 11082
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10606 12480 10950
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12254 9616 12310 9625
rect 12360 9586 12388 10202
rect 13280 10062 13308 11047
rect 13636 11018 13688 11024
rect 13648 10674 13676 11018
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13556 10266 13584 10406
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13360 9988 13412 9994
rect 13360 9930 13412 9936
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12254 9551 12310 9560
rect 12348 9580 12400 9586
rect 11980 9036 12032 9042
rect 12032 8996 12204 9024
rect 11980 8978 12032 8984
rect 11574 8188 11882 8197
rect 11574 8186 11580 8188
rect 11636 8186 11660 8188
rect 11716 8186 11740 8188
rect 11796 8186 11820 8188
rect 11876 8186 11882 8188
rect 11636 8134 11638 8186
rect 11818 8134 11820 8186
rect 11574 8132 11580 8134
rect 11636 8132 11660 8134
rect 11716 8132 11740 8134
rect 11796 8132 11820 8134
rect 11876 8132 11882 8134
rect 11574 8123 11882 8132
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 10888 6854 11192 6882
rect 11440 6866 11468 7142
rect 11574 7100 11882 7109
rect 11574 7098 11580 7100
rect 11636 7098 11660 7100
rect 11716 7098 11740 7100
rect 11796 7098 11820 7100
rect 11876 7098 11882 7100
rect 11636 7046 11638 7098
rect 11818 7046 11820 7098
rect 11574 7044 11580 7046
rect 11636 7044 11660 7046
rect 11716 7044 11740 7046
rect 11796 7044 11820 7046
rect 11876 7044 11882 7046
rect 11574 7035 11882 7044
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11428 6860 11480 6866
rect 10782 6760 10838 6769
rect 10782 6695 10838 6704
rect 10796 6662 10824 6695
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10428 5732 10548 5760
rect 10140 5704 10192 5710
rect 10428 5658 10456 5732
rect 10140 5646 10192 5652
rect 10152 5234 10180 5646
rect 10336 5642 10456 5658
rect 10888 5642 10916 6854
rect 11428 6802 11480 6808
rect 10968 6792 11020 6798
rect 11020 6740 11100 6746
rect 10968 6734 11100 6740
rect 10980 6718 11100 6734
rect 11532 6730 11560 6938
rect 11992 6882 12020 7142
rect 12084 7002 12112 7346
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11796 6860 11848 6866
rect 11992 6854 12112 6882
rect 11796 6802 11848 6808
rect 10966 6624 11022 6633
rect 10966 6559 11022 6568
rect 10980 6322 11008 6559
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 11072 5914 11100 6718
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11164 6322 11192 6598
rect 11152 6316 11204 6322
rect 11204 6276 11284 6304
rect 11152 6258 11204 6264
rect 11152 6180 11204 6186
rect 11152 6122 11204 6128
rect 11164 5914 11192 6122
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 10324 5636 10456 5642
rect 10376 5630 10456 5636
rect 10876 5636 10928 5642
rect 10324 5578 10376 5584
rect 10876 5578 10928 5584
rect 10888 5234 10916 5578
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10152 4826 10180 5170
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10336 4690 10364 4966
rect 11072 4826 11100 5850
rect 11164 5710 11192 5850
rect 11256 5710 11284 6276
rect 11348 5914 11376 6666
rect 11716 6458 11744 6802
rect 11808 6458 11836 6802
rect 12084 6798 12112 6854
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11440 5778 11468 6394
rect 11574 6012 11882 6021
rect 11574 6010 11580 6012
rect 11636 6010 11660 6012
rect 11716 6010 11740 6012
rect 11796 6010 11820 6012
rect 11876 6010 11882 6012
rect 11636 5958 11638 6010
rect 11818 5958 11820 6010
rect 11574 5956 11580 5958
rect 11636 5956 11660 5958
rect 11716 5956 11740 5958
rect 11796 5956 11820 5958
rect 11876 5956 11882 5958
rect 11574 5947 11882 5956
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11428 5636 11480 5642
rect 11428 5578 11480 5584
rect 11348 5166 11376 5578
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 11348 4622 11376 5102
rect 11440 4826 11468 5578
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11808 5234 11836 5510
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 12084 5166 12112 6734
rect 12176 6662 12204 8996
rect 12268 8974 12296 9551
rect 12348 9522 12400 9528
rect 13096 9178 13124 9862
rect 13176 9648 13228 9654
rect 13174 9616 13176 9625
rect 13228 9616 13230 9625
rect 13174 9551 13230 9560
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13280 8634 13308 8842
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13372 8430 13400 9930
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 13464 8430 13492 9590
rect 13740 9382 13768 11698
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13924 10062 13952 10202
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13832 9654 13860 9862
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13648 8566 13676 8774
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12728 7478 12756 8298
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12820 7546 12848 7890
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 13372 7410 13400 7686
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13464 7392 13492 8366
rect 13740 7818 13768 8910
rect 13912 8900 13964 8906
rect 13912 8842 13964 8848
rect 13924 8294 13952 8842
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13544 7404 13596 7410
rect 13464 7364 13544 7392
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 13464 6254 13492 7364
rect 13544 7346 13596 7352
rect 13648 7002 13676 7754
rect 13924 7750 13952 8230
rect 14016 8090 14044 12718
rect 14108 12209 14136 13738
rect 14094 12200 14150 12209
rect 14094 12135 14150 12144
rect 14108 11762 14136 12135
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14108 10606 14136 10746
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14108 9518 14136 10542
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14108 8430 14136 9454
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 14016 7886 14044 8026
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13924 6934 13952 7686
rect 14016 7206 14044 7822
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14108 7018 14136 8366
rect 14200 8022 14228 17546
rect 14292 14414 14320 18278
rect 14372 16720 14424 16726
rect 14372 16662 14424 16668
rect 14384 16522 14412 16662
rect 14372 16516 14424 16522
rect 14372 16458 14424 16464
rect 14476 16402 14504 19306
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14568 16726 14596 18634
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14752 18154 14780 18566
rect 14740 18148 14792 18154
rect 14740 18090 14792 18096
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14660 16794 14688 17478
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14556 16720 14608 16726
rect 14556 16662 14608 16668
rect 14936 16674 14964 19343
rect 15160 19366 15240 19372
rect 15292 19372 15344 19378
rect 15108 19314 15160 19320
rect 15292 19314 15344 19320
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 15304 19258 15332 19314
rect 15856 19292 15884 19722
rect 16132 19514 16160 20810
rect 16120 19508 16172 19514
rect 16120 19450 16172 19456
rect 15936 19304 15988 19310
rect 15856 19264 15936 19292
rect 15304 19230 15608 19258
rect 15936 19246 15988 19252
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15028 18034 15056 19110
rect 15488 18902 15516 19110
rect 15580 18902 15608 19230
rect 15948 18970 15976 19246
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 15115 18524 15423 18533
rect 15115 18522 15121 18524
rect 15177 18522 15201 18524
rect 15257 18522 15281 18524
rect 15337 18522 15361 18524
rect 15417 18522 15423 18524
rect 15177 18470 15179 18522
rect 15359 18470 15361 18522
rect 15115 18468 15121 18470
rect 15177 18468 15201 18470
rect 15257 18468 15281 18470
rect 15337 18468 15361 18470
rect 15417 18468 15423 18470
rect 15115 18459 15423 18468
rect 15488 18358 15516 18634
rect 16132 18630 16160 19450
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 15476 18352 15528 18358
rect 15528 18312 15608 18340
rect 15476 18294 15528 18300
rect 15580 18222 15608 18312
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15568 18216 15620 18222
rect 16132 18170 16160 18566
rect 15568 18158 15620 18164
rect 15028 18006 15240 18034
rect 15212 17921 15240 18006
rect 15198 17912 15254 17921
rect 15198 17847 15254 17856
rect 15115 17436 15423 17445
rect 15115 17434 15121 17436
rect 15177 17434 15201 17436
rect 15257 17434 15281 17436
rect 15337 17434 15361 17436
rect 15417 17434 15423 17436
rect 15177 17382 15179 17434
rect 15359 17382 15361 17434
rect 15115 17380 15121 17382
rect 15177 17380 15201 17382
rect 15257 17380 15281 17382
rect 15337 17380 15361 17382
rect 15417 17380 15423 17382
rect 15115 17371 15423 17380
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15120 16794 15148 17138
rect 15488 17134 15516 18158
rect 16040 18142 16160 18170
rect 16040 17270 16068 18142
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 16132 17678 16160 18022
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 16132 17270 16160 17614
rect 16028 17264 16080 17270
rect 16028 17206 16080 17212
rect 16120 17264 16172 17270
rect 16120 17206 16172 17212
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15108 16788 15160 16794
rect 15108 16730 15160 16736
rect 14936 16646 15056 16674
rect 15028 16590 15056 16646
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 14476 16374 14596 16402
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14384 14958 14412 15438
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14476 12850 14504 13194
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14384 12646 14412 12786
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14278 12336 14334 12345
rect 14278 12271 14334 12280
rect 14292 11830 14320 12271
rect 14280 11824 14332 11830
rect 14280 11766 14332 11772
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14292 10674 14320 11494
rect 14372 11076 14424 11082
rect 14372 11018 14424 11024
rect 14384 10674 14412 11018
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14384 9926 14412 10610
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14292 9382 14320 9590
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14292 8566 14320 9318
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 14188 8016 14240 8022
rect 14188 7958 14240 7964
rect 14292 7478 14320 8502
rect 14476 7970 14504 10406
rect 14384 7942 14504 7970
rect 14384 7886 14412 7942
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14280 7472 14332 7478
rect 14016 6990 14136 7018
rect 14200 7420 14280 7426
rect 14200 7414 14332 7420
rect 14200 7398 14320 7414
rect 13912 6928 13964 6934
rect 13912 6870 13964 6876
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13924 6633 13952 6734
rect 13910 6624 13966 6633
rect 13910 6559 13966 6568
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 13452 6248 13504 6254
rect 13452 6190 13504 6196
rect 12452 5522 12480 6190
rect 14016 5846 14044 6990
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14108 6769 14136 6802
rect 14094 6760 14150 6769
rect 14094 6695 14150 6704
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 6458 14136 6598
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14200 6390 14228 7398
rect 14476 7002 14504 7686
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14188 6384 14240 6390
rect 14188 6326 14240 6332
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 12360 5494 12480 5522
rect 12360 5370 12388 5494
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12452 5166 12480 5306
rect 14200 5234 14228 6326
rect 14568 5370 14596 16374
rect 14660 14414 14688 16526
rect 14924 16516 14976 16522
rect 14924 16458 14976 16464
rect 14832 16448 14884 16454
rect 14832 16390 14884 16396
rect 14844 16114 14872 16390
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14660 13938 14688 14350
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14660 12986 14688 13330
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14752 12782 14780 14758
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14844 13938 14872 14214
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14660 12238 14688 12718
rect 14936 12238 14964 16458
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 15028 16046 15056 16390
rect 15115 16348 15423 16357
rect 15115 16346 15121 16348
rect 15177 16346 15201 16348
rect 15257 16346 15281 16348
rect 15337 16346 15361 16348
rect 15417 16346 15423 16348
rect 15177 16294 15179 16346
rect 15359 16294 15361 16346
rect 15115 16292 15121 16294
rect 15177 16292 15201 16294
rect 15257 16292 15281 16294
rect 15337 16292 15361 16294
rect 15417 16292 15423 16294
rect 15115 16283 15423 16292
rect 15488 16114 15608 16130
rect 15476 16108 15608 16114
rect 15528 16102 15608 16108
rect 15476 16050 15528 16056
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15115 15260 15423 15269
rect 15115 15258 15121 15260
rect 15177 15258 15201 15260
rect 15257 15258 15281 15260
rect 15337 15258 15361 15260
rect 15417 15258 15423 15260
rect 15177 15206 15179 15258
rect 15359 15206 15361 15258
rect 15115 15204 15121 15206
rect 15177 15204 15201 15206
rect 15257 15204 15281 15206
rect 15337 15204 15361 15206
rect 15417 15204 15423 15206
rect 15115 15195 15423 15204
rect 15488 15076 15516 15846
rect 15396 15048 15516 15076
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 15120 14618 15148 14758
rect 15396 14618 15424 15048
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15120 14362 15148 14554
rect 15028 14334 15148 14362
rect 15028 13938 15056 14334
rect 15115 14172 15423 14181
rect 15115 14170 15121 14172
rect 15177 14170 15201 14172
rect 15257 14170 15281 14172
rect 15337 14170 15361 14172
rect 15417 14170 15423 14172
rect 15177 14118 15179 14170
rect 15359 14118 15361 14170
rect 15115 14116 15121 14118
rect 15177 14116 15201 14118
rect 15257 14116 15281 14118
rect 15337 14116 15361 14118
rect 15417 14116 15423 14118
rect 15115 14107 15423 14116
rect 15384 14000 15436 14006
rect 15384 13942 15436 13948
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 15396 13682 15424 13942
rect 15488 13802 15516 14894
rect 15476 13796 15528 13802
rect 15476 13738 15528 13744
rect 15396 13654 15516 13682
rect 15115 13084 15423 13093
rect 15115 13082 15121 13084
rect 15177 13082 15201 13084
rect 15257 13082 15281 13084
rect 15337 13082 15361 13084
rect 15417 13082 15423 13084
rect 15177 13030 15179 13082
rect 15359 13030 15361 13082
rect 15115 13028 15121 13030
rect 15177 13028 15201 13030
rect 15257 13028 15281 13030
rect 15337 13028 15361 13030
rect 15417 13028 15423 13030
rect 15115 13019 15423 13028
rect 15108 12368 15160 12374
rect 15292 12368 15344 12374
rect 15160 12328 15292 12356
rect 15108 12310 15160 12316
rect 15292 12310 15344 12316
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 15115 11996 15423 12005
rect 15115 11994 15121 11996
rect 15177 11994 15201 11996
rect 15257 11994 15281 11996
rect 15337 11994 15361 11996
rect 15417 11994 15423 11996
rect 15177 11942 15179 11994
rect 15359 11942 15361 11994
rect 15115 11940 15121 11942
rect 15177 11940 15201 11942
rect 15257 11940 15281 11942
rect 15337 11940 15361 11942
rect 15417 11940 15423 11942
rect 15115 11931 15423 11940
rect 15488 11762 15516 13654
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 14660 7886 14688 11698
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14752 10810 14780 11494
rect 15115 10908 15423 10917
rect 15115 10906 15121 10908
rect 15177 10906 15201 10908
rect 15257 10906 15281 10908
rect 15337 10906 15361 10908
rect 15417 10906 15423 10908
rect 15177 10854 15179 10906
rect 15359 10854 15361 10906
rect 15115 10852 15121 10854
rect 15177 10852 15201 10854
rect 15257 10852 15281 10854
rect 15337 10852 15361 10854
rect 15417 10852 15423 10854
rect 15115 10843 15423 10852
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 15580 10690 15608 16102
rect 15672 15162 15700 16526
rect 15752 16516 15804 16522
rect 15752 16458 15804 16464
rect 15764 15910 15792 16458
rect 15856 16114 15884 17138
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15764 15094 15792 15438
rect 15856 15314 15884 16050
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 15948 15434 15976 15846
rect 16132 15706 16160 15846
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 15936 15428 15988 15434
rect 15936 15370 15988 15376
rect 15856 15286 15976 15314
rect 15752 15088 15804 15094
rect 15752 15030 15804 15036
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15672 14260 15700 14554
rect 15752 14408 15804 14414
rect 15804 14368 15884 14396
rect 15752 14350 15804 14356
rect 15672 14232 15792 14260
rect 15764 13462 15792 14232
rect 15752 13456 15804 13462
rect 15752 13398 15804 13404
rect 15764 12374 15792 13398
rect 15752 12368 15804 12374
rect 15752 12310 15804 12316
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15396 10662 15608 10690
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 15304 9994 15332 10474
rect 15396 10062 15424 10662
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15672 10062 15700 10406
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15115 9820 15423 9829
rect 15115 9818 15121 9820
rect 15177 9818 15201 9820
rect 15257 9818 15281 9820
rect 15337 9818 15361 9820
rect 15417 9818 15423 9820
rect 15177 9766 15179 9818
rect 15359 9766 15361 9818
rect 15115 9764 15121 9766
rect 15177 9764 15201 9766
rect 15257 9764 15281 9766
rect 15337 9764 15361 9766
rect 15417 9764 15423 9766
rect 15115 9755 15423 9764
rect 15115 8732 15423 8741
rect 15115 8730 15121 8732
rect 15177 8730 15201 8732
rect 15257 8730 15281 8732
rect 15337 8730 15361 8732
rect 15417 8730 15423 8732
rect 15177 8678 15179 8730
rect 15359 8678 15361 8730
rect 15115 8676 15121 8678
rect 15177 8676 15201 8678
rect 15257 8676 15281 8678
rect 15337 8676 15361 8678
rect 15417 8676 15423 8678
rect 15115 8667 15423 8676
rect 14648 7880 14700 7886
rect 15016 7880 15068 7886
rect 14700 7840 14780 7868
rect 14648 7822 14700 7828
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14660 7546 14688 7686
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 14752 6730 14780 7840
rect 15016 7822 15068 7828
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15028 7342 15056 7822
rect 15115 7644 15423 7653
rect 15115 7642 15121 7644
rect 15177 7642 15201 7644
rect 15257 7642 15281 7644
rect 15337 7642 15361 7644
rect 15417 7642 15423 7644
rect 15177 7590 15179 7642
rect 15359 7590 15361 7642
rect 15115 7588 15121 7590
rect 15177 7588 15201 7590
rect 15257 7588 15281 7590
rect 15337 7588 15361 7590
rect 15417 7588 15423 7590
rect 15115 7579 15423 7588
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15488 6866 15516 7822
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 14740 6724 14792 6730
rect 14740 6666 14792 6672
rect 15115 6556 15423 6565
rect 15115 6554 15121 6556
rect 15177 6554 15201 6556
rect 15257 6554 15281 6556
rect 15337 6554 15361 6556
rect 15417 6554 15423 6556
rect 15177 6502 15179 6554
rect 15359 6502 15361 6554
rect 15115 6500 15121 6502
rect 15177 6500 15201 6502
rect 15257 6500 15281 6502
rect 15337 6500 15361 6502
rect 15417 6500 15423 6502
rect 15115 6491 15423 6500
rect 15488 6390 15516 6802
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15115 5468 15423 5477
rect 15115 5466 15121 5468
rect 15177 5466 15201 5468
rect 15257 5466 15281 5468
rect 15337 5466 15361 5468
rect 15417 5466 15423 5468
rect 15177 5414 15179 5466
rect 15359 5414 15361 5466
rect 15115 5412 15121 5414
rect 15177 5412 15201 5414
rect 15257 5412 15281 5414
rect 15337 5412 15361 5414
rect 15417 5412 15423 5414
rect 15115 5403 15423 5412
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 11574 4924 11882 4933
rect 11574 4922 11580 4924
rect 11636 4922 11660 4924
rect 11716 4922 11740 4924
rect 11796 4922 11820 4924
rect 11876 4922 11882 4924
rect 11636 4870 11638 4922
rect 11818 4870 11820 4922
rect 11574 4868 11580 4870
rect 11636 4868 11660 4870
rect 11716 4868 11740 4870
rect 11796 4868 11820 4870
rect 11876 4868 11882 4870
rect 11574 4859 11882 4868
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 8032 4380 8340 4389
rect 8032 4378 8038 4380
rect 8094 4378 8118 4380
rect 8174 4378 8198 4380
rect 8254 4378 8278 4380
rect 8334 4378 8340 4380
rect 8094 4326 8096 4378
rect 8276 4326 8278 4378
rect 8032 4324 8038 4326
rect 8094 4324 8118 4326
rect 8174 4324 8198 4326
rect 8254 4324 8278 4326
rect 8334 4324 8340 4326
rect 8032 4315 8340 4324
rect 13004 4146 13032 4558
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 2410 3975 2466 3984
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2240 3738 2268 3878
rect 4491 3836 4799 3845
rect 4491 3834 4497 3836
rect 4553 3834 4577 3836
rect 4633 3834 4657 3836
rect 4713 3834 4737 3836
rect 4793 3834 4799 3836
rect 4553 3782 4555 3834
rect 4735 3782 4737 3834
rect 4491 3780 4497 3782
rect 4553 3780 4577 3782
rect 4633 3780 4657 3782
rect 4713 3780 4737 3782
rect 4793 3780 4799 3782
rect 4491 3771 4799 3780
rect 11574 3836 11882 3845
rect 11574 3834 11580 3836
rect 11636 3834 11660 3836
rect 11716 3834 11740 3836
rect 11796 3834 11820 3836
rect 11876 3834 11882 3836
rect 11636 3782 11638 3834
rect 11818 3782 11820 3834
rect 11574 3780 11580 3782
rect 11636 3780 11660 3782
rect 11716 3780 11740 3782
rect 11796 3780 11820 3782
rect 11876 3780 11882 3782
rect 11574 3771 11882 3780
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 12900 3528 12952 3534
rect 938 3496 994 3505
rect 12900 3470 12952 3476
rect 938 3431 994 3440
rect 952 3398 980 3431
rect 12912 3398 12940 3470
rect 940 3392 992 3398
rect 940 3334 992 3340
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 2240 2446 2268 3334
rect 8032 3292 8340 3301
rect 8032 3290 8038 3292
rect 8094 3290 8118 3292
rect 8174 3290 8198 3292
rect 8254 3290 8278 3292
rect 8334 3290 8340 3292
rect 8094 3238 8096 3290
rect 8276 3238 8278 3290
rect 8032 3236 8038 3238
rect 8094 3236 8118 3238
rect 8174 3236 8198 3238
rect 8254 3236 8278 3238
rect 8334 3236 8340 3238
rect 8032 3227 8340 3236
rect 4491 2748 4799 2757
rect 4491 2746 4497 2748
rect 4553 2746 4577 2748
rect 4633 2746 4657 2748
rect 4713 2746 4737 2748
rect 4793 2746 4799 2748
rect 4553 2694 4555 2746
rect 4735 2694 4737 2746
rect 4491 2692 4497 2694
rect 4553 2692 4577 2694
rect 4633 2692 4657 2694
rect 4713 2692 4737 2694
rect 4793 2692 4799 2694
rect 4491 2683 4799 2692
rect 11574 2748 11882 2757
rect 11574 2746 11580 2748
rect 11636 2746 11660 2748
rect 11716 2746 11740 2748
rect 11796 2746 11820 2748
rect 11876 2746 11882 2748
rect 11636 2694 11638 2746
rect 11818 2694 11820 2746
rect 11574 2692 11580 2694
rect 11636 2692 11660 2694
rect 11716 2692 11740 2694
rect 11796 2692 11820 2694
rect 11876 2692 11882 2694
rect 11574 2683 11882 2692
rect 12820 2650 12848 3334
rect 13004 3194 13032 4082
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 13096 3194 13124 3878
rect 13188 3738 13216 4218
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13174 3496 13230 3505
rect 13174 3431 13176 3440
rect 13228 3431 13230 3440
rect 13176 3402 13228 3408
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 13188 2446 13216 2790
rect 13280 2650 13308 4558
rect 14004 4548 14056 4554
rect 14004 4490 14056 4496
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 13372 3534 13400 3946
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 13464 3534 13492 3878
rect 13544 3664 13596 3670
rect 13924 3652 13952 3878
rect 14016 3670 14044 4490
rect 15115 4380 15423 4389
rect 15115 4378 15121 4380
rect 15177 4378 15201 4380
rect 15257 4378 15281 4380
rect 15337 4378 15361 4380
rect 15417 4378 15423 4380
rect 15177 4326 15179 4378
rect 15359 4326 15361 4378
rect 15115 4324 15121 4326
rect 15177 4324 15201 4326
rect 15257 4324 15281 4326
rect 15337 4324 15361 4326
rect 15417 4324 15423 4326
rect 15115 4315 15423 4324
rect 15580 4282 15608 9862
rect 15764 9042 15792 11698
rect 15856 11694 15884 14368
rect 15948 13870 15976 15286
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 16132 12850 16160 15438
rect 16224 15162 16252 22918
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16316 20777 16344 21830
rect 16302 20768 16358 20777
rect 16302 20703 16358 20712
rect 16408 17542 16436 23258
rect 16764 23044 16816 23050
rect 16764 22986 16816 22992
rect 16488 22568 16540 22574
rect 16488 22510 16540 22516
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16500 22098 16528 22510
rect 16488 22094 16540 22098
rect 16488 22092 16620 22094
rect 16540 22066 16620 22092
rect 16488 22034 16540 22040
rect 16592 21486 16620 22066
rect 16684 21894 16712 22510
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 16592 20942 16620 21422
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16500 20466 16528 20878
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 16500 18766 16528 20402
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16316 15706 16344 15846
rect 16304 15700 16356 15706
rect 16304 15642 16356 15648
rect 16302 15192 16358 15201
rect 16212 15156 16264 15162
rect 16302 15127 16358 15136
rect 16212 15098 16264 15104
rect 16224 14618 16252 15098
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16316 14482 16344 15127
rect 16408 15094 16436 17478
rect 16500 16998 16528 18702
rect 16592 18426 16620 20878
rect 16776 18766 16804 22986
rect 17236 22030 17264 24074
rect 17420 23322 17448 25162
rect 17500 23792 17552 23798
rect 17500 23734 17552 23740
rect 17408 23316 17460 23322
rect 17408 23258 17460 23264
rect 17512 22964 17540 23734
rect 17592 22976 17644 22982
rect 17512 22936 17592 22964
rect 17592 22918 17644 22924
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 17236 21622 17264 21966
rect 17224 21616 17276 21622
rect 17224 21558 17276 21564
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 16960 21146 16988 21422
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 17132 20868 17184 20874
rect 17132 20810 17184 20816
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 16856 20460 16908 20466
rect 16856 20402 16908 20408
rect 16868 20058 16896 20402
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16960 19961 16988 20538
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 17052 20058 17080 20402
rect 17144 20262 17172 20810
rect 17604 20466 17632 22918
rect 17696 22001 17724 26166
rect 17868 25832 17920 25838
rect 17868 25774 17920 25780
rect 17880 25294 17908 25774
rect 17868 25288 17920 25294
rect 17868 25230 17920 25236
rect 17972 24818 18000 26318
rect 19260 26194 19288 28086
rect 19338 28047 19394 28056
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 19352 27674 19380 27950
rect 19340 27668 19392 27674
rect 19340 27610 19392 27616
rect 19444 27470 19472 28358
rect 19536 27470 19564 28512
rect 19892 27872 19944 27878
rect 19892 27814 19944 27820
rect 19904 27470 19932 27814
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19524 27464 19576 27470
rect 19524 27406 19576 27412
rect 19892 27464 19944 27470
rect 19892 27406 19944 27412
rect 19536 27130 19564 27406
rect 20076 27396 20128 27402
rect 20180 27384 20208 28562
rect 20260 28416 20312 28422
rect 20260 28358 20312 28364
rect 20272 27946 20300 28358
rect 20260 27940 20312 27946
rect 20260 27882 20312 27888
rect 20272 27402 20300 27882
rect 20732 27402 20760 28902
rect 20824 28762 20852 29582
rect 22198 29404 22506 29413
rect 22198 29402 22204 29404
rect 22260 29402 22284 29404
rect 22340 29402 22364 29404
rect 22420 29402 22444 29404
rect 22500 29402 22506 29404
rect 22260 29350 22262 29402
rect 22442 29350 22444 29402
rect 22198 29348 22204 29350
rect 22260 29348 22284 29350
rect 22340 29348 22364 29350
rect 22420 29348 22444 29350
rect 22500 29348 22506 29350
rect 22198 29339 22506 29348
rect 22836 29164 22888 29170
rect 22836 29106 22888 29112
rect 22100 29096 22152 29102
rect 22100 29038 22152 29044
rect 21364 28960 21416 28966
rect 21364 28902 21416 28908
rect 20812 28756 20864 28762
rect 20812 28698 20864 28704
rect 21272 28756 21324 28762
rect 21272 28698 21324 28704
rect 20812 28552 20864 28558
rect 20864 28512 20944 28540
rect 20812 28494 20864 28500
rect 20812 28076 20864 28082
rect 20812 28018 20864 28024
rect 20824 27538 20852 28018
rect 20812 27532 20864 27538
rect 20812 27474 20864 27480
rect 20128 27356 20208 27384
rect 20260 27396 20312 27402
rect 20076 27338 20128 27344
rect 20260 27338 20312 27344
rect 20720 27396 20772 27402
rect 20720 27338 20772 27344
rect 19524 27124 19576 27130
rect 19524 27066 19576 27072
rect 19432 26308 19484 26314
rect 19432 26250 19484 26256
rect 19800 26308 19852 26314
rect 19800 26250 19852 26256
rect 19260 26166 19380 26194
rect 19352 25974 19380 26166
rect 18236 25968 18288 25974
rect 18236 25910 18288 25916
rect 19340 25968 19392 25974
rect 19340 25910 19392 25916
rect 18144 25424 18196 25430
rect 18144 25366 18196 25372
rect 18156 24818 18184 25366
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 17960 24200 18012 24206
rect 17960 24142 18012 24148
rect 17972 23662 18000 24142
rect 18052 24132 18104 24138
rect 18052 24074 18104 24080
rect 18064 23662 18092 24074
rect 17960 23656 18012 23662
rect 17960 23598 18012 23604
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 18064 22982 18092 23598
rect 18156 23254 18184 24754
rect 18248 24682 18276 25910
rect 18657 25596 18965 25605
rect 18657 25594 18663 25596
rect 18719 25594 18743 25596
rect 18799 25594 18823 25596
rect 18879 25594 18903 25596
rect 18959 25594 18965 25596
rect 18719 25542 18721 25594
rect 18901 25542 18903 25594
rect 18657 25540 18663 25542
rect 18719 25540 18743 25542
rect 18799 25540 18823 25542
rect 18879 25540 18903 25542
rect 18959 25540 18965 25542
rect 18657 25531 18965 25540
rect 18880 25492 18932 25498
rect 18880 25434 18932 25440
rect 18892 25294 18920 25434
rect 19248 25356 19300 25362
rect 19248 25298 19300 25304
rect 18880 25288 18932 25294
rect 18340 25226 18828 25242
rect 18880 25230 18932 25236
rect 19064 25288 19116 25294
rect 19064 25230 19116 25236
rect 18340 25220 18840 25226
rect 18340 25214 18788 25220
rect 18340 24886 18368 25214
rect 18788 25162 18840 25168
rect 18420 25152 18472 25158
rect 19076 25106 19104 25230
rect 18420 25094 18472 25100
rect 18432 24886 18460 25094
rect 18984 25078 19104 25106
rect 19156 25152 19208 25158
rect 19156 25094 19208 25100
rect 18328 24880 18380 24886
rect 18328 24822 18380 24828
rect 18420 24880 18472 24886
rect 18420 24822 18472 24828
rect 18984 24834 19012 25078
rect 19168 24970 19196 25094
rect 19076 24954 19196 24970
rect 19064 24948 19196 24954
rect 19116 24942 19196 24948
rect 19064 24890 19116 24896
rect 18236 24676 18288 24682
rect 18236 24618 18288 24624
rect 18144 23248 18196 23254
rect 18144 23190 18196 23196
rect 18340 23118 18368 24822
rect 18984 24806 19104 24834
rect 18657 24508 18965 24517
rect 18657 24506 18663 24508
rect 18719 24506 18743 24508
rect 18799 24506 18823 24508
rect 18879 24506 18903 24508
rect 18959 24506 18965 24508
rect 18719 24454 18721 24506
rect 18901 24454 18903 24506
rect 18657 24452 18663 24454
rect 18719 24452 18743 24454
rect 18799 24452 18823 24454
rect 18879 24452 18903 24454
rect 18959 24452 18965 24454
rect 18657 24443 18965 24452
rect 19076 24206 19104 24806
rect 19260 24410 19288 25298
rect 19352 24886 19380 25910
rect 19444 25294 19472 26250
rect 19812 25294 19840 26250
rect 19892 25356 19944 25362
rect 19892 25298 19944 25304
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19800 25288 19852 25294
rect 19800 25230 19852 25236
rect 19340 24880 19392 24886
rect 19340 24822 19392 24828
rect 19248 24404 19300 24410
rect 19248 24346 19300 24352
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 18657 23420 18965 23429
rect 18657 23418 18663 23420
rect 18719 23418 18743 23420
rect 18799 23418 18823 23420
rect 18879 23418 18903 23420
rect 18959 23418 18965 23420
rect 18719 23366 18721 23418
rect 18901 23366 18903 23418
rect 18657 23364 18663 23366
rect 18719 23364 18743 23366
rect 18799 23364 18823 23366
rect 18879 23364 18903 23366
rect 18959 23364 18965 23366
rect 18657 23355 18965 23364
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 18657 22332 18965 22341
rect 18657 22330 18663 22332
rect 18719 22330 18743 22332
rect 18799 22330 18823 22332
rect 18879 22330 18903 22332
rect 18959 22330 18965 22332
rect 18719 22278 18721 22330
rect 18901 22278 18903 22330
rect 18657 22276 18663 22278
rect 18719 22276 18743 22278
rect 18799 22276 18823 22278
rect 18879 22276 18903 22278
rect 18959 22276 18965 22278
rect 18657 22267 18965 22276
rect 18052 22092 18104 22098
rect 18052 22034 18104 22040
rect 19248 22094 19300 22098
rect 19352 22094 19380 24822
rect 19444 24614 19472 25230
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19444 24342 19472 24550
rect 19432 24336 19484 24342
rect 19432 24278 19484 24284
rect 19812 24290 19840 25230
rect 19904 24410 19932 25298
rect 20088 25226 20116 27338
rect 20732 26042 20760 27338
rect 20824 27062 20852 27474
rect 20916 27130 20944 28512
rect 21284 28422 21312 28698
rect 21376 28558 21404 28902
rect 22006 28656 22062 28665
rect 22006 28591 22062 28600
rect 21364 28552 21416 28558
rect 21364 28494 21416 28500
rect 21640 28552 21692 28558
rect 21640 28494 21692 28500
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 21376 28422 21404 28494
rect 21272 28416 21324 28422
rect 21272 28358 21324 28364
rect 21364 28416 21416 28422
rect 21364 28358 21416 28364
rect 21652 28014 21680 28494
rect 21836 28218 21864 28494
rect 22020 28422 22048 28591
rect 22112 28490 22140 29038
rect 22376 28756 22428 28762
rect 22376 28698 22428 28704
rect 22388 28558 22416 28698
rect 22376 28552 22428 28558
rect 22376 28494 22428 28500
rect 22100 28484 22152 28490
rect 22100 28426 22152 28432
rect 22652 28484 22704 28490
rect 22652 28426 22704 28432
rect 22008 28416 22060 28422
rect 22008 28358 22060 28364
rect 21824 28212 21876 28218
rect 21824 28154 21876 28160
rect 21272 28008 21324 28014
rect 21270 27976 21272 27985
rect 21640 28008 21692 28014
rect 21324 27976 21326 27985
rect 21640 27950 21692 27956
rect 21270 27911 21326 27920
rect 20996 27328 21048 27334
rect 20996 27270 21048 27276
rect 20904 27124 20956 27130
rect 20904 27066 20956 27072
rect 20812 27056 20864 27062
rect 20812 26998 20864 27004
rect 21008 26790 21036 27270
rect 20996 26784 21048 26790
rect 20996 26726 21048 26732
rect 20720 26036 20772 26042
rect 20720 25978 20772 25984
rect 20732 25786 20760 25978
rect 20732 25758 20852 25786
rect 20720 25696 20772 25702
rect 20720 25638 20772 25644
rect 20076 25220 20128 25226
rect 20076 25162 20128 25168
rect 20088 24750 20116 25162
rect 20260 24880 20312 24886
rect 20260 24822 20312 24828
rect 20076 24744 20128 24750
rect 20076 24686 20128 24692
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 19892 24404 19944 24410
rect 19892 24346 19944 24352
rect 19812 24262 19932 24290
rect 19904 24138 19932 24262
rect 20088 24206 20116 24550
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19892 24132 19944 24138
rect 19892 24074 19944 24080
rect 19904 23866 19932 24074
rect 20088 24070 20116 24142
rect 20272 24138 20300 24822
rect 20732 24818 20760 25638
rect 20824 25226 20852 25758
rect 21284 25362 21312 27911
rect 21652 27334 21680 27950
rect 22112 27538 22140 28426
rect 22198 28316 22506 28325
rect 22198 28314 22204 28316
rect 22260 28314 22284 28316
rect 22340 28314 22364 28316
rect 22420 28314 22444 28316
rect 22500 28314 22506 28316
rect 22260 28262 22262 28314
rect 22442 28262 22444 28314
rect 22198 28260 22204 28262
rect 22260 28260 22284 28262
rect 22340 28260 22364 28262
rect 22420 28260 22444 28262
rect 22500 28260 22506 28262
rect 22198 28251 22506 28260
rect 22284 28212 22336 28218
rect 22284 28154 22336 28160
rect 22192 27872 22244 27878
rect 22192 27814 22244 27820
rect 22100 27532 22152 27538
rect 22100 27474 22152 27480
rect 22008 27464 22060 27470
rect 21928 27424 22008 27452
rect 21640 27328 21692 27334
rect 21640 27270 21692 27276
rect 21928 26994 21956 27424
rect 22008 27406 22060 27412
rect 22204 27402 22232 27814
rect 22296 27470 22324 28154
rect 22664 28082 22692 28426
rect 22376 28076 22428 28082
rect 22376 28018 22428 28024
rect 22652 28076 22704 28082
rect 22652 28018 22704 28024
rect 22388 27470 22416 28018
rect 22652 27940 22704 27946
rect 22652 27882 22704 27888
rect 22560 27872 22612 27878
rect 22560 27814 22612 27820
rect 22572 27674 22600 27814
rect 22560 27668 22612 27674
rect 22560 27610 22612 27616
rect 22664 27606 22692 27882
rect 22848 27606 22876 29106
rect 23388 29096 23440 29102
rect 23388 29038 23440 29044
rect 24492 29096 24544 29102
rect 24492 29038 24544 29044
rect 23204 29028 23256 29034
rect 23204 28970 23256 28976
rect 22928 28960 22980 28966
rect 22928 28902 22980 28908
rect 23112 28960 23164 28966
rect 23112 28902 23164 28908
rect 22940 28762 22968 28902
rect 22928 28756 22980 28762
rect 22928 28698 22980 28704
rect 23124 28626 23152 28902
rect 23112 28620 23164 28626
rect 23112 28562 23164 28568
rect 23216 28150 23244 28970
rect 23400 28422 23428 29038
rect 24216 28688 24268 28694
rect 24216 28630 24268 28636
rect 24032 28552 24084 28558
rect 23860 28512 24032 28540
rect 23388 28416 23440 28422
rect 23388 28358 23440 28364
rect 23204 28144 23256 28150
rect 23204 28086 23256 28092
rect 23756 28144 23808 28150
rect 23860 28132 23888 28512
rect 24032 28494 24084 28500
rect 24228 28218 24256 28630
rect 24504 28558 24532 29038
rect 24492 28552 24544 28558
rect 24492 28494 24544 28500
rect 24676 28484 24728 28490
rect 24676 28426 24728 28432
rect 24400 28416 24452 28422
rect 24400 28358 24452 28364
rect 24216 28212 24268 28218
rect 24216 28154 24268 28160
rect 23808 28104 23888 28132
rect 23756 28086 23808 28092
rect 22652 27600 22704 27606
rect 22652 27542 22704 27548
rect 22836 27600 22888 27606
rect 22836 27542 22888 27548
rect 22284 27464 22336 27470
rect 22284 27406 22336 27412
rect 22376 27464 22428 27470
rect 22376 27406 22428 27412
rect 22192 27396 22244 27402
rect 22192 27338 22244 27344
rect 22008 27328 22060 27334
rect 22008 27270 22060 27276
rect 22020 27130 22048 27270
rect 22198 27228 22506 27237
rect 22198 27226 22204 27228
rect 22260 27226 22284 27228
rect 22340 27226 22364 27228
rect 22420 27226 22444 27228
rect 22500 27226 22506 27228
rect 22260 27174 22262 27226
rect 22442 27174 22444 27226
rect 22198 27172 22204 27174
rect 22260 27172 22284 27174
rect 22340 27172 22364 27174
rect 22420 27172 22444 27174
rect 22500 27172 22506 27174
rect 22198 27163 22506 27172
rect 22008 27124 22060 27130
rect 22008 27066 22060 27072
rect 21916 26988 21968 26994
rect 21916 26930 21968 26936
rect 22198 26140 22506 26149
rect 22198 26138 22204 26140
rect 22260 26138 22284 26140
rect 22340 26138 22364 26140
rect 22420 26138 22444 26140
rect 22500 26138 22506 26140
rect 22260 26086 22262 26138
rect 22442 26086 22444 26138
rect 22198 26084 22204 26086
rect 22260 26084 22284 26086
rect 22340 26084 22364 26086
rect 22420 26084 22444 26086
rect 22500 26084 22506 26086
rect 22198 26075 22506 26084
rect 21272 25356 21324 25362
rect 21272 25298 21324 25304
rect 20812 25220 20864 25226
rect 20812 25162 20864 25168
rect 22652 25220 22704 25226
rect 22652 25162 22704 25168
rect 22198 25052 22506 25061
rect 22198 25050 22204 25052
rect 22260 25050 22284 25052
rect 22340 25050 22364 25052
rect 22420 25050 22444 25052
rect 22500 25050 22506 25052
rect 22260 24998 22262 25050
rect 22442 24998 22444 25050
rect 22198 24996 22204 24998
rect 22260 24996 22284 24998
rect 22340 24996 22364 24998
rect 22420 24996 22444 24998
rect 22500 24996 22506 24998
rect 22198 24987 22506 24996
rect 20720 24812 20772 24818
rect 20720 24754 20772 24760
rect 20260 24132 20312 24138
rect 20260 24074 20312 24080
rect 20076 24064 20128 24070
rect 20076 24006 20128 24012
rect 19892 23860 19944 23866
rect 19892 23802 19944 23808
rect 19248 22092 19380 22094
rect 19300 22066 19380 22092
rect 19248 22034 19300 22040
rect 17682 21992 17738 22001
rect 17682 21927 17738 21936
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 17880 21146 17908 21830
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 16946 19952 17002 19961
rect 16946 19887 17002 19896
rect 16856 19780 16908 19786
rect 16856 19722 16908 19728
rect 16868 19514 16896 19722
rect 17236 19514 17264 20402
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 17512 18630 17540 20402
rect 17604 19718 17632 20402
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17972 19854 18000 20334
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17972 19242 18000 19450
rect 17960 19236 18012 19242
rect 17960 19178 18012 19184
rect 17684 18896 17736 18902
rect 17684 18838 17736 18844
rect 17696 18698 17724 18838
rect 17684 18692 17736 18698
rect 17684 18634 17736 18640
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17972 18426 18000 18566
rect 16580 18420 16632 18426
rect 16580 18362 16632 18368
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 18064 18222 18092 22034
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 18432 21690 18460 21966
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18432 21162 18460 21626
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 18657 21244 18965 21253
rect 18657 21242 18663 21244
rect 18719 21242 18743 21244
rect 18799 21242 18823 21244
rect 18879 21242 18903 21244
rect 18959 21242 18965 21244
rect 18719 21190 18721 21242
rect 18901 21190 18903 21242
rect 18657 21188 18663 21190
rect 18719 21188 18743 21190
rect 18799 21188 18823 21190
rect 18879 21188 18903 21190
rect 18959 21188 18965 21190
rect 18657 21179 18965 21188
rect 18340 21134 18460 21162
rect 18144 20868 18196 20874
rect 18144 20810 18196 20816
rect 18156 20466 18184 20810
rect 18340 20466 18368 21134
rect 19076 21128 19104 21490
rect 19168 21146 19196 21490
rect 18984 21100 19104 21128
rect 19156 21140 19208 21146
rect 18984 20874 19012 21100
rect 19156 21082 19208 21088
rect 19352 20942 19380 22066
rect 19616 21616 19668 21622
rect 19616 21558 19668 21564
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 18972 20868 19024 20874
rect 18972 20810 19024 20816
rect 19248 20868 19300 20874
rect 19248 20810 19300 20816
rect 18880 20800 18932 20806
rect 18880 20742 18932 20748
rect 19064 20800 19116 20806
rect 19064 20742 19116 20748
rect 18892 20466 18920 20742
rect 19076 20602 19104 20742
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18156 20058 18184 20402
rect 19260 20330 19288 20810
rect 18512 20324 18564 20330
rect 18512 20266 18564 20272
rect 19248 20324 19300 20330
rect 19248 20266 19300 20272
rect 18524 20058 18552 20266
rect 19444 20262 19472 21490
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19536 21146 19564 21286
rect 19628 21146 19656 21558
rect 19708 21480 19760 21486
rect 19708 21422 19760 21428
rect 19524 21140 19576 21146
rect 19524 21082 19576 21088
rect 19616 21140 19668 21146
rect 19616 21082 19668 21088
rect 19720 21010 19748 21422
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 19892 21004 19944 21010
rect 19892 20946 19944 20952
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 19524 20800 19576 20806
rect 19812 20788 19840 20878
rect 19576 20760 19840 20788
rect 19524 20742 19576 20748
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 18657 20156 18965 20165
rect 18657 20154 18663 20156
rect 18719 20154 18743 20156
rect 18799 20154 18823 20156
rect 18879 20154 18903 20156
rect 18959 20154 18965 20156
rect 18719 20102 18721 20154
rect 18901 20102 18903 20154
rect 18657 20100 18663 20102
rect 18719 20100 18743 20102
rect 18799 20100 18823 20102
rect 18879 20100 18903 20102
rect 18959 20100 18965 20102
rect 18657 20091 18965 20100
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18512 20052 18564 20058
rect 18512 19994 18564 20000
rect 18156 18426 18184 19994
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 19708 19712 19760 19718
rect 19708 19654 19760 19660
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 18657 19068 18965 19077
rect 18657 19066 18663 19068
rect 18719 19066 18743 19068
rect 18799 19066 18823 19068
rect 18879 19066 18903 19068
rect 18959 19066 18965 19068
rect 18719 19014 18721 19066
rect 18901 19014 18903 19066
rect 18657 19012 18663 19014
rect 18719 19012 18743 19014
rect 18799 19012 18823 19014
rect 18879 19012 18903 19014
rect 18959 19012 18965 19014
rect 18657 19003 18965 19012
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18800 18426 18828 18702
rect 18144 18420 18196 18426
rect 18144 18362 18196 18368
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16684 17338 16712 17478
rect 16776 17338 16804 18090
rect 18156 18034 18184 18362
rect 19076 18290 19104 19450
rect 19352 19378 19380 19654
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19444 18970 19472 19382
rect 19536 19378 19564 19654
rect 19628 19446 19656 19654
rect 19720 19514 19748 19654
rect 19904 19514 19932 20946
rect 19708 19508 19760 19514
rect 19708 19450 19760 19456
rect 19892 19508 19944 19514
rect 19892 19450 19944 19456
rect 19616 19440 19668 19446
rect 19616 19382 19668 19388
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 19720 19366 19932 19394
rect 20088 19378 20116 24006
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19156 18896 19208 18902
rect 19156 18838 19208 18844
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18328 18148 18380 18154
rect 18328 18090 18380 18096
rect 17880 18006 18184 18034
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16764 17332 16816 17338
rect 16764 17274 16816 17280
rect 17144 17202 17172 17478
rect 17604 17338 17632 17546
rect 17880 17542 17908 18006
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 18340 17202 18368 18090
rect 18418 17912 18474 17921
rect 18418 17847 18474 17856
rect 18432 17542 18460 17847
rect 18524 17660 18552 18158
rect 18657 17980 18965 17989
rect 18657 17978 18663 17980
rect 18719 17978 18743 17980
rect 18799 17978 18823 17980
rect 18879 17978 18903 17980
rect 18959 17978 18965 17980
rect 18719 17926 18721 17978
rect 18901 17926 18903 17978
rect 18657 17924 18663 17926
rect 18719 17924 18743 17926
rect 18799 17924 18823 17926
rect 18879 17924 18903 17926
rect 18959 17924 18965 17926
rect 18657 17915 18965 17924
rect 18604 17808 18656 17814
rect 18604 17750 18656 17756
rect 18616 17678 18644 17750
rect 18604 17672 18656 17678
rect 18524 17632 18604 17660
rect 18604 17614 18656 17620
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 18328 17196 18380 17202
rect 18432 17184 18460 17478
rect 19076 17338 19104 17478
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 18512 17196 18564 17202
rect 18432 17156 18512 17184
rect 18328 17138 18380 17144
rect 18512 17138 18564 17144
rect 19064 17196 19116 17202
rect 19168 17184 19196 18838
rect 19432 18692 19484 18698
rect 19432 18634 19484 18640
rect 19444 18442 19472 18634
rect 19536 18442 19564 19314
rect 19616 19304 19668 19310
rect 19720 19292 19748 19366
rect 19668 19264 19748 19292
rect 19616 19246 19668 19252
rect 19800 19236 19852 19242
rect 19800 19178 19852 19184
rect 19812 18766 19840 19178
rect 19904 18970 19932 19366
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20168 19372 20220 19378
rect 20168 19314 20220 19320
rect 20272 19334 20300 24074
rect 22198 23964 22506 23973
rect 22198 23962 22204 23964
rect 22260 23962 22284 23964
rect 22340 23962 22364 23964
rect 22420 23962 22444 23964
rect 22500 23962 22506 23964
rect 22260 23910 22262 23962
rect 22442 23910 22444 23962
rect 22198 23908 22204 23910
rect 22260 23908 22284 23910
rect 22340 23908 22364 23910
rect 22420 23908 22444 23910
rect 22500 23908 22506 23910
rect 22198 23899 22506 23908
rect 22664 23866 22692 25162
rect 22652 23860 22704 23866
rect 22652 23802 22704 23808
rect 21640 23180 21692 23186
rect 21640 23122 21692 23128
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 21178 23080 21234 23089
rect 20732 22778 20760 23054
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20824 22642 20852 23054
rect 21178 23015 21180 23024
rect 21232 23015 21234 23024
rect 21180 22986 21232 22992
rect 20996 22976 21048 22982
rect 20996 22918 21048 22924
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 20444 22568 20496 22574
rect 20444 22510 20496 22516
rect 20352 22160 20404 22166
rect 20350 22128 20352 22137
rect 20404 22128 20406 22137
rect 20350 22063 20406 22072
rect 20456 22030 20484 22510
rect 20732 22094 20760 22578
rect 20732 22066 20852 22094
rect 20824 22030 20852 22066
rect 21008 22030 21036 22918
rect 21192 22506 21220 22986
rect 21652 22658 21680 23122
rect 21732 23112 21784 23118
rect 21732 23054 21784 23060
rect 21744 22710 21772 23054
rect 22560 23044 22612 23050
rect 22560 22986 22612 22992
rect 22198 22876 22506 22885
rect 22198 22874 22204 22876
rect 22260 22874 22284 22876
rect 22340 22874 22364 22876
rect 22420 22874 22444 22876
rect 22500 22874 22506 22876
rect 22260 22822 22262 22874
rect 22442 22822 22444 22874
rect 22198 22820 22204 22822
rect 22260 22820 22284 22822
rect 22340 22820 22364 22822
rect 22420 22820 22444 22822
rect 22500 22820 22506 22822
rect 22198 22811 22506 22820
rect 21284 22642 21680 22658
rect 21732 22704 21784 22710
rect 21732 22646 21784 22652
rect 21284 22636 21692 22642
rect 21284 22630 21640 22636
rect 21180 22500 21232 22506
rect 21180 22442 21232 22448
rect 21088 22432 21140 22438
rect 21088 22374 21140 22380
rect 21100 22030 21128 22374
rect 21284 22166 21312 22630
rect 21640 22578 21692 22584
rect 21364 22568 21416 22574
rect 21364 22510 21416 22516
rect 21376 22234 21404 22510
rect 21456 22500 21508 22506
rect 21456 22442 21508 22448
rect 21640 22500 21692 22506
rect 21640 22442 21692 22448
rect 21364 22228 21416 22234
rect 21364 22170 21416 22176
rect 21272 22160 21324 22166
rect 21272 22102 21324 22108
rect 20444 22024 20496 22030
rect 20444 21966 20496 21972
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20812 22024 20864 22030
rect 20812 21966 20864 21972
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 21088 22024 21140 22030
rect 21088 21966 21140 21972
rect 20456 21894 20484 21966
rect 20444 21888 20496 21894
rect 20444 21830 20496 21836
rect 20628 21480 20680 21486
rect 20548 21440 20628 21468
rect 20548 21078 20576 21440
rect 20628 21422 20680 21428
rect 20732 21418 20760 21966
rect 20824 21690 20852 21966
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 21284 21486 21312 22102
rect 21376 21622 21404 22170
rect 21468 22030 21496 22442
rect 21548 22432 21600 22438
rect 21548 22374 21600 22380
rect 21560 22030 21588 22374
rect 21652 22234 21680 22442
rect 21744 22234 21772 22646
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 21640 22228 21692 22234
rect 21640 22170 21692 22176
rect 21732 22228 21784 22234
rect 21732 22170 21784 22176
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 21548 22024 21600 22030
rect 21548 21966 21600 21972
rect 21456 21684 21508 21690
rect 21456 21626 21508 21632
rect 21364 21616 21416 21622
rect 21364 21558 21416 21564
rect 21272 21480 21324 21486
rect 21272 21422 21324 21428
rect 21364 21480 21416 21486
rect 21468 21468 21496 21626
rect 21560 21468 21588 21966
rect 21640 21956 21692 21962
rect 21640 21898 21692 21904
rect 21652 21690 21680 21898
rect 21640 21684 21692 21690
rect 21640 21626 21692 21632
rect 21416 21440 21588 21468
rect 21364 21422 21416 21428
rect 20720 21412 20772 21418
rect 20720 21354 20772 21360
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 21364 21344 21416 21350
rect 21364 21286 21416 21292
rect 20536 21072 20588 21078
rect 20536 21014 20588 21020
rect 20640 20942 20668 21286
rect 21376 20942 21404 21286
rect 21468 21078 21496 21440
rect 21456 21072 21508 21078
rect 21456 21014 21508 21020
rect 20628 20936 20680 20942
rect 20628 20878 20680 20884
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 21364 20936 21416 20942
rect 21364 20878 21416 20884
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20548 19514 20576 20334
rect 20536 19508 20588 19514
rect 20536 19450 20588 19456
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19800 18760 19852 18766
rect 19852 18720 20024 18748
rect 19800 18702 19852 18708
rect 19444 18414 19564 18442
rect 19996 18426 20024 18720
rect 19536 18290 19564 18414
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19524 18284 19576 18290
rect 19524 18226 19576 18232
rect 19800 18284 19852 18290
rect 19800 18226 19852 18232
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19260 17338 19288 18158
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19116 17156 19196 17184
rect 19064 17138 19116 17144
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16500 16114 16528 16934
rect 16592 16658 16620 17070
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 17144 16522 17172 17138
rect 18657 16892 18965 16901
rect 18657 16890 18663 16892
rect 18719 16890 18743 16892
rect 18799 16890 18823 16892
rect 18879 16890 18903 16892
rect 18959 16890 18965 16892
rect 18719 16838 18721 16890
rect 18901 16838 18903 16890
rect 18657 16836 18663 16838
rect 18719 16836 18743 16838
rect 18799 16836 18823 16838
rect 18879 16836 18903 16838
rect 18959 16836 18965 16838
rect 18657 16827 18965 16836
rect 19076 16658 19104 17138
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 17132 16516 17184 16522
rect 17132 16458 17184 16464
rect 16488 16108 16540 16114
rect 16488 16050 16540 16056
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16408 13530 16436 15030
rect 16500 13938 16528 16050
rect 18657 15804 18965 15813
rect 18657 15802 18663 15804
rect 18719 15802 18743 15804
rect 18799 15802 18823 15804
rect 18879 15802 18903 15804
rect 18959 15802 18965 15804
rect 18719 15750 18721 15802
rect 18901 15750 18903 15802
rect 18657 15748 18663 15750
rect 18719 15748 18743 15750
rect 18799 15748 18823 15750
rect 18879 15748 18903 15750
rect 18959 15748 18965 15750
rect 18657 15739 18965 15748
rect 18512 15632 18564 15638
rect 17958 15600 18014 15609
rect 17408 15564 17460 15570
rect 18512 15574 18564 15580
rect 17958 15535 17960 15544
rect 17408 15506 17460 15512
rect 18012 15535 18014 15544
rect 17960 15506 18012 15512
rect 17420 14958 17448 15506
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16592 14414 16620 14758
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 17040 14340 17092 14346
rect 17040 14282 17092 14288
rect 16764 14272 16816 14278
rect 16684 14232 16764 14260
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16132 12646 16160 12786
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 16132 11558 16160 12174
rect 16316 11762 16344 13126
rect 16500 12918 16528 13262
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16592 12918 16620 13126
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16580 12912 16632 12918
rect 16580 12854 16632 12860
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15936 11076 15988 11082
rect 15936 11018 15988 11024
rect 15948 10606 15976 11018
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 16040 9625 16068 11086
rect 16316 10062 16344 11698
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 16408 10674 16436 11630
rect 16592 11218 16620 12718
rect 16684 12345 16712 14232
rect 16764 14214 16816 14220
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16670 12336 16726 12345
rect 16776 12306 16804 13670
rect 16868 12850 16896 13806
rect 17052 13326 17080 14282
rect 17132 13796 17184 13802
rect 17132 13738 17184 13744
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17144 12850 17172 13738
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 16670 12271 16726 12280
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16684 11626 16712 12174
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16672 11620 16724 11626
rect 16672 11562 16724 11568
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16408 10470 16436 10610
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16408 9738 16436 10406
rect 16592 10130 16620 11154
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16408 9710 16620 9738
rect 16026 9616 16082 9625
rect 16026 9551 16082 9560
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 15764 8566 15792 8978
rect 16592 8634 16620 9710
rect 16684 9500 16712 11018
rect 16776 9602 16804 12038
rect 16868 11082 16896 12786
rect 16960 12170 16988 12786
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16960 11218 16988 11494
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 16868 9722 16896 9930
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16776 9574 16896 9602
rect 16764 9512 16816 9518
rect 16684 9472 16764 9500
rect 16684 9042 16712 9472
rect 16764 9454 16816 9460
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 15752 8560 15804 8566
rect 15752 8502 15804 8508
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16408 7886 16436 8230
rect 16592 8022 16620 8570
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 16592 7886 16620 7958
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16776 7546 16804 7686
rect 16868 7546 16896 9574
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16776 7002 16804 7142
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 16868 6934 16896 7482
rect 16960 6934 16988 10406
rect 17038 9616 17094 9625
rect 17144 9602 17172 12786
rect 17328 10674 17356 13126
rect 17420 12918 17448 14894
rect 17972 14890 18000 15506
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18156 15366 18184 15438
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 18156 15026 18184 15302
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 18156 14618 18184 14758
rect 18144 14612 18196 14618
rect 18524 14600 18552 15574
rect 19064 15428 19116 15434
rect 19064 15370 19116 15376
rect 18657 14716 18965 14725
rect 18657 14714 18663 14716
rect 18719 14714 18743 14716
rect 18799 14714 18823 14716
rect 18879 14714 18903 14716
rect 18959 14714 18965 14716
rect 18719 14662 18721 14714
rect 18901 14662 18903 14714
rect 18657 14660 18663 14662
rect 18719 14660 18743 14662
rect 18799 14660 18823 14662
rect 18879 14660 18903 14662
rect 18959 14660 18965 14662
rect 18657 14651 18965 14660
rect 18524 14572 18736 14600
rect 18144 14554 18196 14560
rect 18156 13802 18184 14554
rect 18604 14408 18656 14414
rect 18524 14368 18604 14396
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18340 14074 18368 14214
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18144 13796 18196 13802
rect 18144 13738 18196 13744
rect 17868 13456 17920 13462
rect 17868 13398 17920 13404
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 17880 12434 17908 13398
rect 18156 13326 18184 13738
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 18328 13252 18380 13258
rect 18328 13194 18380 13200
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17788 12406 17908 12434
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17604 11354 17632 11494
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17094 9574 17172 9602
rect 17038 9551 17040 9560
rect 17092 9551 17094 9560
rect 17040 9522 17092 9528
rect 17130 9480 17186 9489
rect 17130 9415 17132 9424
rect 17184 9415 17186 9424
rect 17132 9386 17184 9392
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 17328 7886 17356 9046
rect 17512 8498 17540 9114
rect 17604 8634 17632 9318
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17696 8498 17724 10610
rect 17788 9466 17816 12406
rect 17868 11144 17920 11150
rect 17972 11132 18000 12582
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 18064 11354 18092 11630
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 17920 11104 18000 11132
rect 17868 11086 17920 11092
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17880 10674 17908 10950
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17880 9674 17908 10610
rect 17972 10062 18000 11104
rect 18064 10674 18092 11290
rect 18340 10674 18368 13194
rect 18432 12986 18460 13670
rect 18524 13530 18552 14368
rect 18604 14350 18656 14356
rect 18708 13938 18736 14572
rect 19076 14414 19104 15370
rect 19352 15094 19380 17682
rect 19444 17649 19472 18226
rect 19430 17640 19486 17649
rect 19430 17575 19486 17584
rect 19432 17536 19484 17542
rect 19536 17490 19564 18226
rect 19812 17882 19840 18226
rect 19800 17876 19852 17882
rect 19800 17818 19852 17824
rect 19996 17678 20024 18362
rect 20180 18358 20208 19314
rect 20272 19306 20484 19334
rect 20168 18352 20220 18358
rect 20168 18294 20220 18300
rect 20456 18290 20484 19306
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20258 17776 20314 17785
rect 20258 17711 20314 17720
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19484 17484 19564 17490
rect 19432 17478 19564 17484
rect 19444 17462 19564 17478
rect 19444 17184 19472 17462
rect 19444 17156 19656 17184
rect 19432 15428 19484 15434
rect 19432 15370 19484 15376
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 19444 14906 19472 15370
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19536 15026 19564 15302
rect 19628 15042 19656 17156
rect 19996 17116 20024 17614
rect 20272 17610 20300 17711
rect 20260 17604 20312 17610
rect 20260 17546 20312 17552
rect 20352 17604 20404 17610
rect 20352 17546 20404 17552
rect 20364 17338 20392 17546
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 19996 17088 20300 17116
rect 19984 15632 20036 15638
rect 19984 15574 20036 15580
rect 19524 15020 19576 15026
rect 19628 15020 19932 15042
rect 19628 15014 19708 15020
rect 19524 14962 19576 14968
rect 19760 15014 19932 15020
rect 19708 14962 19760 14968
rect 19352 14890 19472 14906
rect 19340 14884 19472 14890
rect 19392 14878 19472 14884
rect 19340 14826 19392 14832
rect 19352 14550 19380 14826
rect 19536 14618 19564 14962
rect 19800 14952 19852 14958
rect 19800 14894 19852 14900
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 19628 14618 19656 14758
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 19076 13841 19104 14350
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19062 13832 19118 13841
rect 19062 13767 19118 13776
rect 18657 13628 18965 13637
rect 18657 13626 18663 13628
rect 18719 13626 18743 13628
rect 18799 13626 18823 13628
rect 18879 13626 18903 13628
rect 18959 13626 18965 13628
rect 18719 13574 18721 13626
rect 18901 13574 18903 13626
rect 18657 13572 18663 13574
rect 18719 13572 18743 13574
rect 18799 13572 18823 13574
rect 18879 13572 18903 13574
rect 18959 13572 18965 13574
rect 18657 13563 18965 13572
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 18657 12540 18965 12549
rect 18657 12538 18663 12540
rect 18719 12538 18743 12540
rect 18799 12538 18823 12540
rect 18879 12538 18903 12540
rect 18959 12538 18965 12540
rect 18719 12486 18721 12538
rect 18901 12486 18903 12538
rect 18657 12484 18663 12486
rect 18719 12484 18743 12486
rect 18799 12484 18823 12486
rect 18879 12484 18903 12486
rect 18959 12484 18965 12486
rect 18657 12475 18965 12484
rect 19168 12345 19196 13874
rect 19260 13326 19288 14214
rect 19352 13938 19380 14486
rect 19628 14464 19656 14554
rect 19708 14544 19760 14550
rect 19708 14486 19760 14492
rect 19444 14436 19656 14464
rect 19444 14074 19472 14436
rect 19524 14340 19576 14346
rect 19524 14282 19576 14288
rect 19536 14074 19564 14282
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19524 14068 19576 14074
rect 19524 14010 19576 14016
rect 19720 13938 19748 14486
rect 19812 13938 19840 14894
rect 19904 14346 19932 15014
rect 19996 14550 20024 15574
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 19892 14340 19944 14346
rect 19892 14282 19944 14288
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19904 13954 19932 14282
rect 19996 14074 20024 14282
rect 20088 14278 20116 15302
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 20180 14618 20208 14894
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19800 13932 19852 13938
rect 19904 13926 20024 13954
rect 19800 13874 19852 13880
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 19352 13258 19380 13670
rect 19536 13530 19564 13874
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19628 13274 19656 13874
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19154 12336 19210 12345
rect 19154 12271 19210 12280
rect 19352 11762 19380 13194
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 18064 10266 18092 10406
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18432 10198 18460 11086
rect 18524 10810 18552 11698
rect 18657 11452 18965 11461
rect 18657 11450 18663 11452
rect 18719 11450 18743 11452
rect 18799 11450 18823 11452
rect 18879 11450 18903 11452
rect 18959 11450 18965 11452
rect 18719 11398 18721 11450
rect 18901 11398 18903 11450
rect 18657 11396 18663 11398
rect 18719 11396 18743 11398
rect 18799 11396 18823 11398
rect 18879 11396 18903 11398
rect 18959 11396 18965 11398
rect 18657 11387 18965 11396
rect 18696 11144 18748 11150
rect 18694 11112 18696 11121
rect 19248 11144 19300 11150
rect 18748 11112 18750 11121
rect 19248 11086 19300 11092
rect 18694 11047 18750 11056
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18420 10192 18472 10198
rect 18420 10134 18472 10140
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18340 9926 18368 9998
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 17880 9646 18276 9674
rect 17880 9586 17908 9646
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 18052 9580 18104 9586
rect 18104 9540 18184 9568
rect 18052 9522 18104 9528
rect 17788 9438 18092 9466
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17420 8090 17448 8434
rect 17696 8090 17724 8434
rect 17776 8288 17828 8294
rect 17776 8230 17828 8236
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17592 8016 17644 8022
rect 17406 7984 17462 7993
rect 17592 7958 17644 7964
rect 17406 7919 17462 7928
rect 17420 7886 17448 7919
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17224 7812 17276 7818
rect 17224 7754 17276 7760
rect 17236 7449 17264 7754
rect 17222 7440 17278 7449
rect 17040 7404 17092 7410
rect 17222 7375 17278 7384
rect 17328 7392 17356 7822
rect 17408 7404 17460 7410
rect 17040 7346 17092 7352
rect 17052 7274 17080 7346
rect 17040 7268 17092 7274
rect 17040 7210 17092 7216
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 16948 6928 17000 6934
rect 16948 6870 17000 6876
rect 16868 6474 16896 6870
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16776 6446 16896 6474
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 16210 4992 16266 5001
rect 16210 4927 16266 4936
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 16040 4282 16068 4626
rect 16224 4554 16252 4927
rect 16316 4826 16344 5510
rect 16396 5160 16448 5166
rect 16396 5102 16448 5108
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 16408 4622 16436 5102
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16500 4622 16528 4762
rect 16592 4622 16620 6394
rect 16776 5302 16804 6446
rect 16856 6384 16908 6390
rect 16856 6326 16908 6332
rect 16764 5296 16816 5302
rect 16764 5238 16816 5244
rect 16868 5030 16896 6326
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16212 4548 16264 4554
rect 16212 4490 16264 4496
rect 16304 4548 16356 4554
rect 16304 4490 16356 4496
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 15568 4276 15620 4282
rect 15568 4218 15620 4224
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 16028 4276 16080 4282
rect 16028 4218 16080 4224
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 13596 3624 13952 3652
rect 13544 3606 13596 3612
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13452 3528 13504 3534
rect 13820 3528 13872 3534
rect 13452 3470 13504 3476
rect 13556 3476 13820 3482
rect 13556 3470 13872 3476
rect 13372 2922 13400 3470
rect 13556 3454 13860 3470
rect 13924 3466 13952 3624
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 13912 3460 13964 3466
rect 13556 3058 13584 3454
rect 13912 3402 13964 3408
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13360 2916 13412 2922
rect 13360 2858 13412 2864
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13556 2446 13584 2994
rect 13740 2854 13768 3334
rect 13924 3058 13952 3402
rect 14016 3058 14044 3606
rect 14108 3602 14136 4014
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14108 3126 14136 3538
rect 14200 3534 14228 4218
rect 14280 4208 14332 4214
rect 14332 4156 14412 4162
rect 14280 4150 14412 4156
rect 14292 4134 14412 4150
rect 14384 4060 14412 4134
rect 14464 4072 14516 4078
rect 14384 4032 14464 4060
rect 14280 3732 14332 3738
rect 14384 3720 14412 4032
rect 14464 4014 14516 4020
rect 15568 4004 15620 4010
rect 15568 3946 15620 3952
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14568 3754 14596 3878
rect 14332 3692 14412 3720
rect 14280 3674 14332 3680
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14384 3398 14412 3692
rect 14476 3726 14596 3754
rect 15580 3738 15608 3946
rect 15568 3732 15620 3738
rect 14476 3534 14504 3726
rect 15568 3674 15620 3680
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 14556 3664 14608 3670
rect 14556 3606 14608 3612
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 14292 3058 14320 3334
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14476 2854 14504 3470
rect 14568 3194 14596 3606
rect 15212 3505 15240 3606
rect 15198 3496 15254 3505
rect 15198 3431 15254 3440
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 14660 3058 14688 3334
rect 14936 3126 14964 3334
rect 15115 3292 15423 3301
rect 15115 3290 15121 3292
rect 15177 3290 15201 3292
rect 15257 3290 15281 3292
rect 15337 3290 15361 3292
rect 15417 3290 15423 3292
rect 15177 3238 15179 3290
rect 15359 3238 15361 3290
rect 15115 3236 15121 3238
rect 15177 3236 15201 3238
rect 15257 3236 15281 3238
rect 15337 3236 15361 3238
rect 15417 3236 15423 3238
rect 15115 3227 15423 3236
rect 15672 3194 15700 3674
rect 15856 3602 15884 4218
rect 16316 4146 16344 4490
rect 16592 4146 16620 4558
rect 16868 4486 16896 4966
rect 16960 4826 16988 5850
rect 17052 5778 17080 7210
rect 17236 6798 17264 7375
rect 17328 7364 17408 7392
rect 17408 7346 17460 7352
rect 17500 7404 17552 7410
rect 17604 7392 17632 7958
rect 17696 7410 17724 8026
rect 17552 7364 17632 7392
rect 17684 7404 17736 7410
rect 17500 7346 17552 7352
rect 17684 7346 17736 7352
rect 17788 7274 17816 8230
rect 17972 7886 18000 9318
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17972 7546 18000 7822
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17866 7440 17922 7449
rect 18064 7410 18092 9438
rect 18156 9364 18184 9540
rect 18248 9466 18276 9646
rect 18340 9586 18368 9862
rect 18524 9722 18552 10746
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 18708 10452 18736 10610
rect 19064 10464 19116 10470
rect 18708 10424 19064 10452
rect 19064 10406 19116 10412
rect 18657 10364 18965 10373
rect 18657 10362 18663 10364
rect 18719 10362 18743 10364
rect 18799 10362 18823 10364
rect 18879 10362 18903 10364
rect 18959 10362 18965 10364
rect 18719 10310 18721 10362
rect 18901 10310 18903 10362
rect 18657 10308 18663 10310
rect 18719 10308 18743 10310
rect 18799 10308 18823 10310
rect 18879 10308 18903 10310
rect 18959 10308 18965 10310
rect 18657 10299 18965 10308
rect 19168 10130 19196 10610
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 18512 9716 18564 9722
rect 18512 9658 18564 9664
rect 19076 9586 19104 9862
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 18432 9466 18460 9522
rect 18248 9438 18460 9466
rect 18156 9336 18368 9364
rect 18340 8974 18368 9336
rect 18657 9276 18965 9285
rect 18657 9274 18663 9276
rect 18719 9274 18743 9276
rect 18799 9274 18823 9276
rect 18879 9274 18903 9276
rect 18959 9274 18965 9276
rect 18719 9222 18721 9274
rect 18901 9222 18903 9274
rect 18657 9220 18663 9222
rect 18719 9220 18743 9222
rect 18799 9220 18823 9222
rect 18879 9220 18903 9222
rect 18959 9220 18965 9222
rect 18657 9211 18965 9220
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18236 8900 18288 8906
rect 18236 8842 18288 8848
rect 18248 8362 18276 8842
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18524 8634 18552 8774
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 19260 8566 19288 11086
rect 19352 11014 19380 11698
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19444 11150 19472 11494
rect 19536 11286 19564 13262
rect 19628 13246 19932 13274
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19616 12980 19668 12986
rect 19616 12922 19668 12928
rect 19524 11280 19576 11286
rect 19524 11222 19576 11228
rect 19628 11150 19656 12922
rect 19720 12238 19748 13126
rect 19904 12434 19932 13246
rect 19996 12986 20024 13926
rect 20166 13832 20222 13841
rect 20166 13767 20222 13776
rect 20180 13734 20208 13767
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20272 13462 20300 17088
rect 20456 16794 20484 18226
rect 20732 17882 20760 18226
rect 21100 18154 21128 20402
rect 21284 20330 21312 20878
rect 21468 20380 21496 21014
rect 21548 21004 21600 21010
rect 21548 20946 21600 20952
rect 21560 20534 21588 20946
rect 21744 20942 21772 22170
rect 22112 22030 22140 22374
rect 22572 22234 22600 22986
rect 22560 22228 22612 22234
rect 22560 22170 22612 22176
rect 22572 22098 22600 22170
rect 22664 22148 22692 23802
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23492 22778 23520 22918
rect 23480 22772 23532 22778
rect 23480 22714 23532 22720
rect 22836 22704 22888 22710
rect 22836 22646 22888 22652
rect 22848 22438 22876 22646
rect 23020 22636 23072 22642
rect 23296 22636 23348 22642
rect 23020 22578 23072 22584
rect 23124 22596 23296 22624
rect 22744 22432 22796 22438
rect 22744 22374 22796 22380
rect 22836 22432 22888 22438
rect 22836 22374 22888 22380
rect 22756 22250 22784 22374
rect 22756 22222 22876 22250
rect 22664 22120 22784 22148
rect 22560 22092 22612 22098
rect 22560 22034 22612 22040
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 22198 21788 22506 21797
rect 22198 21786 22204 21788
rect 22260 21786 22284 21788
rect 22340 21786 22364 21788
rect 22420 21786 22444 21788
rect 22500 21786 22506 21788
rect 22260 21734 22262 21786
rect 22442 21734 22444 21786
rect 22198 21732 22204 21734
rect 22260 21732 22284 21734
rect 22340 21732 22364 21734
rect 22420 21732 22444 21734
rect 22500 21732 22506 21734
rect 22198 21723 22506 21732
rect 22572 21622 22600 21830
rect 22560 21616 22612 21622
rect 21822 21584 21878 21593
rect 22560 21558 22612 21564
rect 21822 21519 21878 21528
rect 22008 21548 22060 21554
rect 21836 21418 21864 21519
rect 22008 21490 22060 21496
rect 21824 21412 21876 21418
rect 21824 21354 21876 21360
rect 21732 20936 21784 20942
rect 21732 20878 21784 20884
rect 21548 20528 21600 20534
rect 21548 20470 21600 20476
rect 22020 20398 22048 21490
rect 22560 21480 22612 21486
rect 22560 21422 22612 21428
rect 22190 21176 22246 21185
rect 22112 21134 22190 21162
rect 22112 20942 22140 21134
rect 22190 21111 22246 21120
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 22198 20700 22506 20709
rect 22198 20698 22204 20700
rect 22260 20698 22284 20700
rect 22340 20698 22364 20700
rect 22420 20698 22444 20700
rect 22500 20698 22506 20700
rect 22260 20646 22262 20698
rect 22442 20646 22444 20698
rect 22198 20644 22204 20646
rect 22260 20644 22284 20646
rect 22340 20644 22364 20646
rect 22420 20644 22444 20646
rect 22500 20644 22506 20646
rect 22198 20635 22506 20644
rect 22572 20602 22600 21422
rect 22652 21344 22704 21350
rect 22652 21286 22704 21292
rect 22664 20942 22692 21286
rect 22652 20936 22704 20942
rect 22652 20878 22704 20884
rect 22664 20806 22692 20878
rect 22652 20800 22704 20806
rect 22652 20742 22704 20748
rect 22664 20602 22692 20742
rect 22560 20596 22612 20602
rect 22560 20538 22612 20544
rect 22652 20596 22704 20602
rect 22652 20538 22704 20544
rect 21548 20392 21600 20398
rect 21468 20352 21548 20380
rect 21548 20334 21600 20340
rect 22008 20392 22060 20398
rect 22008 20334 22060 20340
rect 21272 20324 21324 20330
rect 21272 20266 21324 20272
rect 21284 19174 21312 20266
rect 22664 20058 22692 20538
rect 22652 20052 22704 20058
rect 22652 19994 22704 20000
rect 22198 19612 22506 19621
rect 22198 19610 22204 19612
rect 22260 19610 22284 19612
rect 22340 19610 22364 19612
rect 22420 19610 22444 19612
rect 22500 19610 22506 19612
rect 22260 19558 22262 19610
rect 22442 19558 22444 19610
rect 22198 19556 22204 19558
rect 22260 19556 22284 19558
rect 22340 19556 22364 19558
rect 22420 19556 22444 19558
rect 22500 19556 22506 19558
rect 22198 19547 22506 19556
rect 22560 19440 22612 19446
rect 22560 19382 22612 19388
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 22198 18524 22506 18533
rect 22198 18522 22204 18524
rect 22260 18522 22284 18524
rect 22340 18522 22364 18524
rect 22420 18522 22444 18524
rect 22500 18522 22506 18524
rect 22260 18470 22262 18522
rect 22442 18470 22444 18522
rect 22198 18468 22204 18470
rect 22260 18468 22284 18470
rect 22340 18468 22364 18470
rect 22420 18468 22444 18470
rect 22500 18468 22506 18470
rect 22198 18459 22506 18468
rect 21088 18148 21140 18154
rect 21088 18090 21140 18096
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 21824 17876 21876 17882
rect 21824 17818 21876 17824
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 21836 17610 21864 17818
rect 22480 17678 22508 17818
rect 22572 17678 22600 19382
rect 22756 17954 22784 22120
rect 22848 21978 22876 22222
rect 22848 21962 22968 21978
rect 22848 21956 22980 21962
rect 22848 21950 22928 21956
rect 22848 21622 22876 21950
rect 22928 21898 22980 21904
rect 22836 21616 22888 21622
rect 22836 21558 22888 21564
rect 22928 21480 22980 21486
rect 22928 21422 22980 21428
rect 22836 21412 22888 21418
rect 22836 21354 22888 21360
rect 22848 20602 22876 21354
rect 22940 21185 22968 21422
rect 22926 21176 22982 21185
rect 22926 21111 22982 21120
rect 23032 21010 23060 22578
rect 23020 21004 23072 21010
rect 23020 20946 23072 20952
rect 23020 20868 23072 20874
rect 23124 20856 23152 22596
rect 23296 22578 23348 22584
rect 23388 22568 23440 22574
rect 23388 22510 23440 22516
rect 23204 22432 23256 22438
rect 23204 22374 23256 22380
rect 23216 22030 23244 22374
rect 23400 22098 23428 22510
rect 23388 22092 23440 22098
rect 23388 22034 23440 22040
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 23216 21418 23244 21966
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23308 21690 23336 21830
rect 23492 21690 23520 22714
rect 23572 22636 23624 22642
rect 23572 22578 23624 22584
rect 23584 22098 23612 22578
rect 23572 22092 23624 22098
rect 23572 22034 23624 22040
rect 23296 21684 23348 21690
rect 23296 21626 23348 21632
rect 23480 21684 23532 21690
rect 23480 21626 23532 21632
rect 23204 21412 23256 21418
rect 23204 21354 23256 21360
rect 23072 20828 23152 20856
rect 23020 20810 23072 20816
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 23124 20330 23152 20828
rect 23308 20602 23336 21626
rect 23388 21480 23440 21486
rect 23388 21422 23440 21428
rect 23480 21480 23532 21486
rect 23480 21422 23532 21428
rect 23400 21146 23428 21422
rect 23492 21185 23520 21422
rect 23478 21176 23534 21185
rect 23388 21140 23440 21146
rect 23478 21111 23534 21120
rect 23388 21082 23440 21088
rect 23584 21078 23612 22034
rect 23768 21162 23796 28086
rect 24412 27470 24440 28358
rect 24688 28218 24716 28426
rect 24676 28212 24728 28218
rect 24676 28154 24728 28160
rect 24400 27464 24452 27470
rect 24400 27406 24452 27412
rect 25240 23322 25268 29582
rect 25228 23316 25280 23322
rect 25228 23258 25280 23264
rect 24308 23180 24360 23186
rect 24308 23122 24360 23128
rect 25044 23180 25096 23186
rect 25044 23122 25096 23128
rect 24124 22976 24176 22982
rect 24124 22918 24176 22924
rect 24136 22642 24164 22918
rect 24320 22642 24348 23122
rect 24492 23112 24544 23118
rect 24492 23054 24544 23060
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 24308 22636 24360 22642
rect 24308 22578 24360 22584
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24216 22568 24268 22574
rect 24412 22545 24440 22578
rect 24216 22510 24268 22516
rect 24398 22536 24454 22545
rect 24032 22500 24084 22506
rect 24032 22442 24084 22448
rect 23848 22160 23900 22166
rect 23848 22102 23900 22108
rect 23860 21350 23888 22102
rect 24044 21622 24072 22442
rect 24228 22234 24256 22510
rect 24398 22471 24454 22480
rect 24216 22228 24268 22234
rect 24216 22170 24268 22176
rect 24228 21894 24256 22170
rect 24308 22160 24360 22166
rect 24308 22102 24360 22108
rect 24216 21888 24268 21894
rect 24216 21830 24268 21836
rect 24124 21684 24176 21690
rect 24124 21626 24176 21632
rect 24032 21616 24084 21622
rect 24032 21558 24084 21564
rect 23848 21344 23900 21350
rect 23848 21286 23900 21292
rect 23768 21134 23888 21162
rect 23572 21072 23624 21078
rect 23572 21014 23624 21020
rect 23756 20936 23808 20942
rect 23756 20878 23808 20884
rect 23296 20596 23348 20602
rect 23296 20538 23348 20544
rect 23768 20466 23796 20878
rect 23756 20460 23808 20466
rect 23756 20402 23808 20408
rect 23112 20324 23164 20330
rect 23112 20266 23164 20272
rect 23768 20262 23796 20402
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23388 19780 23440 19786
rect 23388 19722 23440 19728
rect 23296 18692 23348 18698
rect 23296 18634 23348 18640
rect 23204 18216 23256 18222
rect 23204 18158 23256 18164
rect 22664 17926 22784 17954
rect 22664 17882 22692 17926
rect 23216 17882 23244 18158
rect 22652 17876 22704 17882
rect 22652 17818 22704 17824
rect 22836 17876 22888 17882
rect 22836 17818 22888 17824
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 22468 17672 22520 17678
rect 22468 17614 22520 17620
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 21824 17604 21876 17610
rect 21824 17546 21876 17552
rect 21836 17202 21864 17546
rect 22198 17436 22506 17445
rect 22198 17434 22204 17436
rect 22260 17434 22284 17436
rect 22340 17434 22364 17436
rect 22420 17434 22444 17436
rect 22500 17434 22506 17436
rect 22260 17382 22262 17434
rect 22442 17382 22444 17434
rect 22198 17380 22204 17382
rect 22260 17380 22284 17382
rect 22340 17380 22364 17382
rect 22420 17380 22444 17382
rect 22500 17380 22506 17382
rect 22198 17371 22506 17380
rect 22572 17270 22600 17614
rect 22560 17264 22612 17270
rect 22560 17206 22612 17212
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 21836 16658 21864 17138
rect 22204 16794 22232 17138
rect 22284 17060 22336 17066
rect 22284 17002 22336 17008
rect 22296 16794 22324 17002
rect 22572 16794 22600 17206
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22560 16788 22612 16794
rect 22560 16730 22612 16736
rect 21824 16652 21876 16658
rect 21824 16594 21876 16600
rect 22664 16590 22692 17682
rect 22848 17354 22876 17818
rect 23308 17678 23336 18634
rect 23400 17882 23428 19722
rect 23860 18612 23888 21134
rect 23940 21140 23992 21146
rect 23940 21082 23992 21088
rect 23952 20466 23980 21082
rect 24136 21026 24164 21626
rect 24228 21146 24256 21830
rect 24216 21140 24268 21146
rect 24216 21082 24268 21088
rect 24136 20998 24256 21026
rect 24124 20936 24176 20942
rect 24124 20878 24176 20884
rect 24032 20800 24084 20806
rect 24032 20742 24084 20748
rect 24044 20466 24072 20742
rect 24136 20466 24164 20878
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 24032 20460 24084 20466
rect 24032 20402 24084 20408
rect 24124 20460 24176 20466
rect 24124 20402 24176 20408
rect 23940 18624 23992 18630
rect 23860 18584 23940 18612
rect 23940 18566 23992 18572
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 23388 17876 23440 17882
rect 23388 17818 23440 17824
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 23112 17536 23164 17542
rect 23112 17478 23164 17484
rect 22848 17338 22968 17354
rect 22836 17332 22968 17338
rect 22888 17326 22968 17332
rect 22836 17274 22888 17280
rect 22836 17196 22888 17202
rect 22836 17138 22888 17144
rect 22848 16794 22876 17138
rect 22836 16788 22888 16794
rect 22836 16730 22888 16736
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22198 16348 22506 16357
rect 22198 16346 22204 16348
rect 22260 16346 22284 16348
rect 22340 16346 22364 16348
rect 22420 16346 22444 16348
rect 22500 16346 22506 16348
rect 22260 16294 22262 16346
rect 22442 16294 22444 16346
rect 22198 16292 22204 16294
rect 22260 16292 22284 16294
rect 22340 16292 22364 16294
rect 22420 16292 22444 16294
rect 22500 16292 22506 16294
rect 22198 16283 22506 16292
rect 22848 16250 22876 16730
rect 22836 16244 22888 16250
rect 22836 16186 22888 16192
rect 22652 15564 22704 15570
rect 22652 15506 22704 15512
rect 22198 15260 22506 15269
rect 22198 15258 22204 15260
rect 22260 15258 22284 15260
rect 22340 15258 22364 15260
rect 22420 15258 22444 15260
rect 22500 15258 22506 15260
rect 22260 15206 22262 15258
rect 22442 15206 22444 15258
rect 22198 15204 22204 15206
rect 22260 15204 22284 15206
rect 22340 15204 22364 15206
rect 22420 15204 22444 15206
rect 22500 15204 22506 15206
rect 22198 15195 22506 15204
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20536 14408 20588 14414
rect 20588 14368 20668 14396
rect 20536 14350 20588 14356
rect 20640 14090 20668 14368
rect 20456 14074 20668 14090
rect 20456 14068 20680 14074
rect 20456 14062 20628 14068
rect 20456 13530 20484 14062
rect 20628 14010 20680 14016
rect 20824 13938 20852 15098
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20812 13932 20864 13938
rect 20812 13874 20864 13880
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20260 13456 20312 13462
rect 20260 13398 20312 13404
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 20732 12850 20760 13874
rect 20824 12918 20852 13874
rect 20812 12912 20864 12918
rect 20812 12854 20864 12860
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 21468 12730 21496 14962
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21560 14414 21588 14758
rect 22664 14550 22692 15506
rect 22940 15026 22968 17326
rect 23124 16998 23152 17478
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 23308 16726 23336 17614
rect 23492 17202 23520 18294
rect 23664 18216 23716 18222
rect 23664 18158 23716 18164
rect 23572 17604 23624 17610
rect 23572 17546 23624 17552
rect 23584 17338 23612 17546
rect 23572 17332 23624 17338
rect 23572 17274 23624 17280
rect 23676 17270 23704 18158
rect 23756 17740 23808 17746
rect 23756 17682 23808 17688
rect 23664 17264 23716 17270
rect 23664 17206 23716 17212
rect 23480 17196 23532 17202
rect 23480 17138 23532 17144
rect 23388 17128 23440 17134
rect 23388 17070 23440 17076
rect 23296 16720 23348 16726
rect 23296 16662 23348 16668
rect 23112 16448 23164 16454
rect 23112 16390 23164 16396
rect 23204 16448 23256 16454
rect 23204 16390 23256 16396
rect 23124 15570 23152 16390
rect 23216 16182 23244 16390
rect 23204 16176 23256 16182
rect 23204 16118 23256 16124
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 22928 15020 22980 15026
rect 22928 14962 22980 14968
rect 23020 14816 23072 14822
rect 23020 14758 23072 14764
rect 23124 14770 23152 15506
rect 23216 15502 23244 16118
rect 23400 15978 23428 17070
rect 23388 15972 23440 15978
rect 23388 15914 23440 15920
rect 23296 15632 23348 15638
rect 23296 15574 23348 15580
rect 23204 15496 23256 15502
rect 23204 15438 23256 15444
rect 23308 15026 23336 15574
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 22652 14544 22704 14550
rect 22652 14486 22704 14492
rect 22836 14476 22888 14482
rect 22836 14418 22888 14424
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 22560 14408 22612 14414
rect 22560 14350 22612 14356
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 21560 12850 21588 14350
rect 21652 12986 21680 14350
rect 21916 14340 21968 14346
rect 21916 14282 21968 14288
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21744 13326 21772 13670
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21824 13184 21876 13190
rect 21824 13126 21876 13132
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 21548 12844 21600 12850
rect 21548 12786 21600 12792
rect 19904 12406 20024 12434
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19812 11354 19840 12038
rect 19996 11898 20024 12406
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19616 11144 19668 11150
rect 19616 11086 19668 11092
rect 19996 11082 20024 11834
rect 20272 11626 20300 12718
rect 21468 12702 21588 12730
rect 21560 12646 21588 12702
rect 21652 12646 21680 12922
rect 21836 12850 21864 13126
rect 21824 12844 21876 12850
rect 21824 12786 21876 12792
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20076 11620 20128 11626
rect 20076 11562 20128 11568
rect 20260 11620 20312 11626
rect 20260 11562 20312 11568
rect 19984 11076 20036 11082
rect 19984 11018 20036 11024
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 20088 10742 20116 11562
rect 19892 10736 19944 10742
rect 19892 10678 19944 10684
rect 20076 10736 20128 10742
rect 20076 10678 20128 10684
rect 19904 10169 19932 10678
rect 19890 10160 19946 10169
rect 19890 10095 19946 10104
rect 20088 10062 20116 10678
rect 20272 10674 20300 11562
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 20272 10470 20300 10610
rect 20364 10606 20392 11698
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 20536 11008 20588 11014
rect 20536 10950 20588 10956
rect 20352 10600 20404 10606
rect 20352 10542 20404 10548
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20272 10130 20300 10406
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20364 10062 20392 10542
rect 20548 10266 20576 10950
rect 21468 10810 21496 11494
rect 21560 11150 21588 12582
rect 21732 11824 21784 11830
rect 21732 11766 21784 11772
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 21548 11144 21600 11150
rect 21546 11112 21548 11121
rect 21600 11112 21602 11121
rect 21546 11047 21602 11056
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 21652 10062 21680 11290
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 21640 10056 21692 10062
rect 21640 9998 21692 10004
rect 21744 9722 21772 11766
rect 21928 11354 21956 14282
rect 22198 14172 22506 14181
rect 22198 14170 22204 14172
rect 22260 14170 22284 14172
rect 22340 14170 22364 14172
rect 22420 14170 22444 14172
rect 22500 14170 22506 14172
rect 22260 14118 22262 14170
rect 22442 14118 22444 14170
rect 22198 14116 22204 14118
rect 22260 14116 22284 14118
rect 22340 14116 22364 14118
rect 22420 14116 22444 14118
rect 22500 14116 22506 14118
rect 22198 14107 22506 14116
rect 22572 14074 22600 14350
rect 22560 14068 22612 14074
rect 22560 14010 22612 14016
rect 22192 13864 22244 13870
rect 22192 13806 22244 13812
rect 22204 13394 22232 13806
rect 22664 13394 22692 14350
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22198 13084 22506 13093
rect 22198 13082 22204 13084
rect 22260 13082 22284 13084
rect 22340 13082 22364 13084
rect 22420 13082 22444 13084
rect 22500 13082 22506 13084
rect 22260 13030 22262 13082
rect 22442 13030 22444 13082
rect 22198 13028 22204 13030
rect 22260 13028 22284 13030
rect 22340 13028 22364 13030
rect 22420 13028 22444 13030
rect 22500 13028 22506 13030
rect 22198 13019 22506 13028
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22744 12776 22796 12782
rect 22744 12718 22796 12724
rect 22204 12238 22232 12718
rect 22652 12708 22704 12714
rect 22652 12650 22704 12656
rect 22664 12238 22692 12650
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22198 11996 22506 12005
rect 22198 11994 22204 11996
rect 22260 11994 22284 11996
rect 22340 11994 22364 11996
rect 22420 11994 22444 11996
rect 22500 11994 22506 11996
rect 22260 11942 22262 11994
rect 22442 11942 22444 11994
rect 22198 11940 22204 11942
rect 22260 11940 22284 11942
rect 22340 11940 22364 11942
rect 22420 11940 22444 11942
rect 22500 11940 22506 11942
rect 22198 11931 22506 11940
rect 22664 11762 22692 12038
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 22652 11756 22704 11762
rect 22652 11698 22704 11704
rect 21916 11348 21968 11354
rect 21916 11290 21968 11296
rect 22112 11150 22140 11698
rect 22572 11626 22600 11698
rect 22560 11620 22612 11626
rect 22560 11562 22612 11568
rect 22572 11150 22600 11562
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22008 11076 22060 11082
rect 22008 11018 22060 11024
rect 22020 10810 22048 11018
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 22112 10674 22140 11086
rect 22198 10908 22506 10917
rect 22198 10906 22204 10908
rect 22260 10906 22284 10908
rect 22340 10906 22364 10908
rect 22420 10906 22444 10908
rect 22500 10906 22506 10908
rect 22260 10854 22262 10906
rect 22442 10854 22444 10906
rect 22198 10852 22204 10854
rect 22260 10852 22284 10854
rect 22340 10852 22364 10854
rect 22420 10852 22444 10854
rect 22500 10852 22506 10854
rect 22198 10843 22506 10852
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 22572 10470 22600 11086
rect 22664 10606 22692 11698
rect 22756 11082 22784 12718
rect 22848 12345 22876 14418
rect 22928 14408 22980 14414
rect 22928 14350 22980 14356
rect 22940 13530 22968 14350
rect 22928 13524 22980 13530
rect 22928 13466 22980 13472
rect 23032 13410 23060 14758
rect 23124 14742 23336 14770
rect 23112 14340 23164 14346
rect 23112 14282 23164 14288
rect 23124 14074 23152 14282
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 23124 13546 23152 14010
rect 23124 13518 23244 13546
rect 23032 13382 23152 13410
rect 22928 12776 22980 12782
rect 22928 12718 22980 12724
rect 22940 12434 22968 12718
rect 22940 12406 23060 12434
rect 22928 12368 22980 12374
rect 22834 12336 22890 12345
rect 22928 12310 22980 12316
rect 22834 12271 22890 12280
rect 22848 12102 22876 12271
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22940 11694 22968 12310
rect 23032 12306 23060 12406
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 23020 12164 23072 12170
rect 23020 12106 23072 12112
rect 22928 11688 22980 11694
rect 22928 11630 22980 11636
rect 22744 11076 22796 11082
rect 22744 11018 22796 11024
rect 22836 11076 22888 11082
rect 22836 11018 22888 11024
rect 22652 10600 22704 10606
rect 22652 10542 22704 10548
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22652 10464 22704 10470
rect 22652 10406 22704 10412
rect 22756 10418 22784 11018
rect 22848 10538 22876 11018
rect 23032 10810 23060 12106
rect 23020 10804 23072 10810
rect 23020 10746 23072 10752
rect 22836 10532 22888 10538
rect 22836 10474 22888 10480
rect 22928 10464 22980 10470
rect 22756 10412 22928 10418
rect 22756 10406 22980 10412
rect 22112 10266 22140 10406
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 22388 10198 22416 10406
rect 22664 10266 22692 10406
rect 22756 10390 22968 10406
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22376 10192 22428 10198
rect 22376 10134 22428 10140
rect 22560 10192 22612 10198
rect 22560 10134 22612 10140
rect 22650 10160 22706 10169
rect 22572 9994 22600 10134
rect 22650 10095 22706 10104
rect 22664 10062 22692 10095
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22560 9988 22612 9994
rect 22560 9930 22612 9936
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 21732 9716 21784 9722
rect 21732 9658 21784 9664
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19352 8974 19380 9318
rect 22112 8974 22140 9862
rect 22198 9820 22506 9829
rect 22198 9818 22204 9820
rect 22260 9818 22284 9820
rect 22340 9818 22364 9820
rect 22420 9818 22444 9820
rect 22500 9818 22506 9820
rect 22260 9766 22262 9818
rect 22442 9766 22444 9818
rect 22198 9764 22204 9766
rect 22260 9764 22284 9766
rect 22340 9764 22364 9766
rect 22420 9764 22444 9766
rect 22500 9764 22506 9766
rect 22198 9755 22506 9764
rect 22572 9042 22600 9930
rect 22652 9580 22704 9586
rect 22652 9522 22704 9528
rect 22664 9042 22692 9522
rect 22376 9036 22428 9042
rect 22376 8978 22428 8984
rect 22560 9036 22612 9042
rect 22560 8978 22612 8984
rect 22652 9036 22704 9042
rect 22652 8978 22704 8984
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 22100 8968 22152 8974
rect 22100 8910 22152 8916
rect 22388 8838 22416 8978
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 21732 8832 21784 8838
rect 21732 8774 21784 8780
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 22376 8832 22428 8838
rect 22376 8774 22428 8780
rect 20640 8634 20668 8774
rect 21744 8634 21772 8774
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 20812 8288 20864 8294
rect 20812 8230 20864 8236
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 18657 8188 18965 8197
rect 18657 8186 18663 8188
rect 18719 8186 18743 8188
rect 18799 8186 18823 8188
rect 18879 8186 18903 8188
rect 18959 8186 18965 8188
rect 18719 8134 18721 8186
rect 18901 8134 18903 8186
rect 18657 8132 18663 8134
rect 18719 8132 18743 8134
rect 18799 8132 18823 8134
rect 18879 8132 18903 8134
rect 18959 8132 18965 8134
rect 18657 8123 18965 8132
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 17866 7375 17868 7384
rect 17920 7375 17922 7384
rect 18052 7404 18104 7410
rect 17868 7346 17920 7352
rect 18052 7346 18104 7352
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17420 6798 17448 7142
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 17500 6928 17552 6934
rect 17500 6870 17552 6876
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 17052 5137 17080 5170
rect 17038 5128 17094 5137
rect 17038 5063 17094 5072
rect 17144 5030 17172 6598
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17236 5370 17264 5782
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16868 4282 16896 4422
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16960 4146 16988 4762
rect 17052 4690 17080 4966
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 17328 4570 17356 5306
rect 17420 5234 17448 5714
rect 17512 5642 17540 6870
rect 17604 6730 17632 6938
rect 17592 6724 17644 6730
rect 17592 6666 17644 6672
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17788 6458 17816 6598
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17880 6390 17908 7142
rect 18064 6662 18092 7346
rect 18340 7206 18368 7686
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 17972 6458 18000 6598
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17868 6384 17920 6390
rect 17868 6326 17920 6332
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17500 5636 17552 5642
rect 17500 5578 17552 5584
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17604 4826 17632 6054
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17684 5296 17736 5302
rect 17684 5238 17736 5244
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17052 4542 17356 4570
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 16028 4140 16080 4146
rect 16028 4082 16080 4088
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16040 3942 16068 4082
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 16592 3534 16620 4082
rect 17052 3942 17080 4542
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 17236 4146 17264 4422
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17420 4078 17448 4558
rect 17592 4548 17644 4554
rect 17592 4490 17644 4496
rect 17408 4072 17460 4078
rect 17408 4014 17460 4020
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 17052 3534 17080 3878
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17144 3380 17172 3878
rect 17052 3352 17172 3380
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 17052 3058 17080 3352
rect 17420 3074 17448 4014
rect 17604 3602 17632 4490
rect 17696 4486 17724 5238
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17788 4282 17816 5510
rect 17880 5234 17908 6326
rect 18340 5710 18368 7142
rect 18657 7100 18965 7109
rect 18657 7098 18663 7100
rect 18719 7098 18743 7100
rect 18799 7098 18823 7100
rect 18879 7098 18903 7100
rect 18959 7098 18965 7100
rect 18719 7046 18721 7098
rect 18901 7046 18903 7098
rect 18657 7044 18663 7046
rect 18719 7044 18743 7046
rect 18799 7044 18823 7046
rect 18879 7044 18903 7046
rect 18959 7044 18965 7046
rect 18657 7035 18965 7044
rect 20088 6866 20116 7822
rect 20824 7818 20852 8230
rect 20916 7954 20944 8230
rect 22112 8090 22140 8774
rect 22198 8732 22506 8741
rect 22198 8730 22204 8732
rect 22260 8730 22284 8732
rect 22340 8730 22364 8732
rect 22420 8730 22444 8732
rect 22500 8730 22506 8732
rect 22260 8678 22262 8730
rect 22442 8678 22444 8730
rect 22198 8676 22204 8678
rect 22260 8676 22284 8678
rect 22340 8676 22364 8678
rect 22420 8676 22444 8678
rect 22500 8676 22506 8678
rect 22198 8667 22506 8676
rect 22572 8616 22600 8978
rect 22296 8588 22600 8616
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 22204 7834 22232 8026
rect 22296 7886 22324 8588
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 22468 8288 22520 8294
rect 22468 8230 22520 8236
rect 22480 7954 22508 8230
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 22572 7886 22600 8434
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 22020 7806 22232 7834
rect 22284 7880 22336 7886
rect 22560 7880 22612 7886
rect 22284 7822 22336 7828
rect 22480 7828 22560 7834
rect 22480 7822 22612 7828
rect 22480 7806 22600 7822
rect 22652 7812 22704 7818
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 20074 6760 20130 6769
rect 20824 6730 20852 7754
rect 22020 7002 22048 7806
rect 22480 7750 22508 7806
rect 22652 7754 22704 7760
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22112 7410 22140 7686
rect 22198 7644 22506 7653
rect 22198 7642 22204 7644
rect 22260 7642 22284 7644
rect 22340 7642 22364 7644
rect 22420 7642 22444 7644
rect 22500 7642 22506 7644
rect 22260 7590 22262 7642
rect 22442 7590 22444 7642
rect 22198 7588 22204 7590
rect 22260 7588 22284 7590
rect 22340 7588 22364 7590
rect 22420 7588 22444 7590
rect 22500 7588 22506 7590
rect 22198 7579 22506 7588
rect 22664 7546 22692 7754
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 22296 7002 22324 7278
rect 22008 6996 22060 7002
rect 22008 6938 22060 6944
rect 22284 6996 22336 7002
rect 22284 6938 22336 6944
rect 22756 6866 22784 10390
rect 23124 10266 23152 13382
rect 23216 10266 23244 13518
rect 23308 13410 23336 14742
rect 23400 14618 23428 14962
rect 23388 14612 23440 14618
rect 23388 14554 23440 14560
rect 23492 13938 23520 17138
rect 23572 16992 23624 16998
rect 23572 16934 23624 16940
rect 23584 15706 23612 16934
rect 23676 16590 23704 17206
rect 23768 16794 23796 17682
rect 24032 17604 24084 17610
rect 24032 17546 24084 17552
rect 23756 16788 23808 16794
rect 23756 16730 23808 16736
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 23940 16584 23992 16590
rect 23940 16526 23992 16532
rect 23756 16516 23808 16522
rect 23756 16458 23808 16464
rect 23664 15972 23716 15978
rect 23664 15914 23716 15920
rect 23572 15700 23624 15706
rect 23572 15642 23624 15648
rect 23584 14618 23612 15642
rect 23572 14612 23624 14618
rect 23572 14554 23624 14560
rect 23676 14414 23704 15914
rect 23768 15570 23796 16458
rect 23952 16114 23980 16526
rect 23940 16108 23992 16114
rect 23940 16050 23992 16056
rect 23756 15564 23808 15570
rect 23756 15506 23808 15512
rect 23952 15502 23980 16050
rect 24044 15570 24072 17546
rect 24032 15564 24084 15570
rect 24032 15506 24084 15512
rect 23940 15496 23992 15502
rect 23940 15438 23992 15444
rect 23952 15042 23980 15438
rect 24044 15094 24072 15506
rect 24124 15428 24176 15434
rect 24124 15370 24176 15376
rect 23768 15014 23980 15042
rect 24032 15088 24084 15094
rect 24032 15030 24084 15036
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 23572 14000 23624 14006
rect 23572 13942 23624 13948
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23308 13382 23428 13410
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 23308 12374 23336 13262
rect 23400 12850 23428 13382
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 23400 12730 23428 12786
rect 23400 12702 23520 12730
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 23296 12368 23348 12374
rect 23296 12310 23348 12316
rect 23400 12306 23428 12582
rect 23388 12300 23440 12306
rect 23388 12242 23440 12248
rect 23296 12232 23348 12238
rect 23492 12186 23520 12702
rect 23296 12174 23348 12180
rect 23308 11898 23336 12174
rect 23400 12158 23520 12186
rect 23296 11892 23348 11898
rect 23296 11834 23348 11840
rect 23296 11756 23348 11762
rect 23296 11698 23348 11704
rect 23308 11150 23336 11698
rect 23296 11144 23348 11150
rect 23296 11086 23348 11092
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 23204 10260 23256 10266
rect 23204 10202 23256 10208
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 22836 9988 22888 9994
rect 22836 9930 22888 9936
rect 22848 9178 22876 9930
rect 23124 9674 23152 9998
rect 23400 9704 23428 12158
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 23492 11014 23520 12038
rect 23584 11082 23612 13942
rect 23768 13326 23796 15014
rect 23940 14884 23992 14890
rect 23940 14826 23992 14832
rect 23952 14482 23980 14826
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23940 14272 23992 14278
rect 23940 14214 23992 14220
rect 23860 14074 23888 14214
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 23768 12170 23796 13262
rect 23756 12164 23808 12170
rect 23756 12106 23808 12112
rect 23848 12096 23900 12102
rect 23848 12038 23900 12044
rect 23664 11688 23716 11694
rect 23664 11630 23716 11636
rect 23676 11218 23704 11630
rect 23664 11212 23716 11218
rect 23664 11154 23716 11160
rect 23572 11076 23624 11082
rect 23572 11018 23624 11024
rect 23480 11008 23532 11014
rect 23480 10950 23532 10956
rect 23676 10606 23704 11154
rect 23860 10810 23888 12038
rect 23952 11642 23980 14214
rect 24136 14006 24164 15370
rect 24124 14000 24176 14006
rect 24124 13942 24176 13948
rect 24136 13870 24164 13942
rect 24124 13864 24176 13870
rect 24124 13806 24176 13812
rect 24124 11824 24176 11830
rect 24124 11766 24176 11772
rect 24032 11756 24084 11762
rect 24032 11698 24084 11704
rect 24044 11642 24072 11698
rect 23952 11614 24072 11642
rect 24136 11558 24164 11766
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24136 11082 24164 11494
rect 24124 11076 24176 11082
rect 24124 11018 24176 11024
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 23032 9646 23152 9674
rect 23308 9676 23428 9704
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 22848 8634 22876 8910
rect 22836 8628 22888 8634
rect 22836 8570 22888 8576
rect 22848 7993 22876 8570
rect 23032 8498 23060 9646
rect 23308 8616 23336 9676
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23400 8906 23428 9522
rect 24032 9104 24084 9110
rect 24032 9046 24084 9052
rect 23388 8900 23440 8906
rect 23388 8842 23440 8848
rect 23308 8588 23428 8616
rect 23020 8492 23072 8498
rect 23020 8434 23072 8440
rect 23296 8492 23348 8498
rect 23296 8434 23348 8440
rect 23112 8424 23164 8430
rect 23112 8366 23164 8372
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 22834 7984 22890 7993
rect 22834 7919 22890 7928
rect 22836 7880 22888 7886
rect 22836 7822 22888 7828
rect 22848 6866 22876 7822
rect 22940 7546 22968 8230
rect 23020 7882 23072 7888
rect 23124 7886 23152 8366
rect 23308 7886 23336 8434
rect 23400 8430 23428 8588
rect 23572 8560 23624 8566
rect 23572 8502 23624 8508
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 23492 8090 23520 8434
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 23020 7824 23072 7830
rect 23112 7880 23164 7886
rect 23296 7880 23348 7886
rect 23032 7546 23060 7824
rect 23112 7822 23164 7828
rect 23216 7840 23296 7868
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 23112 7336 23164 7342
rect 23216 7324 23244 7840
rect 23296 7822 23348 7828
rect 23492 7868 23520 8026
rect 23584 8022 23612 8502
rect 24044 8498 24072 9046
rect 24032 8492 24084 8498
rect 24084 8452 24164 8480
rect 24032 8434 24084 8440
rect 23756 8424 23808 8430
rect 23756 8366 23808 8372
rect 23664 8356 23716 8362
rect 23664 8298 23716 8304
rect 23572 8016 23624 8022
rect 23572 7958 23624 7964
rect 23676 7886 23704 8298
rect 23768 7970 23796 8366
rect 24032 8016 24084 8022
rect 23768 7954 23980 7970
rect 24032 7958 24084 7964
rect 23768 7948 23992 7954
rect 23768 7942 23940 7948
rect 23768 7886 23796 7942
rect 23940 7890 23992 7896
rect 23572 7880 23624 7886
rect 23492 7840 23572 7868
rect 23388 7812 23440 7818
rect 23388 7754 23440 7760
rect 23400 7546 23428 7754
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23492 7478 23520 7840
rect 23572 7822 23624 7828
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 23756 7880 23808 7886
rect 23756 7822 23808 7828
rect 24044 7750 24072 7958
rect 24136 7886 24164 8452
rect 24124 7880 24176 7886
rect 24124 7822 24176 7828
rect 24032 7744 24084 7750
rect 24032 7686 24084 7692
rect 23480 7472 23532 7478
rect 23480 7414 23532 7420
rect 24044 7410 24072 7686
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 23164 7296 23244 7324
rect 23112 7278 23164 7284
rect 24044 6934 24072 7346
rect 24136 7206 24164 7822
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 24136 6934 24164 7142
rect 24032 6928 24084 6934
rect 24032 6870 24084 6876
rect 24124 6928 24176 6934
rect 24124 6870 24176 6876
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 22836 6860 22888 6866
rect 22836 6802 22888 6808
rect 20074 6695 20130 6704
rect 20812 6724 20864 6730
rect 20088 6458 20116 6695
rect 20812 6666 20864 6672
rect 22198 6556 22506 6565
rect 22198 6554 22204 6556
rect 22260 6554 22284 6556
rect 22340 6554 22364 6556
rect 22420 6554 22444 6556
rect 22500 6554 22506 6556
rect 22260 6502 22262 6554
rect 22442 6502 22444 6554
rect 22198 6500 22204 6502
rect 22260 6500 22284 6502
rect 22340 6500 22364 6502
rect 22420 6500 22444 6502
rect 22500 6500 22506 6502
rect 22198 6491 22506 6500
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20258 6352 20314 6361
rect 20258 6287 20260 6296
rect 20312 6287 20314 6296
rect 20260 6258 20312 6264
rect 18657 6012 18965 6021
rect 18657 6010 18663 6012
rect 18719 6010 18743 6012
rect 18799 6010 18823 6012
rect 18879 6010 18903 6012
rect 18959 6010 18965 6012
rect 18719 5958 18721 6010
rect 18901 5958 18903 6010
rect 18657 5956 18663 5958
rect 18719 5956 18743 5958
rect 18799 5956 18823 5958
rect 18879 5956 18903 5958
rect 18959 5956 18965 5958
rect 18657 5947 18965 5956
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 17972 5030 18000 5510
rect 18248 5234 18276 5510
rect 18340 5234 18368 5646
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18524 5234 18552 5510
rect 20272 5370 20300 6258
rect 20548 6186 20576 6394
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18234 5128 18290 5137
rect 18052 5092 18104 5098
rect 18052 5034 18104 5040
rect 18144 5092 18196 5098
rect 18234 5063 18290 5072
rect 18144 5034 18196 5040
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 17880 4826 17908 4966
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 17880 4486 17908 4558
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 17592 3596 17644 3602
rect 17592 3538 17644 3544
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17512 3194 17540 3334
rect 17604 3194 17632 3334
rect 17788 3194 17816 3402
rect 17500 3188 17552 3194
rect 17500 3130 17552 3136
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17132 3052 17184 3058
rect 17420 3046 17540 3074
rect 17132 2994 17184 3000
rect 17144 2854 17172 2994
rect 17512 2990 17540 3046
rect 17972 2990 18000 4966
rect 18064 4622 18092 5034
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 18156 3058 18184 5034
rect 18248 4570 18276 5063
rect 18340 5001 18368 5170
rect 18326 4992 18382 5001
rect 18326 4927 18382 4936
rect 18248 4542 18368 4570
rect 18340 4486 18368 4542
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18248 3058 18276 4422
rect 18524 3942 18552 5170
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 18657 4924 18965 4933
rect 18657 4922 18663 4924
rect 18719 4922 18743 4924
rect 18799 4922 18823 4924
rect 18879 4922 18903 4924
rect 18959 4922 18965 4924
rect 18719 4870 18721 4922
rect 18901 4870 18903 4922
rect 18657 4868 18663 4870
rect 18719 4868 18743 4870
rect 18799 4868 18823 4870
rect 18879 4868 18903 4870
rect 18959 4868 18965 4870
rect 18657 4859 18965 4868
rect 19340 4752 19392 4758
rect 19340 4694 19392 4700
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19260 4146 19288 4558
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18524 3534 18552 3878
rect 18657 3836 18965 3845
rect 18657 3834 18663 3836
rect 18719 3834 18743 3836
rect 18799 3834 18823 3836
rect 18879 3834 18903 3836
rect 18959 3834 18965 3836
rect 18719 3782 18721 3834
rect 18901 3782 18903 3834
rect 18657 3780 18663 3782
rect 18719 3780 18743 3782
rect 18799 3780 18823 3782
rect 18879 3780 18903 3782
rect 18959 3780 18965 3782
rect 18657 3771 18965 3780
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18800 3194 18828 3334
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 17132 2848 17184 2854
rect 17132 2790 17184 2796
rect 13740 2446 13768 2790
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 17512 2378 17540 2926
rect 18657 2748 18965 2757
rect 18657 2746 18663 2748
rect 18719 2746 18743 2748
rect 18799 2746 18823 2748
rect 18879 2746 18903 2748
rect 18959 2746 18965 2748
rect 18719 2694 18721 2746
rect 18901 2694 18903 2746
rect 18657 2692 18663 2694
rect 18719 2692 18743 2694
rect 18799 2692 18823 2694
rect 18879 2692 18903 2694
rect 18959 2692 18965 2694
rect 18657 2683 18965 2692
rect 19352 2446 19380 4694
rect 19536 4690 19564 4966
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19524 4684 19576 4690
rect 19524 4626 19576 4632
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19444 4162 19472 4558
rect 19536 4282 19564 4626
rect 19812 4622 19840 4762
rect 20456 4622 20484 6054
rect 20548 4758 20576 6122
rect 22198 5468 22506 5477
rect 22198 5466 22204 5468
rect 22260 5466 22284 5468
rect 22340 5466 22364 5468
rect 22420 5466 22444 5468
rect 22500 5466 22506 5468
rect 22260 5414 22262 5466
rect 22442 5414 22444 5466
rect 22198 5412 22204 5414
rect 22260 5412 22284 5414
rect 22340 5412 22364 5414
rect 22420 5412 22444 5414
rect 22500 5412 22506 5414
rect 22198 5403 22506 5412
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20536 4752 20588 4758
rect 20536 4694 20588 4700
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 19444 4146 19656 4162
rect 19812 4146 19840 4558
rect 19432 4140 19656 4146
rect 19484 4134 19656 4140
rect 19432 4082 19484 4088
rect 19628 4078 19656 4134
rect 19800 4140 19852 4146
rect 19800 4082 19852 4088
rect 19524 4072 19576 4078
rect 19524 4014 19576 4020
rect 19616 4072 19668 4078
rect 19616 4014 19668 4020
rect 19536 3738 19564 4014
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19812 2854 19840 4082
rect 20180 3942 20208 4558
rect 20456 4282 20484 4558
rect 20548 4282 20576 4694
rect 20732 4622 20760 4966
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 22198 4380 22506 4389
rect 22198 4378 22204 4380
rect 22260 4378 22284 4380
rect 22340 4378 22364 4380
rect 22420 4378 22444 4380
rect 22500 4378 22506 4380
rect 22260 4326 22262 4378
rect 22442 4326 22444 4378
rect 22198 4324 22204 4326
rect 22260 4324 22284 4326
rect 22340 4324 22364 4326
rect 22420 4324 22444 4326
rect 22500 4324 22506 4326
rect 22198 4315 22506 4324
rect 20444 4276 20496 4282
rect 20444 4218 20496 4224
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 24228 4049 24256 20998
rect 24320 19334 24348 22102
rect 24504 22030 24532 23054
rect 24676 23044 24728 23050
rect 24676 22986 24728 22992
rect 24584 22636 24636 22642
rect 24584 22578 24636 22584
rect 24492 22024 24544 22030
rect 24492 21966 24544 21972
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24412 21554 24440 21830
rect 24400 21548 24452 21554
rect 24400 21490 24452 21496
rect 24596 21350 24624 22578
rect 24688 22234 24716 22986
rect 24768 22976 24820 22982
rect 24768 22918 24820 22924
rect 24952 22976 25004 22982
rect 24952 22918 25004 22924
rect 24780 22234 24808 22918
rect 24964 22710 24992 22918
rect 24952 22704 25004 22710
rect 24952 22646 25004 22652
rect 25056 22642 25084 23122
rect 25332 22778 25360 30194
rect 28540 30048 28592 30054
rect 28540 29990 28592 29996
rect 25740 29948 26048 29957
rect 25740 29946 25746 29948
rect 25802 29946 25826 29948
rect 25882 29946 25906 29948
rect 25962 29946 25986 29948
rect 26042 29946 26048 29948
rect 25802 29894 25804 29946
rect 25984 29894 25986 29946
rect 25740 29892 25746 29894
rect 25802 29892 25826 29894
rect 25882 29892 25906 29894
rect 25962 29892 25986 29894
rect 26042 29892 26048 29894
rect 25740 29883 26048 29892
rect 28552 29306 28580 29990
rect 28540 29300 28592 29306
rect 28540 29242 28592 29248
rect 28736 29073 28764 30194
rect 28920 30190 28948 30631
rect 29012 30326 29040 31925
rect 29281 30492 29589 30501
rect 29281 30490 29287 30492
rect 29343 30490 29367 30492
rect 29423 30490 29447 30492
rect 29503 30490 29527 30492
rect 29583 30490 29589 30492
rect 29343 30438 29345 30490
rect 29525 30438 29527 30490
rect 29281 30436 29287 30438
rect 29343 30436 29367 30438
rect 29423 30436 29447 30438
rect 29503 30436 29527 30438
rect 29583 30436 29589 30438
rect 29281 30427 29589 30436
rect 29000 30320 29052 30326
rect 29000 30262 29052 30268
rect 28908 30184 28960 30190
rect 28908 30126 28960 30132
rect 29281 29404 29589 29413
rect 29281 29402 29287 29404
rect 29343 29402 29367 29404
rect 29423 29402 29447 29404
rect 29503 29402 29527 29404
rect 29583 29402 29589 29404
rect 29343 29350 29345 29402
rect 29525 29350 29527 29402
rect 29281 29348 29287 29350
rect 29343 29348 29367 29350
rect 29423 29348 29447 29350
rect 29503 29348 29527 29350
rect 29583 29348 29589 29350
rect 29281 29339 29589 29348
rect 28722 29064 28778 29073
rect 28722 28999 28778 29008
rect 25740 28860 26048 28869
rect 25740 28858 25746 28860
rect 25802 28858 25826 28860
rect 25882 28858 25906 28860
rect 25962 28858 25986 28860
rect 26042 28858 26048 28860
rect 25802 28806 25804 28858
rect 25984 28806 25986 28858
rect 25740 28804 25746 28806
rect 25802 28804 25826 28806
rect 25882 28804 25906 28806
rect 25962 28804 25986 28806
rect 26042 28804 26048 28806
rect 25740 28795 26048 28804
rect 29281 28316 29589 28325
rect 29281 28314 29287 28316
rect 29343 28314 29367 28316
rect 29423 28314 29447 28316
rect 29503 28314 29527 28316
rect 29583 28314 29589 28316
rect 29343 28262 29345 28314
rect 29525 28262 29527 28314
rect 29281 28260 29287 28262
rect 29343 28260 29367 28262
rect 29423 28260 29447 28262
rect 29503 28260 29527 28262
rect 29583 28260 29589 28262
rect 29281 28251 29589 28260
rect 25740 27772 26048 27781
rect 25740 27770 25746 27772
rect 25802 27770 25826 27772
rect 25882 27770 25906 27772
rect 25962 27770 25986 27772
rect 26042 27770 26048 27772
rect 25802 27718 25804 27770
rect 25984 27718 25986 27770
rect 25740 27716 25746 27718
rect 25802 27716 25826 27718
rect 25882 27716 25906 27718
rect 25962 27716 25986 27718
rect 26042 27716 26048 27718
rect 25740 27707 26048 27716
rect 29281 27228 29589 27237
rect 29281 27226 29287 27228
rect 29343 27226 29367 27228
rect 29423 27226 29447 27228
rect 29503 27226 29527 27228
rect 29583 27226 29589 27228
rect 29343 27174 29345 27226
rect 29525 27174 29527 27226
rect 29281 27172 29287 27174
rect 29343 27172 29367 27174
rect 29423 27172 29447 27174
rect 29503 27172 29527 27174
rect 29583 27172 29589 27174
rect 29281 27163 29589 27172
rect 28264 26988 28316 26994
rect 28264 26930 28316 26936
rect 25740 26684 26048 26693
rect 25740 26682 25746 26684
rect 25802 26682 25826 26684
rect 25882 26682 25906 26684
rect 25962 26682 25986 26684
rect 26042 26682 26048 26684
rect 25802 26630 25804 26682
rect 25984 26630 25986 26682
rect 25740 26628 25746 26630
rect 25802 26628 25826 26630
rect 25882 26628 25906 26630
rect 25962 26628 25986 26630
rect 26042 26628 26048 26630
rect 25740 26619 26048 26628
rect 25740 25596 26048 25605
rect 25740 25594 25746 25596
rect 25802 25594 25826 25596
rect 25882 25594 25906 25596
rect 25962 25594 25986 25596
rect 26042 25594 26048 25596
rect 25802 25542 25804 25594
rect 25984 25542 25986 25594
rect 25740 25540 25746 25542
rect 25802 25540 25826 25542
rect 25882 25540 25906 25542
rect 25962 25540 25986 25542
rect 26042 25540 26048 25542
rect 25740 25531 26048 25540
rect 25740 24508 26048 24517
rect 25740 24506 25746 24508
rect 25802 24506 25826 24508
rect 25882 24506 25906 24508
rect 25962 24506 25986 24508
rect 26042 24506 26048 24508
rect 25802 24454 25804 24506
rect 25984 24454 25986 24506
rect 25740 24452 25746 24454
rect 25802 24452 25826 24454
rect 25882 24452 25906 24454
rect 25962 24452 25986 24454
rect 26042 24452 26048 24454
rect 25740 24443 26048 24452
rect 25740 23420 26048 23429
rect 25740 23418 25746 23420
rect 25802 23418 25826 23420
rect 25882 23418 25906 23420
rect 25962 23418 25986 23420
rect 26042 23418 26048 23420
rect 25802 23366 25804 23418
rect 25984 23366 25986 23418
rect 25740 23364 25746 23366
rect 25802 23364 25826 23366
rect 25882 23364 25906 23366
rect 25962 23364 25986 23366
rect 26042 23364 26048 23366
rect 25740 23355 26048 23364
rect 25504 23044 25556 23050
rect 25504 22986 25556 22992
rect 25320 22772 25372 22778
rect 25320 22714 25372 22720
rect 24860 22636 24912 22642
rect 24860 22578 24912 22584
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 24676 22228 24728 22234
rect 24676 22170 24728 22176
rect 24768 22228 24820 22234
rect 24768 22170 24820 22176
rect 24674 22128 24730 22137
rect 24674 22063 24730 22072
rect 24688 22030 24716 22063
rect 24676 22024 24728 22030
rect 24676 21966 24728 21972
rect 24872 21622 24900 22578
rect 24952 22500 25004 22506
rect 24952 22442 25004 22448
rect 24860 21616 24912 21622
rect 24860 21558 24912 21564
rect 24964 21554 24992 22442
rect 25056 22030 25084 22578
rect 25240 22098 25268 22578
rect 25228 22092 25280 22098
rect 25228 22034 25280 22040
rect 25516 22030 25544 22986
rect 25596 22568 25648 22574
rect 25596 22510 25648 22516
rect 25608 22216 25636 22510
rect 25740 22332 26048 22341
rect 25740 22330 25746 22332
rect 25802 22330 25826 22332
rect 25882 22330 25906 22332
rect 25962 22330 25986 22332
rect 26042 22330 26048 22332
rect 25802 22278 25804 22330
rect 25984 22278 25986 22330
rect 25740 22276 25746 22278
rect 25802 22276 25826 22278
rect 25882 22276 25906 22278
rect 25962 22276 25986 22278
rect 26042 22276 26048 22278
rect 25740 22267 26048 22276
rect 25608 22188 25728 22216
rect 25044 22024 25096 22030
rect 25044 21966 25096 21972
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 25504 22024 25556 22030
rect 25504 21966 25556 21972
rect 25148 21622 25176 21966
rect 25136 21616 25188 21622
rect 25136 21558 25188 21564
rect 25318 21584 25374 21593
rect 24676 21548 24728 21554
rect 24676 21490 24728 21496
rect 24952 21548 25004 21554
rect 25516 21554 25544 21966
rect 25700 21894 25728 22188
rect 26146 21992 26202 22001
rect 26146 21927 26202 21936
rect 25596 21888 25648 21894
rect 25596 21830 25648 21836
rect 25688 21888 25740 21894
rect 25688 21830 25740 21836
rect 25318 21519 25320 21528
rect 24952 21490 25004 21496
rect 25372 21519 25374 21528
rect 25504 21548 25556 21554
rect 25320 21490 25372 21496
rect 25504 21490 25556 21496
rect 24584 21344 24636 21350
rect 24584 21286 24636 21292
rect 24688 20602 24716 21490
rect 25608 21185 25636 21830
rect 25740 21244 26048 21253
rect 25740 21242 25746 21244
rect 25802 21242 25826 21244
rect 25882 21242 25906 21244
rect 25962 21242 25986 21244
rect 26042 21242 26048 21244
rect 25802 21190 25804 21242
rect 25984 21190 25986 21242
rect 25740 21188 25746 21190
rect 25802 21188 25826 21190
rect 25882 21188 25906 21190
rect 25962 21188 25986 21190
rect 26042 21188 26048 21190
rect 25594 21176 25650 21185
rect 25740 21179 26048 21188
rect 26160 21146 26188 21927
rect 26976 21548 27028 21554
rect 26976 21490 27028 21496
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 27804 21548 27856 21554
rect 27804 21490 27856 21496
rect 26240 21412 26292 21418
rect 26240 21354 26292 21360
rect 25594 21111 25650 21120
rect 26148 21140 26200 21146
rect 25608 21010 25636 21111
rect 26148 21082 26200 21088
rect 25596 21004 25648 21010
rect 25596 20946 25648 20952
rect 26252 20942 26280 21354
rect 26988 21146 27016 21490
rect 27066 21448 27122 21457
rect 27066 21383 27068 21392
rect 27120 21383 27122 21392
rect 27068 21354 27120 21360
rect 27252 21344 27304 21350
rect 27252 21286 27304 21292
rect 26976 21140 27028 21146
rect 26976 21082 27028 21088
rect 27068 21004 27120 21010
rect 27068 20946 27120 20952
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 26608 20936 26660 20942
rect 26608 20878 26660 20884
rect 25320 20868 25372 20874
rect 25320 20810 25372 20816
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 25332 20466 25360 20810
rect 26620 20466 26648 20878
rect 27080 20602 27108 20946
rect 27068 20596 27120 20602
rect 27068 20538 27120 20544
rect 25320 20460 25372 20466
rect 25320 20402 25372 20408
rect 26608 20460 26660 20466
rect 26608 20402 26660 20408
rect 24320 19306 24440 19334
rect 24412 12434 24440 19306
rect 24492 18624 24544 18630
rect 24492 18566 24544 18572
rect 24504 18358 24532 18566
rect 25332 18426 25360 20402
rect 27264 20330 27292 21286
rect 27540 21010 27568 21490
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 27528 21004 27580 21010
rect 27356 20964 27528 20992
rect 27356 20466 27384 20964
rect 27528 20946 27580 20952
rect 27436 20800 27488 20806
rect 27436 20742 27488 20748
rect 27448 20466 27476 20742
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 27436 20460 27488 20466
rect 27436 20402 27488 20408
rect 27252 20324 27304 20330
rect 27252 20266 27304 20272
rect 25740 20156 26048 20165
rect 25740 20154 25746 20156
rect 25802 20154 25826 20156
rect 25882 20154 25906 20156
rect 25962 20154 25986 20156
rect 26042 20154 26048 20156
rect 25802 20102 25804 20154
rect 25984 20102 25986 20154
rect 25740 20100 25746 20102
rect 25802 20100 25826 20102
rect 25882 20100 25906 20102
rect 25962 20100 25986 20102
rect 26042 20100 26048 20102
rect 25740 20091 26048 20100
rect 27264 19854 27292 20266
rect 27356 20262 27384 20402
rect 27344 20256 27396 20262
rect 27344 20198 27396 20204
rect 27356 19854 27384 20198
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 27344 19848 27396 19854
rect 27344 19790 27396 19796
rect 26976 19712 27028 19718
rect 26976 19654 27028 19660
rect 27068 19712 27120 19718
rect 27068 19654 27120 19660
rect 25740 19068 26048 19077
rect 25740 19066 25746 19068
rect 25802 19066 25826 19068
rect 25882 19066 25906 19068
rect 25962 19066 25986 19068
rect 26042 19066 26048 19068
rect 25802 19014 25804 19066
rect 25984 19014 25986 19066
rect 25740 19012 25746 19014
rect 25802 19012 25826 19014
rect 25882 19012 25906 19014
rect 25962 19012 25986 19014
rect 26042 19012 26048 19014
rect 25740 19003 26048 19012
rect 25320 18420 25372 18426
rect 25320 18362 25372 18368
rect 24492 18352 24544 18358
rect 24492 18294 24544 18300
rect 24952 18352 25004 18358
rect 24952 18294 25004 18300
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 24872 17746 24900 18022
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24780 17202 24808 17614
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 24768 17196 24820 17202
rect 24768 17138 24820 17144
rect 24872 16998 24900 17478
rect 24964 17134 24992 18294
rect 25504 18216 25556 18222
rect 25504 18158 25556 18164
rect 26884 18216 26936 18222
rect 26884 18158 26936 18164
rect 25228 18148 25280 18154
rect 25228 18090 25280 18096
rect 25240 17898 25268 18090
rect 25148 17882 25268 17898
rect 25136 17876 25268 17882
rect 25188 17870 25268 17876
rect 25136 17818 25188 17824
rect 25136 17672 25188 17678
rect 25136 17614 25188 17620
rect 25148 17338 25176 17614
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25240 17202 25268 17870
rect 25516 17814 25544 18158
rect 26424 18148 26476 18154
rect 26424 18090 26476 18096
rect 25740 17980 26048 17989
rect 25740 17978 25746 17980
rect 25802 17978 25826 17980
rect 25882 17978 25906 17980
rect 25962 17978 25986 17980
rect 26042 17978 26048 17980
rect 25802 17926 25804 17978
rect 25984 17926 25986 17978
rect 25740 17924 25746 17926
rect 25802 17924 25826 17926
rect 25882 17924 25906 17926
rect 25962 17924 25986 17926
rect 26042 17924 26048 17926
rect 25740 17915 26048 17924
rect 25872 17876 25924 17882
rect 25872 17818 25924 17824
rect 25504 17808 25556 17814
rect 25504 17750 25556 17756
rect 25320 17672 25372 17678
rect 25320 17614 25372 17620
rect 25228 17196 25280 17202
rect 25228 17138 25280 17144
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 24860 16992 24912 16998
rect 24860 16934 24912 16940
rect 24676 16584 24728 16590
rect 24676 16526 24728 16532
rect 24688 15570 24716 16526
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24872 15162 24900 16934
rect 25332 16794 25360 17614
rect 25412 17604 25464 17610
rect 25412 17546 25464 17552
rect 25424 17338 25452 17546
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 25516 17270 25544 17750
rect 25884 17678 25912 17818
rect 26240 17808 26292 17814
rect 26146 17776 26202 17785
rect 26202 17756 26240 17762
rect 26202 17750 26292 17756
rect 26202 17734 26280 17750
rect 26436 17746 26464 18090
rect 26792 17876 26844 17882
rect 26792 17818 26844 17824
rect 26700 17808 26752 17814
rect 26700 17750 26752 17756
rect 26146 17711 26202 17720
rect 25872 17672 25924 17678
rect 25872 17614 25924 17620
rect 25964 17672 26016 17678
rect 25964 17614 26016 17620
rect 25504 17264 25556 17270
rect 25504 17206 25556 17212
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25320 16788 25372 16794
rect 25320 16730 25372 16736
rect 25424 16572 25452 17138
rect 25516 16674 25544 17206
rect 25884 17066 25912 17614
rect 25976 17134 26004 17614
rect 26252 17542 26280 17734
rect 26424 17740 26476 17746
rect 26424 17682 26476 17688
rect 26516 17740 26568 17746
rect 26516 17682 26568 17688
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 26240 17536 26292 17542
rect 26240 17478 26292 17484
rect 26424 17536 26476 17542
rect 26424 17478 26476 17484
rect 26054 17232 26110 17241
rect 26054 17167 26056 17176
rect 26108 17167 26110 17176
rect 26056 17138 26108 17144
rect 25964 17128 26016 17134
rect 25964 17070 26016 17076
rect 25872 17060 25924 17066
rect 25872 17002 25924 17008
rect 25740 16892 26048 16901
rect 25740 16890 25746 16892
rect 25802 16890 25826 16892
rect 25882 16890 25906 16892
rect 25962 16890 25986 16892
rect 26042 16890 26048 16892
rect 25802 16838 25804 16890
rect 25984 16838 25986 16890
rect 25740 16836 25746 16838
rect 25802 16836 25826 16838
rect 25882 16836 25906 16838
rect 25962 16836 25986 16838
rect 26042 16836 26048 16838
rect 25740 16827 26048 16836
rect 25516 16658 25636 16674
rect 25516 16652 25648 16658
rect 25516 16646 25596 16652
rect 25596 16594 25648 16600
rect 26160 16590 26188 17478
rect 26240 17332 26292 17338
rect 26240 17274 26292 17280
rect 25504 16584 25556 16590
rect 25424 16544 25504 16572
rect 25504 16526 25556 16532
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 25516 16046 25544 16526
rect 26056 16448 26108 16454
rect 26054 16416 26056 16425
rect 26108 16416 26110 16425
rect 26054 16351 26110 16360
rect 25504 16040 25556 16046
rect 25504 15982 25556 15988
rect 25134 15464 25190 15473
rect 25056 15422 25134 15450
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24860 15156 24912 15162
rect 24860 15098 24912 15104
rect 24780 15026 24808 15098
rect 24676 15020 24728 15026
rect 24676 14962 24728 14968
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24688 14906 24716 14962
rect 25056 14906 25084 15422
rect 25134 15399 25190 15408
rect 25516 14958 25544 15982
rect 26148 15904 26200 15910
rect 26148 15846 26200 15852
rect 25740 15804 26048 15813
rect 25740 15802 25746 15804
rect 25802 15802 25826 15804
rect 25882 15802 25906 15804
rect 25962 15802 25986 15804
rect 26042 15802 26048 15804
rect 25802 15750 25804 15802
rect 25984 15750 25986 15802
rect 25740 15748 25746 15750
rect 25802 15748 25826 15750
rect 25882 15748 25906 15750
rect 25962 15748 25986 15750
rect 26042 15748 26048 15750
rect 25740 15739 26048 15748
rect 26160 15706 26188 15846
rect 26148 15700 26200 15706
rect 26148 15642 26200 15648
rect 26252 15570 26280 17274
rect 26436 16998 26464 17478
rect 26528 16998 26556 17682
rect 26608 17672 26660 17678
rect 26712 17649 26740 17750
rect 26608 17614 26660 17620
rect 26698 17640 26754 17649
rect 26620 17338 26648 17614
rect 26804 17610 26832 17818
rect 26698 17575 26754 17584
rect 26792 17604 26844 17610
rect 26608 17332 26660 17338
rect 26608 17274 26660 17280
rect 26712 17134 26740 17575
rect 26792 17546 26844 17552
rect 26700 17128 26752 17134
rect 26700 17070 26752 17076
rect 26424 16992 26476 16998
rect 26424 16934 26476 16940
rect 26516 16992 26568 16998
rect 26516 16934 26568 16940
rect 26436 16726 26464 16934
rect 26792 16788 26844 16794
rect 26792 16730 26844 16736
rect 26424 16720 26476 16726
rect 26424 16662 26476 16668
rect 26436 16454 26464 16662
rect 26700 16516 26752 16522
rect 26700 16458 26752 16464
rect 26424 16448 26476 16454
rect 26424 16390 26476 16396
rect 26608 16448 26660 16454
rect 26608 16390 26660 16396
rect 26620 16114 26648 16390
rect 26712 16250 26740 16458
rect 26700 16244 26752 16250
rect 26700 16186 26752 16192
rect 26608 16108 26660 16114
rect 26608 16050 26660 16056
rect 26804 15638 26832 16730
rect 26516 15632 26568 15638
rect 26516 15574 26568 15580
rect 26792 15632 26844 15638
rect 26792 15574 26844 15580
rect 26240 15564 26292 15570
rect 26240 15506 26292 15512
rect 26528 15473 26556 15574
rect 26514 15464 26570 15473
rect 26514 15399 26570 15408
rect 26148 15360 26200 15366
rect 26148 15302 26200 15308
rect 26516 15360 26568 15366
rect 26516 15302 26568 15308
rect 26160 15178 26188 15302
rect 26528 15178 26556 15302
rect 26160 15150 26556 15178
rect 24688 14878 25084 14906
rect 25504 14952 25556 14958
rect 25504 14894 25556 14900
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24504 14618 24532 14758
rect 24492 14612 24544 14618
rect 24492 14554 24544 14560
rect 24492 14476 24544 14482
rect 24492 14418 24544 14424
rect 24504 13938 24532 14418
rect 25516 14278 25544 14894
rect 25740 14716 26048 14725
rect 25740 14714 25746 14716
rect 25802 14714 25826 14716
rect 25882 14714 25906 14716
rect 25962 14714 25986 14716
rect 26042 14714 26048 14716
rect 25802 14662 25804 14714
rect 25984 14662 25986 14714
rect 25740 14660 25746 14662
rect 25802 14660 25826 14662
rect 25882 14660 25906 14662
rect 25962 14660 25986 14662
rect 26042 14660 26048 14662
rect 25740 14651 26048 14660
rect 26896 14618 26924 18158
rect 26988 17814 27016 19654
rect 26976 17808 27028 17814
rect 26976 17750 27028 17756
rect 26976 17128 27028 17134
rect 26976 17070 27028 17076
rect 26988 16794 27016 17070
rect 26976 16788 27028 16794
rect 26976 16730 27028 16736
rect 26988 15706 27016 16730
rect 26976 15700 27028 15706
rect 26976 15642 27028 15648
rect 27080 14906 27108 19654
rect 27448 19378 27476 20402
rect 27528 20256 27580 20262
rect 27528 20198 27580 20204
rect 27540 19854 27568 20198
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 27632 19718 27660 21286
rect 27816 21010 27844 21490
rect 27988 21072 28040 21078
rect 27988 21014 28040 21020
rect 27804 21004 27856 21010
rect 27804 20946 27856 20952
rect 28000 20874 28028 21014
rect 27988 20868 28040 20874
rect 27988 20810 28040 20816
rect 27712 20256 27764 20262
rect 27712 20198 27764 20204
rect 27620 19712 27672 19718
rect 27620 19654 27672 19660
rect 27436 19372 27488 19378
rect 27436 19314 27488 19320
rect 27724 18766 27752 20198
rect 28000 19854 28028 20810
rect 28172 20800 28224 20806
rect 28172 20742 28224 20748
rect 28080 20460 28132 20466
rect 28080 20402 28132 20408
rect 28092 20058 28120 20402
rect 28080 20052 28132 20058
rect 28080 19994 28132 20000
rect 27988 19848 28040 19854
rect 27988 19790 28040 19796
rect 28092 19514 28120 19994
rect 28184 19854 28212 20742
rect 28172 19848 28224 19854
rect 28172 19790 28224 19796
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 27804 19304 27856 19310
rect 27804 19246 27856 19252
rect 27712 18760 27764 18766
rect 27712 18702 27764 18708
rect 27252 18216 27304 18222
rect 27252 18158 27304 18164
rect 27264 17882 27292 18158
rect 27252 17876 27304 17882
rect 27252 17818 27304 17824
rect 27160 17672 27212 17678
rect 27160 17614 27212 17620
rect 27526 17640 27582 17649
rect 27172 17066 27200 17614
rect 27526 17575 27528 17584
rect 27580 17575 27582 17584
rect 27528 17546 27580 17552
rect 27540 17270 27568 17546
rect 27712 17536 27764 17542
rect 27632 17484 27712 17490
rect 27632 17478 27764 17484
rect 27632 17462 27752 17478
rect 27528 17264 27580 17270
rect 27250 17232 27306 17241
rect 27528 17206 27580 17212
rect 27306 17176 27384 17184
rect 27250 17167 27252 17176
rect 27304 17156 27384 17176
rect 27252 17138 27304 17144
rect 27160 17060 27212 17066
rect 27160 17002 27212 17008
rect 27252 16448 27304 16454
rect 27252 16390 27304 16396
rect 27264 15502 27292 16390
rect 27356 16250 27384 17156
rect 27528 17128 27580 17134
rect 27528 17070 27580 17076
rect 27540 16794 27568 17070
rect 27528 16788 27580 16794
rect 27528 16730 27580 16736
rect 27632 16590 27660 17462
rect 27816 17354 27844 19246
rect 27896 17808 27948 17814
rect 27896 17750 27948 17756
rect 27724 17326 27844 17354
rect 27724 17241 27752 17326
rect 27710 17232 27766 17241
rect 27908 17202 27936 17750
rect 27988 17536 28040 17542
rect 27988 17478 28040 17484
rect 28080 17536 28132 17542
rect 28080 17478 28132 17484
rect 27710 17167 27766 17176
rect 27804 17196 27856 17202
rect 27804 17138 27856 17144
rect 27896 17196 27948 17202
rect 27896 17138 27948 17144
rect 27816 16794 27844 17138
rect 28000 16998 28028 17478
rect 27988 16992 28040 16998
rect 27988 16934 28040 16940
rect 27804 16788 27856 16794
rect 27804 16730 27856 16736
rect 27896 16788 27948 16794
rect 27896 16730 27948 16736
rect 27908 16590 27936 16730
rect 28092 16674 28120 17478
rect 28000 16658 28120 16674
rect 27988 16652 28120 16658
rect 28040 16646 28120 16652
rect 27988 16594 28040 16600
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27896 16584 27948 16590
rect 27896 16526 27948 16532
rect 27988 16448 28040 16454
rect 27986 16416 27988 16425
rect 28040 16416 28042 16425
rect 27986 16351 28042 16360
rect 27344 16244 27396 16250
rect 27344 16186 27396 16192
rect 27804 16244 27856 16250
rect 27804 16186 27856 16192
rect 27344 15700 27396 15706
rect 27344 15642 27396 15648
rect 27252 15496 27304 15502
rect 27252 15438 27304 15444
rect 27160 15360 27212 15366
rect 27160 15302 27212 15308
rect 27252 15360 27304 15366
rect 27252 15302 27304 15308
rect 27172 15162 27200 15302
rect 27160 15156 27212 15162
rect 27160 15098 27212 15104
rect 27160 15020 27212 15026
rect 27264 15008 27292 15302
rect 27356 15162 27384 15642
rect 27712 15564 27764 15570
rect 27712 15506 27764 15512
rect 27344 15156 27396 15162
rect 27344 15098 27396 15104
rect 27212 14980 27292 15008
rect 27160 14962 27212 14968
rect 27080 14878 27200 14906
rect 27724 14890 27752 15506
rect 27816 15094 27844 16186
rect 28172 15632 28224 15638
rect 28172 15574 28224 15580
rect 27804 15088 27856 15094
rect 27804 15030 27856 15036
rect 28184 15026 28212 15574
rect 28172 15020 28224 15026
rect 28172 14962 28224 14968
rect 27068 14816 27120 14822
rect 27068 14758 27120 14764
rect 26884 14612 26936 14618
rect 26884 14554 26936 14560
rect 27080 14482 27108 14758
rect 27068 14476 27120 14482
rect 27068 14418 27120 14424
rect 25872 14408 25924 14414
rect 25872 14350 25924 14356
rect 25504 14272 25556 14278
rect 25504 14214 25556 14220
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 24492 13932 24544 13938
rect 24492 13874 24544 13880
rect 25148 13394 25176 14010
rect 25884 13938 25912 14350
rect 25872 13932 25924 13938
rect 25872 13874 25924 13880
rect 26332 13864 26384 13870
rect 26332 13806 26384 13812
rect 25320 13728 25372 13734
rect 25320 13670 25372 13676
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 25332 13530 25360 13670
rect 25740 13628 26048 13637
rect 25740 13626 25746 13628
rect 25802 13626 25826 13628
rect 25882 13626 25906 13628
rect 25962 13626 25986 13628
rect 26042 13626 26048 13628
rect 25802 13574 25804 13626
rect 25984 13574 25986 13626
rect 25740 13572 25746 13574
rect 25802 13572 25826 13574
rect 25882 13572 25906 13574
rect 25962 13572 25986 13574
rect 26042 13572 26048 13574
rect 25740 13563 26048 13572
rect 25320 13524 25372 13530
rect 25320 13466 25372 13472
rect 26252 13394 26280 13670
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 26240 13388 26292 13394
rect 26240 13330 26292 13336
rect 25740 12540 26048 12549
rect 25740 12538 25746 12540
rect 25802 12538 25826 12540
rect 25882 12538 25906 12540
rect 25962 12538 25986 12540
rect 26042 12538 26048 12540
rect 25802 12486 25804 12538
rect 25984 12486 25986 12538
rect 25740 12484 25746 12486
rect 25802 12484 25826 12486
rect 25882 12484 25906 12486
rect 25962 12484 25986 12486
rect 26042 12484 26048 12486
rect 25740 12475 26048 12484
rect 24412 12406 24532 12434
rect 24308 12096 24360 12102
rect 24308 12038 24360 12044
rect 24320 11694 24348 12038
rect 24308 11688 24360 11694
rect 24308 11630 24360 11636
rect 24400 11212 24452 11218
rect 24400 11154 24452 11160
rect 24412 11121 24440 11154
rect 24398 11112 24454 11121
rect 24398 11047 24454 11056
rect 24412 10742 24440 11047
rect 24400 10736 24452 10742
rect 24400 10678 24452 10684
rect 24308 8832 24360 8838
rect 24308 8774 24360 8780
rect 24320 7818 24348 8774
rect 24308 7812 24360 7818
rect 24308 7754 24360 7760
rect 24320 7410 24348 7754
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 24320 6798 24348 7346
rect 24400 7200 24452 7206
rect 24400 7142 24452 7148
rect 24412 7002 24440 7142
rect 24400 6996 24452 7002
rect 24400 6938 24452 6944
rect 24308 6792 24360 6798
rect 24308 6734 24360 6740
rect 24306 5536 24362 5545
rect 24306 5471 24362 5480
rect 24320 4214 24348 5471
rect 24308 4208 24360 4214
rect 24308 4150 24360 4156
rect 24504 4146 24532 12406
rect 25596 11552 25648 11558
rect 25596 11494 25648 11500
rect 26240 11552 26292 11558
rect 26240 11494 26292 11500
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 24768 11076 24820 11082
rect 24768 11018 24820 11024
rect 24780 10538 24808 11018
rect 24768 10532 24820 10538
rect 24768 10474 24820 10480
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24596 7886 24624 8366
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 24688 7886 24716 8230
rect 24584 7880 24636 7886
rect 24584 7822 24636 7828
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24688 7562 24716 7822
rect 24596 7534 24716 7562
rect 24596 7478 24624 7534
rect 24584 7472 24636 7478
rect 24584 7414 24636 7420
rect 24780 6798 24808 10474
rect 24964 10470 24992 11086
rect 25228 11076 25280 11082
rect 25608 11054 25636 11494
rect 25740 11452 26048 11461
rect 25740 11450 25746 11452
rect 25802 11450 25826 11452
rect 25882 11450 25906 11452
rect 25962 11450 25986 11452
rect 26042 11450 26048 11452
rect 25802 11398 25804 11450
rect 25984 11398 25986 11450
rect 25740 11396 25746 11398
rect 25802 11396 25826 11398
rect 25882 11396 25906 11398
rect 25962 11396 25986 11398
rect 26042 11396 26048 11398
rect 25740 11387 26048 11396
rect 25608 11026 25912 11054
rect 25228 11018 25280 11024
rect 25240 10810 25268 11018
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25884 10606 25912 11026
rect 26056 11008 26108 11014
rect 26056 10950 26108 10956
rect 26068 10742 26096 10950
rect 26252 10742 26280 11494
rect 26344 11150 26372 13806
rect 26700 11620 26752 11626
rect 26700 11562 26752 11568
rect 26712 11354 26740 11562
rect 26700 11348 26752 11354
rect 26700 11290 26752 11296
rect 26332 11144 26384 11150
rect 26332 11086 26384 11092
rect 27068 11144 27120 11150
rect 27068 11086 27120 11092
rect 26056 10736 26108 10742
rect 26056 10678 26108 10684
rect 26240 10736 26292 10742
rect 26240 10678 26292 10684
rect 25596 10600 25648 10606
rect 25596 10542 25648 10548
rect 25872 10600 25924 10606
rect 25872 10542 25924 10548
rect 26148 10600 26200 10606
rect 26148 10542 26200 10548
rect 24952 10464 25004 10470
rect 24952 10406 25004 10412
rect 24964 8974 24992 10406
rect 25608 10266 25636 10542
rect 25740 10364 26048 10373
rect 25740 10362 25746 10364
rect 25802 10362 25826 10364
rect 25882 10362 25906 10364
rect 25962 10362 25986 10364
rect 26042 10362 26048 10364
rect 25802 10310 25804 10362
rect 25984 10310 25986 10362
rect 25740 10308 25746 10310
rect 25802 10308 25826 10310
rect 25882 10308 25906 10310
rect 25962 10308 25986 10310
rect 26042 10308 26048 10310
rect 25740 10299 26048 10308
rect 25596 10260 25648 10266
rect 25596 10202 25648 10208
rect 26160 9874 26188 10542
rect 26252 9994 26280 10678
rect 26424 10668 26476 10674
rect 26424 10610 26476 10616
rect 26516 10668 26568 10674
rect 26516 10610 26568 10616
rect 26436 10062 26464 10610
rect 26424 10056 26476 10062
rect 26424 9998 26476 10004
rect 26240 9988 26292 9994
rect 26240 9930 26292 9936
rect 26160 9846 26280 9874
rect 25596 9648 25648 9654
rect 25596 9590 25648 9596
rect 25504 9580 25556 9586
rect 25504 9522 25556 9528
rect 24952 8968 25004 8974
rect 24952 8910 25004 8916
rect 24964 7410 24992 8910
rect 25516 8498 25544 9522
rect 25608 8974 25636 9590
rect 26148 9444 26200 9450
rect 26148 9386 26200 9392
rect 25740 9276 26048 9285
rect 25740 9274 25746 9276
rect 25802 9274 25826 9276
rect 25882 9274 25906 9276
rect 25962 9274 25986 9276
rect 26042 9274 26048 9276
rect 25802 9222 25804 9274
rect 25984 9222 25986 9274
rect 25740 9220 25746 9222
rect 25802 9220 25826 9222
rect 25882 9220 25906 9222
rect 25962 9220 25986 9222
rect 26042 9220 26048 9222
rect 25740 9211 26048 9220
rect 26160 8974 26188 9386
rect 25596 8968 25648 8974
rect 25596 8910 25648 8916
rect 26148 8968 26200 8974
rect 26148 8910 26200 8916
rect 26252 8906 26280 9846
rect 26436 9674 26464 9998
rect 26528 9926 26556 10610
rect 26516 9920 26568 9926
rect 26516 9862 26568 9868
rect 26344 9646 26464 9674
rect 26528 9674 26556 9862
rect 26528 9646 26648 9674
rect 25780 8900 25832 8906
rect 25780 8842 25832 8848
rect 25872 8900 25924 8906
rect 25872 8842 25924 8848
rect 26240 8900 26292 8906
rect 26240 8842 26292 8848
rect 25792 8566 25820 8842
rect 25780 8560 25832 8566
rect 25780 8502 25832 8508
rect 25504 8492 25556 8498
rect 25504 8434 25556 8440
rect 25228 8356 25280 8362
rect 25228 8298 25280 8304
rect 25240 8090 25268 8298
rect 25884 8276 25912 8842
rect 26240 8628 26292 8634
rect 26240 8570 26292 8576
rect 26146 8528 26202 8537
rect 26146 8463 26148 8472
rect 26200 8463 26202 8472
rect 26148 8434 26200 8440
rect 26252 8430 26280 8570
rect 26344 8566 26372 9646
rect 26620 9382 26648 9646
rect 26884 9512 26936 9518
rect 26884 9454 26936 9460
rect 26608 9376 26660 9382
rect 26608 9318 26660 9324
rect 26424 8900 26476 8906
rect 26424 8842 26476 8848
rect 26332 8560 26384 8566
rect 26332 8502 26384 8508
rect 26240 8424 26292 8430
rect 26240 8366 26292 8372
rect 25884 8248 26188 8276
rect 25740 8188 26048 8197
rect 25740 8186 25746 8188
rect 25802 8186 25826 8188
rect 25882 8186 25906 8188
rect 25962 8186 25986 8188
rect 26042 8186 26048 8188
rect 25802 8134 25804 8186
rect 25984 8134 25986 8186
rect 25740 8132 25746 8134
rect 25802 8132 25826 8134
rect 25882 8132 25906 8134
rect 25962 8132 25986 8134
rect 26042 8132 26048 8134
rect 25740 8123 26048 8132
rect 26160 8090 26188 8248
rect 25228 8084 25280 8090
rect 25228 8026 25280 8032
rect 26148 8084 26200 8090
rect 26148 8026 26200 8032
rect 26160 7954 26188 8026
rect 26148 7948 26200 7954
rect 26148 7890 26200 7896
rect 26252 7818 26280 8366
rect 25872 7812 25924 7818
rect 25872 7754 25924 7760
rect 26240 7812 26292 7818
rect 26240 7754 26292 7760
rect 25596 7744 25648 7750
rect 25596 7686 25648 7692
rect 25608 7546 25636 7686
rect 25884 7546 25912 7754
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25872 7540 25924 7546
rect 25872 7482 25924 7488
rect 26252 7410 26280 7754
rect 26436 7750 26464 8842
rect 26620 8498 26648 9318
rect 26896 9178 26924 9454
rect 26884 9172 26936 9178
rect 26884 9114 26936 9120
rect 27080 8906 27108 11086
rect 27068 8900 27120 8906
rect 27068 8842 27120 8848
rect 26608 8492 26660 8498
rect 26608 8434 26660 8440
rect 26608 8356 26660 8362
rect 26608 8298 26660 8304
rect 26620 7886 26648 8298
rect 26608 7880 26660 7886
rect 26608 7822 26660 7828
rect 26424 7744 26476 7750
rect 26424 7686 26476 7692
rect 26516 7472 26568 7478
rect 26516 7414 26568 7420
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 26240 7404 26292 7410
rect 26240 7346 26292 7352
rect 25740 7100 26048 7109
rect 25740 7098 25746 7100
rect 25802 7098 25826 7100
rect 25882 7098 25906 7100
rect 25962 7098 25986 7100
rect 26042 7098 26048 7100
rect 25802 7046 25804 7098
rect 25984 7046 25986 7098
rect 25740 7044 25746 7046
rect 25802 7044 25826 7046
rect 25882 7044 25906 7046
rect 25962 7044 25986 7046
rect 26042 7044 26048 7046
rect 25740 7035 26048 7044
rect 24768 6792 24820 6798
rect 24768 6734 24820 6740
rect 26528 6662 26556 7414
rect 26620 7410 26648 7822
rect 27080 7478 27108 8842
rect 27068 7472 27120 7478
rect 27068 7414 27120 7420
rect 26608 7404 26660 7410
rect 26608 7346 26660 7352
rect 26516 6656 26568 6662
rect 26516 6598 26568 6604
rect 25740 6012 26048 6021
rect 25740 6010 25746 6012
rect 25802 6010 25826 6012
rect 25882 6010 25906 6012
rect 25962 6010 25986 6012
rect 26042 6010 26048 6012
rect 25802 5958 25804 6010
rect 25984 5958 25986 6010
rect 25740 5956 25746 5958
rect 25802 5956 25826 5958
rect 25882 5956 25906 5958
rect 25962 5956 25986 5958
rect 26042 5956 26048 5958
rect 25740 5947 26048 5956
rect 25740 4924 26048 4933
rect 25740 4922 25746 4924
rect 25802 4922 25826 4924
rect 25882 4922 25906 4924
rect 25962 4922 25986 4924
rect 26042 4922 26048 4924
rect 25802 4870 25804 4922
rect 25984 4870 25986 4922
rect 25740 4868 25746 4870
rect 25802 4868 25826 4870
rect 25882 4868 25906 4870
rect 25962 4868 25986 4870
rect 26042 4868 26048 4870
rect 25740 4859 26048 4868
rect 24492 4140 24544 4146
rect 24492 4082 24544 4088
rect 24214 4040 24270 4049
rect 22100 4004 22152 4010
rect 24214 3975 24270 3984
rect 22100 3946 22152 3952
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20180 3602 20208 3878
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 22112 2446 22140 3946
rect 24400 3936 24452 3942
rect 24400 3878 24452 3884
rect 24952 3936 25004 3942
rect 24952 3878 25004 3884
rect 24412 3738 24440 3878
rect 24964 3738 24992 3878
rect 25740 3836 26048 3845
rect 25740 3834 25746 3836
rect 25802 3834 25826 3836
rect 25882 3834 25906 3836
rect 25962 3834 25986 3836
rect 26042 3834 26048 3836
rect 25802 3782 25804 3834
rect 25984 3782 25986 3834
rect 25740 3780 25746 3782
rect 25802 3780 25826 3782
rect 25882 3780 25906 3782
rect 25962 3780 25986 3782
rect 26042 3780 26048 3782
rect 25740 3771 26048 3780
rect 24400 3732 24452 3738
rect 24400 3674 24452 3680
rect 24952 3732 25004 3738
rect 24952 3674 25004 3680
rect 25228 3392 25280 3398
rect 25228 3334 25280 3340
rect 22198 3292 22506 3301
rect 22198 3290 22204 3292
rect 22260 3290 22284 3292
rect 22340 3290 22364 3292
rect 22420 3290 22444 3292
rect 22500 3290 22506 3292
rect 22260 3238 22262 3290
rect 22442 3238 22444 3290
rect 22198 3236 22204 3238
rect 22260 3236 22284 3238
rect 22340 3236 22364 3238
rect 22420 3236 22444 3238
rect 22500 3236 22506 3238
rect 22198 3227 22506 3236
rect 25240 2446 25268 3334
rect 27172 2774 27200 14878
rect 27712 14884 27764 14890
rect 27712 14826 27764 14832
rect 28184 14550 28212 14962
rect 28172 14544 28224 14550
rect 28172 14486 28224 14492
rect 28080 14340 28132 14346
rect 28080 14282 28132 14288
rect 28092 13870 28120 14282
rect 28080 13864 28132 13870
rect 28080 13806 28132 13812
rect 28172 9580 28224 9586
rect 28172 9522 28224 9528
rect 28080 9512 28132 9518
rect 28080 9454 28132 9460
rect 27896 9444 27948 9450
rect 27896 9386 27948 9392
rect 27252 9036 27304 9042
rect 27252 8978 27304 8984
rect 27264 8498 27292 8978
rect 27908 8974 27936 9386
rect 27896 8968 27948 8974
rect 27896 8910 27948 8916
rect 27804 8900 27856 8906
rect 27804 8842 27856 8848
rect 27816 8537 27844 8842
rect 28092 8566 28120 9454
rect 28184 8634 28212 9522
rect 28172 8628 28224 8634
rect 28172 8570 28224 8576
rect 28080 8560 28132 8566
rect 27802 8528 27858 8537
rect 27252 8492 27304 8498
rect 28080 8502 28132 8508
rect 27802 8463 27858 8472
rect 27252 8434 27304 8440
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27344 8288 27396 8294
rect 27344 8230 27396 8236
rect 27356 8090 27384 8230
rect 27344 8084 27396 8090
rect 27344 8026 27396 8032
rect 27356 7410 27384 8026
rect 27540 7954 27568 8366
rect 27528 7948 27580 7954
rect 27528 7890 27580 7896
rect 27540 7546 27568 7890
rect 27528 7540 27580 7546
rect 27528 7482 27580 7488
rect 27816 7410 27844 8463
rect 28092 8090 28120 8502
rect 28080 8084 28132 8090
rect 28080 8026 28132 8032
rect 27344 7404 27396 7410
rect 27344 7346 27396 7352
rect 27804 7404 27856 7410
rect 27804 7346 27856 7352
rect 28276 5370 28304 26930
rect 29000 26784 29052 26790
rect 29000 26726 29052 26732
rect 29012 26625 29040 26726
rect 28998 26616 29054 26625
rect 28998 26551 29054 26560
rect 29281 26140 29589 26149
rect 29281 26138 29287 26140
rect 29343 26138 29367 26140
rect 29423 26138 29447 26140
rect 29503 26138 29527 26140
rect 29583 26138 29589 26140
rect 29343 26086 29345 26138
rect 29525 26086 29527 26138
rect 29281 26084 29287 26086
rect 29343 26084 29367 26086
rect 29423 26084 29447 26086
rect 29503 26084 29527 26086
rect 29583 26084 29589 26086
rect 29281 26075 29589 26084
rect 29281 25052 29589 25061
rect 29281 25050 29287 25052
rect 29343 25050 29367 25052
rect 29423 25050 29447 25052
rect 29503 25050 29527 25052
rect 29583 25050 29589 25052
rect 29343 24998 29345 25050
rect 29525 24998 29527 25050
rect 29281 24996 29287 24998
rect 29343 24996 29367 24998
rect 29423 24996 29447 24998
rect 29503 24996 29527 24998
rect 29583 24996 29589 24998
rect 29281 24987 29589 24996
rect 29281 23964 29589 23973
rect 29281 23962 29287 23964
rect 29343 23962 29367 23964
rect 29423 23962 29447 23964
rect 29503 23962 29527 23964
rect 29583 23962 29589 23964
rect 29343 23910 29345 23962
rect 29525 23910 29527 23962
rect 29281 23908 29287 23910
rect 29343 23908 29367 23910
rect 29423 23908 29447 23910
rect 29503 23908 29527 23910
rect 29583 23908 29589 23910
rect 29281 23899 29589 23908
rect 29281 22876 29589 22885
rect 29281 22874 29287 22876
rect 29343 22874 29367 22876
rect 29423 22874 29447 22876
rect 29503 22874 29527 22876
rect 29583 22874 29589 22876
rect 29343 22822 29345 22874
rect 29525 22822 29527 22874
rect 29281 22820 29287 22822
rect 29343 22820 29367 22822
rect 29423 22820 29447 22822
rect 29503 22820 29527 22822
rect 29583 22820 29589 22822
rect 29281 22811 29589 22820
rect 28816 22636 28868 22642
rect 28816 22578 28868 22584
rect 28828 22030 28856 22578
rect 28998 22536 29054 22545
rect 28998 22471 29000 22480
rect 29052 22471 29054 22480
rect 29000 22442 29052 22448
rect 28816 22024 28868 22030
rect 28816 21966 28868 21972
rect 29281 21788 29589 21797
rect 29281 21786 29287 21788
rect 29343 21786 29367 21788
rect 29423 21786 29447 21788
rect 29503 21786 29527 21788
rect 29583 21786 29589 21788
rect 29343 21734 29345 21786
rect 29525 21734 29527 21786
rect 29281 21732 29287 21734
rect 29343 21732 29367 21734
rect 29423 21732 29447 21734
rect 29503 21732 29527 21734
rect 29583 21732 29589 21734
rect 29281 21723 29589 21732
rect 28908 21004 28960 21010
rect 28908 20946 28960 20952
rect 28540 20800 28592 20806
rect 28540 20742 28592 20748
rect 28552 20534 28580 20742
rect 28540 20528 28592 20534
rect 28540 20470 28592 20476
rect 28920 20466 28948 20946
rect 29281 20700 29589 20709
rect 29281 20698 29287 20700
rect 29343 20698 29367 20700
rect 29423 20698 29447 20700
rect 29503 20698 29527 20700
rect 29583 20698 29589 20700
rect 29343 20646 29345 20698
rect 29525 20646 29527 20698
rect 29281 20644 29287 20646
rect 29343 20644 29367 20646
rect 29423 20644 29447 20646
rect 29503 20644 29527 20646
rect 29583 20644 29589 20646
rect 29281 20635 29589 20644
rect 28908 20460 28960 20466
rect 28908 20402 28960 20408
rect 28356 20256 28408 20262
rect 28356 20198 28408 20204
rect 28368 19334 28396 20198
rect 28724 19712 28776 19718
rect 28724 19654 28776 19660
rect 28368 19306 28580 19334
rect 28448 17740 28500 17746
rect 28448 17682 28500 17688
rect 28356 17536 28408 17542
rect 28356 17478 28408 17484
rect 28368 17202 28396 17478
rect 28460 17270 28488 17682
rect 28448 17264 28500 17270
rect 28448 17206 28500 17212
rect 28356 17196 28408 17202
rect 28356 17138 28408 17144
rect 28448 17128 28500 17134
rect 28448 17070 28500 17076
rect 28356 16992 28408 16998
rect 28356 16934 28408 16940
rect 28368 16590 28396 16934
rect 28356 16584 28408 16590
rect 28356 16526 28408 16532
rect 28368 15638 28396 16526
rect 28356 15632 28408 15638
rect 28356 15574 28408 15580
rect 28460 13938 28488 17070
rect 28448 13932 28500 13938
rect 28448 13874 28500 13880
rect 28264 5364 28316 5370
rect 28264 5306 28316 5312
rect 28080 5228 28132 5234
rect 28080 5170 28132 5176
rect 28092 4826 28120 5170
rect 28080 4820 28132 4826
rect 28080 4762 28132 4768
rect 25740 2748 26048 2757
rect 25740 2746 25746 2748
rect 25802 2746 25826 2748
rect 25882 2746 25906 2748
rect 25962 2746 25986 2748
rect 26042 2746 26048 2748
rect 25802 2694 25804 2746
rect 25984 2694 25986 2746
rect 25740 2692 25746 2694
rect 25802 2692 25826 2694
rect 25882 2692 25906 2694
rect 25962 2692 25986 2694
rect 26042 2692 26048 2694
rect 25740 2683 26048 2692
rect 27080 2746 27200 2774
rect 27080 2582 27108 2746
rect 27068 2576 27120 2582
rect 27068 2518 27120 2524
rect 28552 2446 28580 19306
rect 28632 18284 28684 18290
rect 28632 18226 28684 18232
rect 28644 17134 28672 18226
rect 28632 17128 28684 17134
rect 28632 17070 28684 17076
rect 28632 16992 28684 16998
rect 28632 16934 28684 16940
rect 28644 16590 28672 16934
rect 28632 16584 28684 16590
rect 28632 16526 28684 16532
rect 28736 11150 28764 19654
rect 29281 19612 29589 19621
rect 29281 19610 29287 19612
rect 29343 19610 29367 19612
rect 29423 19610 29447 19612
rect 29503 19610 29527 19612
rect 29583 19610 29589 19612
rect 29343 19558 29345 19610
rect 29525 19558 29527 19610
rect 29281 19556 29287 19558
rect 29343 19556 29367 19558
rect 29423 19556 29447 19558
rect 29503 19556 29527 19558
rect 29583 19556 29589 19558
rect 29281 19547 29589 19556
rect 29460 18896 29512 18902
rect 29460 18838 29512 18844
rect 29472 18737 29500 18838
rect 29458 18728 29514 18737
rect 29458 18663 29514 18672
rect 29281 18524 29589 18533
rect 29281 18522 29287 18524
rect 29343 18522 29367 18524
rect 29423 18522 29447 18524
rect 29503 18522 29527 18524
rect 29583 18522 29589 18524
rect 29343 18470 29345 18522
rect 29525 18470 29527 18522
rect 29281 18468 29287 18470
rect 29343 18468 29367 18470
rect 29423 18468 29447 18470
rect 29503 18468 29527 18470
rect 29583 18468 29589 18470
rect 29281 18459 29589 18468
rect 29000 18216 29052 18222
rect 29000 18158 29052 18164
rect 29012 17746 29040 18158
rect 29000 17740 29052 17746
rect 29000 17682 29052 17688
rect 29281 17436 29589 17445
rect 29281 17434 29287 17436
rect 29343 17434 29367 17436
rect 29423 17434 29447 17436
rect 29503 17434 29527 17436
rect 29583 17434 29589 17436
rect 29343 17382 29345 17434
rect 29525 17382 29527 17434
rect 29281 17380 29287 17382
rect 29343 17380 29367 17382
rect 29423 17380 29447 17382
rect 29503 17380 29527 17382
rect 29583 17380 29589 17382
rect 29281 17371 29589 17380
rect 29281 16348 29589 16357
rect 29281 16346 29287 16348
rect 29343 16346 29367 16348
rect 29423 16346 29447 16348
rect 29503 16346 29527 16348
rect 29583 16346 29589 16348
rect 29343 16294 29345 16346
rect 29525 16294 29527 16346
rect 29281 16292 29287 16294
rect 29343 16292 29367 16294
rect 29423 16292 29447 16294
rect 29503 16292 29527 16294
rect 29583 16292 29589 16294
rect 29281 16283 29589 16292
rect 29281 15260 29589 15269
rect 29281 15258 29287 15260
rect 29343 15258 29367 15260
rect 29423 15258 29447 15260
rect 29503 15258 29527 15260
rect 29583 15258 29589 15260
rect 29343 15206 29345 15258
rect 29525 15206 29527 15258
rect 29281 15204 29287 15206
rect 29343 15204 29367 15206
rect 29423 15204 29447 15206
rect 29503 15204 29527 15206
rect 29583 15204 29589 15206
rect 29281 15195 29589 15204
rect 28998 14376 29054 14385
rect 28998 14311 29054 14320
rect 29012 13530 29040 14311
rect 29281 14172 29589 14181
rect 29281 14170 29287 14172
rect 29343 14170 29367 14172
rect 29423 14170 29447 14172
rect 29503 14170 29527 14172
rect 29583 14170 29589 14172
rect 29343 14118 29345 14170
rect 29525 14118 29527 14170
rect 29281 14116 29287 14118
rect 29343 14116 29367 14118
rect 29423 14116 29447 14118
rect 29503 14116 29527 14118
rect 29583 14116 29589 14118
rect 29281 14107 29589 14116
rect 29000 13524 29052 13530
rect 29000 13466 29052 13472
rect 29281 13084 29589 13093
rect 29281 13082 29287 13084
rect 29343 13082 29367 13084
rect 29423 13082 29447 13084
rect 29503 13082 29527 13084
rect 29583 13082 29589 13084
rect 29343 13030 29345 13082
rect 29525 13030 29527 13082
rect 29281 13028 29287 13030
rect 29343 13028 29367 13030
rect 29423 13028 29447 13030
rect 29503 13028 29527 13030
rect 29583 13028 29589 13030
rect 29281 13019 29589 13028
rect 29281 11996 29589 12005
rect 29281 11994 29287 11996
rect 29343 11994 29367 11996
rect 29423 11994 29447 11996
rect 29503 11994 29527 11996
rect 29583 11994 29589 11996
rect 29343 11942 29345 11994
rect 29525 11942 29527 11994
rect 29281 11940 29287 11942
rect 29343 11940 29367 11942
rect 29423 11940 29447 11942
rect 29503 11940 29527 11942
rect 29583 11940 29589 11942
rect 29281 11931 29589 11940
rect 28724 11144 28776 11150
rect 28724 11086 28776 11092
rect 29090 11112 29146 11121
rect 29090 11047 29092 11056
rect 29144 11047 29146 11056
rect 29092 11018 29144 11024
rect 29281 10908 29589 10917
rect 29281 10906 29287 10908
rect 29343 10906 29367 10908
rect 29423 10906 29447 10908
rect 29503 10906 29527 10908
rect 29583 10906 29589 10908
rect 29343 10854 29345 10906
rect 29525 10854 29527 10906
rect 29281 10852 29287 10854
rect 29343 10852 29367 10854
rect 29423 10852 29447 10854
rect 29503 10852 29527 10854
rect 29583 10852 29589 10854
rect 29281 10843 29589 10852
rect 29281 9820 29589 9829
rect 29281 9818 29287 9820
rect 29343 9818 29367 9820
rect 29423 9818 29447 9820
rect 29503 9818 29527 9820
rect 29583 9818 29589 9820
rect 29343 9766 29345 9818
rect 29525 9766 29527 9818
rect 29281 9764 29287 9766
rect 29343 9764 29367 9766
rect 29423 9764 29447 9766
rect 29503 9764 29527 9766
rect 29583 9764 29589 9766
rect 29281 9755 29589 9764
rect 29281 8732 29589 8741
rect 29281 8730 29287 8732
rect 29343 8730 29367 8732
rect 29423 8730 29447 8732
rect 29503 8730 29527 8732
rect 29583 8730 29589 8732
rect 29343 8678 29345 8730
rect 29525 8678 29527 8730
rect 29281 8676 29287 8678
rect 29343 8676 29367 8678
rect 29423 8676 29447 8678
rect 29503 8676 29527 8678
rect 29583 8676 29589 8678
rect 29281 8667 29589 8676
rect 29281 7644 29589 7653
rect 29281 7642 29287 7644
rect 29343 7642 29367 7644
rect 29423 7642 29447 7644
rect 29503 7642 29527 7644
rect 29583 7642 29589 7644
rect 29343 7590 29345 7642
rect 29525 7590 29527 7642
rect 29281 7588 29287 7590
rect 29343 7588 29367 7590
rect 29423 7588 29447 7590
rect 29503 7588 29527 7590
rect 29583 7588 29589 7590
rect 29281 7579 29589 7588
rect 28724 7404 28776 7410
rect 28724 7346 28776 7352
rect 28736 6458 28764 7346
rect 29000 7200 29052 7206
rect 29000 7142 29052 7148
rect 29012 6914 29040 7142
rect 29012 6905 29132 6914
rect 29012 6896 29146 6905
rect 29012 6886 29090 6896
rect 29090 6831 29146 6840
rect 29281 6556 29589 6565
rect 29281 6554 29287 6556
rect 29343 6554 29367 6556
rect 29423 6554 29447 6556
rect 29503 6554 29527 6556
rect 29583 6554 29589 6556
rect 29343 6502 29345 6554
rect 29525 6502 29527 6554
rect 29281 6500 29287 6502
rect 29343 6500 29367 6502
rect 29423 6500 29447 6502
rect 29503 6500 29527 6502
rect 29583 6500 29589 6502
rect 29281 6491 29589 6500
rect 28724 6452 28776 6458
rect 28724 6394 28776 6400
rect 29281 5468 29589 5477
rect 29281 5466 29287 5468
rect 29343 5466 29367 5468
rect 29423 5466 29447 5468
rect 29503 5466 29527 5468
rect 29583 5466 29589 5468
rect 29343 5414 29345 5466
rect 29525 5414 29527 5466
rect 29281 5412 29287 5414
rect 29343 5412 29367 5414
rect 29423 5412 29447 5414
rect 29503 5412 29527 5414
rect 29583 5412 29589 5414
rect 29281 5403 29589 5412
rect 29281 4380 29589 4389
rect 29281 4378 29287 4380
rect 29343 4378 29367 4380
rect 29423 4378 29447 4380
rect 29503 4378 29527 4380
rect 29583 4378 29589 4380
rect 29343 4326 29345 4378
rect 29525 4326 29527 4378
rect 29281 4324 29287 4326
rect 29343 4324 29367 4326
rect 29423 4324 29447 4326
rect 29503 4324 29527 4326
rect 29583 4324 29589 4326
rect 29281 4315 29589 4324
rect 29281 3292 29589 3301
rect 29281 3290 29287 3292
rect 29343 3290 29367 3292
rect 29423 3290 29447 3292
rect 29503 3290 29527 3292
rect 29583 3290 29589 3292
rect 29343 3238 29345 3290
rect 29525 3238 29527 3290
rect 29281 3236 29287 3238
rect 29343 3236 29367 3238
rect 29423 3236 29447 3238
rect 29503 3236 29527 3238
rect 29583 3236 29589 3238
rect 29281 3227 29589 3236
rect 29000 2848 29052 2854
rect 28998 2816 29000 2825
rect 29052 2816 29054 2825
rect 28998 2751 29054 2760
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 28540 2440 28592 2446
rect 28540 2382 28592 2388
rect 17500 2372 17552 2378
rect 17500 2314 17552 2320
rect 29644 2372 29696 2378
rect 29644 2314 29696 2320
rect 20 2304 72 2310
rect 3424 2304 3476 2310
rect 20 2246 72 2252
rect 3252 2264 3424 2292
rect 32 800 60 2246
rect 3252 800 3280 2264
rect 3424 2246 3476 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 22008 2304 22060 2310
rect 22008 2246 22060 2252
rect 26148 2304 26200 2310
rect 26148 2246 26200 2252
rect 7116 800 7144 2246
rect 8032 2204 8340 2213
rect 8032 2202 8038 2204
rect 8094 2202 8118 2204
rect 8174 2202 8198 2204
rect 8254 2202 8278 2204
rect 8334 2202 8340 2204
rect 8094 2150 8096 2202
rect 8276 2150 8278 2202
rect 8032 2148 8038 2150
rect 8094 2148 8118 2150
rect 8174 2148 8198 2150
rect 8254 2148 8278 2150
rect 8334 2148 8340 2150
rect 8032 2139 8340 2148
rect 11164 1442 11192 2246
rect 10980 1414 11192 1442
rect 10980 800 11008 1414
rect 14936 1170 14964 2246
rect 15115 2204 15423 2213
rect 15115 2202 15121 2204
rect 15177 2202 15201 2204
rect 15257 2202 15281 2204
rect 15337 2202 15361 2204
rect 15417 2202 15423 2204
rect 15177 2150 15179 2202
rect 15359 2150 15361 2202
rect 15115 2148 15121 2150
rect 15177 2148 15201 2150
rect 15257 2148 15281 2150
rect 15337 2148 15361 2150
rect 15417 2148 15423 2150
rect 15115 2139 15423 2148
rect 14844 1142 14964 1170
rect 14844 800 14872 1142
rect 18708 870 18828 898
rect 18708 800 18736 870
rect 18 0 74 800
rect 3238 0 3294 800
rect 7102 0 7158 800
rect 10966 0 11022 800
rect 14830 0 14886 800
rect 18694 0 18750 800
rect 18800 762 18828 870
rect 19076 762 19104 2246
rect 22020 1170 22048 2246
rect 22198 2204 22506 2213
rect 22198 2202 22204 2204
rect 22260 2202 22284 2204
rect 22340 2202 22364 2204
rect 22420 2202 22444 2204
rect 22500 2202 22506 2204
rect 22260 2150 22262 2202
rect 22442 2150 22444 2202
rect 22198 2148 22204 2150
rect 22260 2148 22284 2150
rect 22340 2148 22364 2150
rect 22420 2148 22444 2150
rect 22500 2148 22506 2150
rect 22198 2139 22506 2148
rect 21928 1142 22048 1170
rect 21928 800 21956 1142
rect 25792 870 25912 898
rect 25792 800 25820 870
rect 18800 734 19104 762
rect 21914 0 21970 800
rect 25778 0 25834 800
rect 25884 762 25912 870
rect 26160 762 26188 2246
rect 29281 2204 29589 2213
rect 29281 2202 29287 2204
rect 29343 2202 29367 2204
rect 29423 2202 29447 2204
rect 29503 2202 29527 2204
rect 29583 2202 29589 2204
rect 29343 2150 29345 2202
rect 29525 2150 29527 2202
rect 29281 2148 29287 2150
rect 29343 2148 29367 2150
rect 29423 2148 29447 2150
rect 29503 2148 29527 2150
rect 29583 2148 29589 2150
rect 29281 2139 29589 2148
rect 29656 800 29684 2314
rect 25884 734 26188 762
rect 29642 0 29698 800
<< via2 >>
rect 1582 30912 1638 30968
rect 8038 30490 8094 30492
rect 8118 30490 8174 30492
rect 8198 30490 8254 30492
rect 8278 30490 8334 30492
rect 8038 30438 8084 30490
rect 8084 30438 8094 30490
rect 8118 30438 8148 30490
rect 8148 30438 8160 30490
rect 8160 30438 8174 30490
rect 8198 30438 8212 30490
rect 8212 30438 8224 30490
rect 8224 30438 8254 30490
rect 8278 30438 8288 30490
rect 8288 30438 8334 30490
rect 8038 30436 8094 30438
rect 8118 30436 8174 30438
rect 8198 30436 8254 30438
rect 8278 30436 8334 30438
rect 15121 30490 15177 30492
rect 15201 30490 15257 30492
rect 15281 30490 15337 30492
rect 15361 30490 15417 30492
rect 15121 30438 15167 30490
rect 15167 30438 15177 30490
rect 15201 30438 15231 30490
rect 15231 30438 15243 30490
rect 15243 30438 15257 30490
rect 15281 30438 15295 30490
rect 15295 30438 15307 30490
rect 15307 30438 15337 30490
rect 15361 30438 15371 30490
rect 15371 30438 15417 30490
rect 15121 30436 15177 30438
rect 15201 30436 15257 30438
rect 15281 30436 15337 30438
rect 15361 30436 15417 30438
rect 938 27276 940 27296
rect 940 27276 992 27296
rect 992 27276 994 27296
rect 938 27240 994 27276
rect 1582 23468 1584 23488
rect 1584 23468 1636 23488
rect 1636 23468 1638 23488
rect 1582 23432 1638 23468
rect 1490 23024 1546 23080
rect 1582 19508 1638 19544
rect 1582 19488 1584 19508
rect 1584 19488 1636 19508
rect 1636 19488 1638 19508
rect 938 15680 994 15736
rect 938 11600 994 11656
rect 4497 29946 4553 29948
rect 4577 29946 4633 29948
rect 4657 29946 4713 29948
rect 4737 29946 4793 29948
rect 4497 29894 4543 29946
rect 4543 29894 4553 29946
rect 4577 29894 4607 29946
rect 4607 29894 4619 29946
rect 4619 29894 4633 29946
rect 4657 29894 4671 29946
rect 4671 29894 4683 29946
rect 4683 29894 4713 29946
rect 4737 29894 4747 29946
rect 4747 29894 4793 29946
rect 4497 29892 4553 29894
rect 4577 29892 4633 29894
rect 4657 29892 4713 29894
rect 4737 29892 4793 29894
rect 4497 28858 4553 28860
rect 4577 28858 4633 28860
rect 4657 28858 4713 28860
rect 4737 28858 4793 28860
rect 4497 28806 4543 28858
rect 4543 28806 4553 28858
rect 4577 28806 4607 28858
rect 4607 28806 4619 28858
rect 4619 28806 4633 28858
rect 4657 28806 4671 28858
rect 4671 28806 4683 28858
rect 4683 28806 4713 28858
rect 4737 28806 4747 28858
rect 4747 28806 4793 28858
rect 4497 28804 4553 28806
rect 4577 28804 4633 28806
rect 4657 28804 4713 28806
rect 4737 28804 4793 28806
rect 4497 27770 4553 27772
rect 4577 27770 4633 27772
rect 4657 27770 4713 27772
rect 4737 27770 4793 27772
rect 4497 27718 4543 27770
rect 4543 27718 4553 27770
rect 4577 27718 4607 27770
rect 4607 27718 4619 27770
rect 4619 27718 4633 27770
rect 4657 27718 4671 27770
rect 4671 27718 4683 27770
rect 4683 27718 4713 27770
rect 4737 27718 4747 27770
rect 4747 27718 4793 27770
rect 4497 27716 4553 27718
rect 4577 27716 4633 27718
rect 4657 27716 4713 27718
rect 4737 27716 4793 27718
rect 4497 26682 4553 26684
rect 4577 26682 4633 26684
rect 4657 26682 4713 26684
rect 4737 26682 4793 26684
rect 4497 26630 4543 26682
rect 4543 26630 4553 26682
rect 4577 26630 4607 26682
rect 4607 26630 4619 26682
rect 4619 26630 4633 26682
rect 4657 26630 4671 26682
rect 4671 26630 4683 26682
rect 4683 26630 4713 26682
rect 4737 26630 4747 26682
rect 4747 26630 4793 26682
rect 4497 26628 4553 26630
rect 4577 26628 4633 26630
rect 4657 26628 4713 26630
rect 4737 26628 4793 26630
rect 2226 11756 2282 11792
rect 2226 11736 2228 11756
rect 2228 11736 2280 11756
rect 2280 11736 2282 11756
rect 3054 12280 3110 12336
rect 1490 6296 1546 6352
rect 2410 3984 2466 4040
rect 4497 25594 4553 25596
rect 4577 25594 4633 25596
rect 4657 25594 4713 25596
rect 4737 25594 4793 25596
rect 4497 25542 4543 25594
rect 4543 25542 4553 25594
rect 4577 25542 4607 25594
rect 4607 25542 4619 25594
rect 4619 25542 4633 25594
rect 4657 25542 4671 25594
rect 4671 25542 4683 25594
rect 4683 25542 4713 25594
rect 4737 25542 4747 25594
rect 4747 25542 4793 25594
rect 4497 25540 4553 25542
rect 4577 25540 4633 25542
rect 4657 25540 4713 25542
rect 4737 25540 4793 25542
rect 4497 24506 4553 24508
rect 4577 24506 4633 24508
rect 4657 24506 4713 24508
rect 4737 24506 4793 24508
rect 4497 24454 4543 24506
rect 4543 24454 4553 24506
rect 4577 24454 4607 24506
rect 4607 24454 4619 24506
rect 4619 24454 4633 24506
rect 4657 24454 4671 24506
rect 4671 24454 4683 24506
rect 4683 24454 4713 24506
rect 4737 24454 4747 24506
rect 4747 24454 4793 24506
rect 4497 24452 4553 24454
rect 4577 24452 4633 24454
rect 4657 24452 4713 24454
rect 4737 24452 4793 24454
rect 4497 23418 4553 23420
rect 4577 23418 4633 23420
rect 4657 23418 4713 23420
rect 4737 23418 4793 23420
rect 4497 23366 4543 23418
rect 4543 23366 4553 23418
rect 4577 23366 4607 23418
rect 4607 23366 4619 23418
rect 4619 23366 4633 23418
rect 4657 23366 4671 23418
rect 4671 23366 4683 23418
rect 4683 23366 4713 23418
rect 4737 23366 4747 23418
rect 4747 23366 4793 23418
rect 4497 23364 4553 23366
rect 4577 23364 4633 23366
rect 4657 23364 4713 23366
rect 4737 23364 4793 23366
rect 4497 22330 4553 22332
rect 4577 22330 4633 22332
rect 4657 22330 4713 22332
rect 4737 22330 4793 22332
rect 4497 22278 4543 22330
rect 4543 22278 4553 22330
rect 4577 22278 4607 22330
rect 4607 22278 4619 22330
rect 4619 22278 4633 22330
rect 4657 22278 4671 22330
rect 4671 22278 4683 22330
rect 4683 22278 4713 22330
rect 4737 22278 4747 22330
rect 4747 22278 4793 22330
rect 4497 22276 4553 22278
rect 4577 22276 4633 22278
rect 4657 22276 4713 22278
rect 4737 22276 4793 22278
rect 4158 21528 4214 21584
rect 5446 21972 5448 21992
rect 5448 21972 5500 21992
rect 5500 21972 5502 21992
rect 5446 21936 5502 21972
rect 4497 21242 4553 21244
rect 4577 21242 4633 21244
rect 4657 21242 4713 21244
rect 4737 21242 4793 21244
rect 4497 21190 4543 21242
rect 4543 21190 4553 21242
rect 4577 21190 4607 21242
rect 4607 21190 4619 21242
rect 4619 21190 4633 21242
rect 4657 21190 4671 21242
rect 4671 21190 4683 21242
rect 4683 21190 4713 21242
rect 4737 21190 4747 21242
rect 4747 21190 4793 21242
rect 4497 21188 4553 21190
rect 4577 21188 4633 21190
rect 4657 21188 4713 21190
rect 4737 21188 4793 21190
rect 5814 21392 5870 21448
rect 5906 21256 5962 21312
rect 4894 20340 4896 20360
rect 4896 20340 4948 20360
rect 4948 20340 4950 20360
rect 4894 20304 4950 20340
rect 4497 20154 4553 20156
rect 4577 20154 4633 20156
rect 4657 20154 4713 20156
rect 4737 20154 4793 20156
rect 4497 20102 4543 20154
rect 4543 20102 4553 20154
rect 4577 20102 4607 20154
rect 4607 20102 4619 20154
rect 4619 20102 4633 20154
rect 4657 20102 4671 20154
rect 4671 20102 4683 20154
rect 4683 20102 4713 20154
rect 4737 20102 4747 20154
rect 4747 20102 4793 20154
rect 4497 20100 4553 20102
rect 4577 20100 4633 20102
rect 4657 20100 4713 20102
rect 4737 20100 4793 20102
rect 4497 19066 4553 19068
rect 4577 19066 4633 19068
rect 4657 19066 4713 19068
rect 4737 19066 4793 19068
rect 4497 19014 4543 19066
rect 4543 19014 4553 19066
rect 4577 19014 4607 19066
rect 4607 19014 4619 19066
rect 4619 19014 4633 19066
rect 4657 19014 4671 19066
rect 4671 19014 4683 19066
rect 4683 19014 4713 19066
rect 4737 19014 4747 19066
rect 4747 19014 4793 19066
rect 4497 19012 4553 19014
rect 4577 19012 4633 19014
rect 4657 19012 4713 19014
rect 4737 19012 4793 19014
rect 4497 17978 4553 17980
rect 4577 17978 4633 17980
rect 4657 17978 4713 17980
rect 4737 17978 4793 17980
rect 4497 17926 4543 17978
rect 4543 17926 4553 17978
rect 4577 17926 4607 17978
rect 4607 17926 4619 17978
rect 4619 17926 4633 17978
rect 4657 17926 4671 17978
rect 4671 17926 4683 17978
rect 4683 17926 4713 17978
rect 4737 17926 4747 17978
rect 4747 17926 4793 17978
rect 4497 17924 4553 17926
rect 4577 17924 4633 17926
rect 4657 17924 4713 17926
rect 4737 17924 4793 17926
rect 4618 17040 4674 17096
rect 4497 16890 4553 16892
rect 4577 16890 4633 16892
rect 4657 16890 4713 16892
rect 4737 16890 4793 16892
rect 4497 16838 4543 16890
rect 4543 16838 4553 16890
rect 4577 16838 4607 16890
rect 4607 16838 4619 16890
rect 4619 16838 4633 16890
rect 4657 16838 4671 16890
rect 4671 16838 4683 16890
rect 4683 16838 4713 16890
rect 4737 16838 4747 16890
rect 4747 16838 4793 16890
rect 4497 16836 4553 16838
rect 4577 16836 4633 16838
rect 4657 16836 4713 16838
rect 4737 16836 4793 16838
rect 5262 17060 5318 17096
rect 5262 17040 5264 17060
rect 5264 17040 5316 17060
rect 5316 17040 5318 17060
rect 4497 15802 4553 15804
rect 4577 15802 4633 15804
rect 4657 15802 4713 15804
rect 4737 15802 4793 15804
rect 4497 15750 4543 15802
rect 4543 15750 4553 15802
rect 4577 15750 4607 15802
rect 4607 15750 4619 15802
rect 4619 15750 4633 15802
rect 4657 15750 4671 15802
rect 4671 15750 4683 15802
rect 4683 15750 4713 15802
rect 4737 15750 4747 15802
rect 4747 15750 4793 15802
rect 4497 15748 4553 15750
rect 4577 15748 4633 15750
rect 4657 15748 4713 15750
rect 4737 15748 4793 15750
rect 4066 15444 4068 15464
rect 4068 15444 4120 15464
rect 4120 15444 4122 15464
rect 4066 15408 4122 15444
rect 4497 14714 4553 14716
rect 4577 14714 4633 14716
rect 4657 14714 4713 14716
rect 4737 14714 4793 14716
rect 4497 14662 4543 14714
rect 4543 14662 4553 14714
rect 4577 14662 4607 14714
rect 4607 14662 4619 14714
rect 4619 14662 4633 14714
rect 4657 14662 4671 14714
rect 4671 14662 4683 14714
rect 4683 14662 4713 14714
rect 4737 14662 4747 14714
rect 4747 14662 4793 14714
rect 4497 14660 4553 14662
rect 4577 14660 4633 14662
rect 4657 14660 4713 14662
rect 4737 14660 4793 14662
rect 3790 12144 3846 12200
rect 4497 13626 4553 13628
rect 4577 13626 4633 13628
rect 4657 13626 4713 13628
rect 4737 13626 4793 13628
rect 4497 13574 4543 13626
rect 4543 13574 4553 13626
rect 4577 13574 4607 13626
rect 4607 13574 4619 13626
rect 4619 13574 4633 13626
rect 4657 13574 4671 13626
rect 4671 13574 4683 13626
rect 4683 13574 4713 13626
rect 4737 13574 4747 13626
rect 4747 13574 4793 13626
rect 4497 13572 4553 13574
rect 4577 13572 4633 13574
rect 4657 13572 4713 13574
rect 4737 13572 4793 13574
rect 4497 12538 4553 12540
rect 4577 12538 4633 12540
rect 4657 12538 4713 12540
rect 4737 12538 4793 12540
rect 4497 12486 4543 12538
rect 4543 12486 4553 12538
rect 4577 12486 4607 12538
rect 4607 12486 4619 12538
rect 4619 12486 4633 12538
rect 4657 12486 4671 12538
rect 4671 12486 4683 12538
rect 4683 12486 4713 12538
rect 4737 12486 4747 12538
rect 4747 12486 4793 12538
rect 4497 12484 4553 12486
rect 4577 12484 4633 12486
rect 4657 12484 4713 12486
rect 4737 12484 4793 12486
rect 4497 11450 4553 11452
rect 4577 11450 4633 11452
rect 4657 11450 4713 11452
rect 4737 11450 4793 11452
rect 4497 11398 4543 11450
rect 4543 11398 4553 11450
rect 4577 11398 4607 11450
rect 4607 11398 4619 11450
rect 4619 11398 4633 11450
rect 4657 11398 4671 11450
rect 4671 11398 4683 11450
rect 4683 11398 4713 11450
rect 4737 11398 4747 11450
rect 4747 11398 4793 11450
rect 4497 11396 4553 11398
rect 4577 11396 4633 11398
rect 4657 11396 4713 11398
rect 4737 11396 4793 11398
rect 4066 9424 4122 9480
rect 4497 10362 4553 10364
rect 4577 10362 4633 10364
rect 4657 10362 4713 10364
rect 4737 10362 4793 10364
rect 4497 10310 4543 10362
rect 4543 10310 4553 10362
rect 4577 10310 4607 10362
rect 4607 10310 4619 10362
rect 4619 10310 4633 10362
rect 4657 10310 4671 10362
rect 4671 10310 4683 10362
rect 4683 10310 4713 10362
rect 4737 10310 4747 10362
rect 4747 10310 4793 10362
rect 4497 10308 4553 10310
rect 4577 10308 4633 10310
rect 4657 10308 4713 10310
rect 4737 10308 4793 10310
rect 4497 9274 4553 9276
rect 4577 9274 4633 9276
rect 4657 9274 4713 9276
rect 4737 9274 4793 9276
rect 4497 9222 4543 9274
rect 4543 9222 4553 9274
rect 4577 9222 4607 9274
rect 4607 9222 4619 9274
rect 4619 9222 4633 9274
rect 4657 9222 4671 9274
rect 4671 9222 4683 9274
rect 4683 9222 4713 9274
rect 4737 9222 4747 9274
rect 4747 9222 4793 9274
rect 4497 9220 4553 9222
rect 4577 9220 4633 9222
rect 4657 9220 4713 9222
rect 4737 9220 4793 9222
rect 5170 12144 5226 12200
rect 4497 8186 4553 8188
rect 4577 8186 4633 8188
rect 4657 8186 4713 8188
rect 4737 8186 4793 8188
rect 4497 8134 4543 8186
rect 4543 8134 4553 8186
rect 4577 8134 4607 8186
rect 4607 8134 4619 8186
rect 4619 8134 4633 8186
rect 4657 8134 4671 8186
rect 4671 8134 4683 8186
rect 4683 8134 4713 8186
rect 4737 8134 4747 8186
rect 4747 8134 4793 8186
rect 4497 8132 4553 8134
rect 4577 8132 4633 8134
rect 4657 8132 4713 8134
rect 4737 8132 4793 8134
rect 8038 29402 8094 29404
rect 8118 29402 8174 29404
rect 8198 29402 8254 29404
rect 8278 29402 8334 29404
rect 8038 29350 8084 29402
rect 8084 29350 8094 29402
rect 8118 29350 8148 29402
rect 8148 29350 8160 29402
rect 8160 29350 8174 29402
rect 8198 29350 8212 29402
rect 8212 29350 8224 29402
rect 8224 29350 8254 29402
rect 8278 29350 8288 29402
rect 8288 29350 8334 29402
rect 8038 29348 8094 29350
rect 8118 29348 8174 29350
rect 8198 29348 8254 29350
rect 8278 29348 8334 29350
rect 8038 28314 8094 28316
rect 8118 28314 8174 28316
rect 8198 28314 8254 28316
rect 8278 28314 8334 28316
rect 8038 28262 8084 28314
rect 8084 28262 8094 28314
rect 8118 28262 8148 28314
rect 8148 28262 8160 28314
rect 8160 28262 8174 28314
rect 8198 28262 8212 28314
rect 8212 28262 8224 28314
rect 8224 28262 8254 28314
rect 8278 28262 8288 28314
rect 8288 28262 8334 28314
rect 8038 28260 8094 28262
rect 8118 28260 8174 28262
rect 8198 28260 8254 28262
rect 8278 28260 8334 28262
rect 8038 27226 8094 27228
rect 8118 27226 8174 27228
rect 8198 27226 8254 27228
rect 8278 27226 8334 27228
rect 8038 27174 8084 27226
rect 8084 27174 8094 27226
rect 8118 27174 8148 27226
rect 8148 27174 8160 27226
rect 8160 27174 8174 27226
rect 8198 27174 8212 27226
rect 8212 27174 8224 27226
rect 8224 27174 8254 27226
rect 8278 27174 8288 27226
rect 8288 27174 8334 27226
rect 8038 27172 8094 27174
rect 8118 27172 8174 27174
rect 8198 27172 8254 27174
rect 8278 27172 8334 27174
rect 8038 26138 8094 26140
rect 8118 26138 8174 26140
rect 8198 26138 8254 26140
rect 8278 26138 8334 26140
rect 8038 26086 8084 26138
rect 8084 26086 8094 26138
rect 8118 26086 8148 26138
rect 8148 26086 8160 26138
rect 8160 26086 8174 26138
rect 8198 26086 8212 26138
rect 8212 26086 8224 26138
rect 8224 26086 8254 26138
rect 8278 26086 8288 26138
rect 8288 26086 8334 26138
rect 8038 26084 8094 26086
rect 8118 26084 8174 26086
rect 8198 26084 8254 26086
rect 8278 26084 8334 26086
rect 8038 25050 8094 25052
rect 8118 25050 8174 25052
rect 8198 25050 8254 25052
rect 8278 25050 8334 25052
rect 8038 24998 8084 25050
rect 8084 24998 8094 25050
rect 8118 24998 8148 25050
rect 8148 24998 8160 25050
rect 8160 24998 8174 25050
rect 8198 24998 8212 25050
rect 8212 24998 8224 25050
rect 8224 24998 8254 25050
rect 8278 24998 8288 25050
rect 8288 24998 8334 25050
rect 8038 24996 8094 24998
rect 8118 24996 8174 24998
rect 8198 24996 8254 24998
rect 8278 24996 8334 24998
rect 8038 23962 8094 23964
rect 8118 23962 8174 23964
rect 8198 23962 8254 23964
rect 8278 23962 8334 23964
rect 8038 23910 8084 23962
rect 8084 23910 8094 23962
rect 8118 23910 8148 23962
rect 8148 23910 8160 23962
rect 8160 23910 8174 23962
rect 8198 23910 8212 23962
rect 8212 23910 8224 23962
rect 8224 23910 8254 23962
rect 8278 23910 8288 23962
rect 8288 23910 8334 23962
rect 8038 23908 8094 23910
rect 8118 23908 8174 23910
rect 8198 23908 8254 23910
rect 8278 23908 8334 23910
rect 8038 22874 8094 22876
rect 8118 22874 8174 22876
rect 8198 22874 8254 22876
rect 8278 22874 8334 22876
rect 8038 22822 8084 22874
rect 8084 22822 8094 22874
rect 8118 22822 8148 22874
rect 8148 22822 8160 22874
rect 8160 22822 8174 22874
rect 8198 22822 8212 22874
rect 8212 22822 8224 22874
rect 8224 22822 8254 22874
rect 8278 22822 8288 22874
rect 8288 22822 8334 22874
rect 8038 22820 8094 22822
rect 8118 22820 8174 22822
rect 8198 22820 8254 22822
rect 8278 22820 8334 22822
rect 7286 21936 7342 21992
rect 6918 21528 6974 21584
rect 8114 22208 8170 22264
rect 6642 15444 6644 15464
rect 6644 15444 6696 15464
rect 6696 15444 6698 15464
rect 6642 15408 6698 15444
rect 8038 21786 8094 21788
rect 8118 21786 8174 21788
rect 8198 21786 8254 21788
rect 8278 21786 8334 21788
rect 8038 21734 8084 21786
rect 8084 21734 8094 21786
rect 8118 21734 8148 21786
rect 8148 21734 8160 21786
rect 8160 21734 8174 21786
rect 8198 21734 8212 21786
rect 8212 21734 8224 21786
rect 8224 21734 8254 21786
rect 8278 21734 8288 21786
rect 8288 21734 8334 21786
rect 8038 21732 8094 21734
rect 8118 21732 8174 21734
rect 8198 21732 8254 21734
rect 8278 21732 8334 21734
rect 7102 17604 7158 17640
rect 7102 17584 7104 17604
rect 7104 17584 7156 17604
rect 7156 17584 7158 17604
rect 8390 21392 8446 21448
rect 8574 21256 8630 21312
rect 8038 20698 8094 20700
rect 8118 20698 8174 20700
rect 8198 20698 8254 20700
rect 8278 20698 8334 20700
rect 8038 20646 8084 20698
rect 8084 20646 8094 20698
rect 8118 20646 8148 20698
rect 8148 20646 8160 20698
rect 8160 20646 8174 20698
rect 8198 20646 8212 20698
rect 8212 20646 8224 20698
rect 8224 20646 8254 20698
rect 8278 20646 8288 20698
rect 8288 20646 8334 20698
rect 8038 20644 8094 20646
rect 8118 20644 8174 20646
rect 8198 20644 8254 20646
rect 8278 20644 8334 20646
rect 8038 19610 8094 19612
rect 8118 19610 8174 19612
rect 8198 19610 8254 19612
rect 8278 19610 8334 19612
rect 8038 19558 8084 19610
rect 8084 19558 8094 19610
rect 8118 19558 8148 19610
rect 8148 19558 8160 19610
rect 8160 19558 8174 19610
rect 8198 19558 8212 19610
rect 8212 19558 8224 19610
rect 8224 19558 8254 19610
rect 8278 19558 8288 19610
rect 8288 19558 8334 19610
rect 8038 19556 8094 19558
rect 8118 19556 8174 19558
rect 8198 19556 8254 19558
rect 8278 19556 8334 19558
rect 8038 18522 8094 18524
rect 8118 18522 8174 18524
rect 8198 18522 8254 18524
rect 8278 18522 8334 18524
rect 8038 18470 8084 18522
rect 8084 18470 8094 18522
rect 8118 18470 8148 18522
rect 8148 18470 8160 18522
rect 8160 18470 8174 18522
rect 8198 18470 8212 18522
rect 8212 18470 8224 18522
rect 8224 18470 8254 18522
rect 8278 18470 8288 18522
rect 8288 18470 8334 18522
rect 8038 18468 8094 18470
rect 8118 18468 8174 18470
rect 8198 18468 8254 18470
rect 8278 18468 8334 18470
rect 5446 9560 5502 9616
rect 5446 8492 5502 8528
rect 5446 8472 5448 8492
rect 5448 8472 5500 8492
rect 5500 8472 5502 8492
rect 4066 7520 4122 7576
rect 4497 7098 4553 7100
rect 4577 7098 4633 7100
rect 4657 7098 4713 7100
rect 4737 7098 4793 7100
rect 4497 7046 4543 7098
rect 4543 7046 4553 7098
rect 4577 7046 4607 7098
rect 4607 7046 4619 7098
rect 4619 7046 4633 7098
rect 4657 7046 4671 7098
rect 4671 7046 4683 7098
rect 4683 7046 4713 7098
rect 4737 7046 4747 7098
rect 4747 7046 4793 7098
rect 4497 7044 4553 7046
rect 4577 7044 4633 7046
rect 4657 7044 4713 7046
rect 4737 7044 4793 7046
rect 6918 9424 6974 9480
rect 5998 6740 6000 6760
rect 6000 6740 6052 6760
rect 6052 6740 6054 6760
rect 5998 6704 6054 6740
rect 4497 6010 4553 6012
rect 4577 6010 4633 6012
rect 4657 6010 4713 6012
rect 4737 6010 4793 6012
rect 4497 5958 4543 6010
rect 4543 5958 4553 6010
rect 4577 5958 4607 6010
rect 4607 5958 4619 6010
rect 4619 5958 4633 6010
rect 4657 5958 4671 6010
rect 4671 5958 4683 6010
rect 4683 5958 4713 6010
rect 4737 5958 4747 6010
rect 4747 5958 4793 6010
rect 4497 5956 4553 5958
rect 4577 5956 4633 5958
rect 4657 5956 4713 5958
rect 4737 5956 4793 5958
rect 4497 4922 4553 4924
rect 4577 4922 4633 4924
rect 4657 4922 4713 4924
rect 4737 4922 4793 4924
rect 4497 4870 4543 4922
rect 4543 4870 4553 4922
rect 4577 4870 4607 4922
rect 4607 4870 4619 4922
rect 4619 4870 4633 4922
rect 4657 4870 4671 4922
rect 4671 4870 4683 4922
rect 4683 4870 4713 4922
rect 4737 4870 4747 4922
rect 4747 4870 4793 4922
rect 4497 4868 4553 4870
rect 4577 4868 4633 4870
rect 4657 4868 4713 4870
rect 4737 4868 4793 4870
rect 8038 17434 8094 17436
rect 8118 17434 8174 17436
rect 8198 17434 8254 17436
rect 8278 17434 8334 17436
rect 8038 17382 8084 17434
rect 8084 17382 8094 17434
rect 8118 17382 8148 17434
rect 8148 17382 8160 17434
rect 8160 17382 8174 17434
rect 8198 17382 8212 17434
rect 8212 17382 8224 17434
rect 8224 17382 8254 17434
rect 8278 17382 8288 17434
rect 8288 17382 8334 17434
rect 8038 17380 8094 17382
rect 8118 17380 8174 17382
rect 8198 17380 8254 17382
rect 8278 17380 8334 17382
rect 8038 16346 8094 16348
rect 8118 16346 8174 16348
rect 8198 16346 8254 16348
rect 8278 16346 8334 16348
rect 8038 16294 8084 16346
rect 8084 16294 8094 16346
rect 8118 16294 8148 16346
rect 8148 16294 8160 16346
rect 8160 16294 8174 16346
rect 8198 16294 8212 16346
rect 8212 16294 8224 16346
rect 8224 16294 8254 16346
rect 8278 16294 8288 16346
rect 8288 16294 8334 16346
rect 8038 16292 8094 16294
rect 8118 16292 8174 16294
rect 8198 16292 8254 16294
rect 8278 16292 8334 16294
rect 8038 15258 8094 15260
rect 8118 15258 8174 15260
rect 8198 15258 8254 15260
rect 8278 15258 8334 15260
rect 8038 15206 8084 15258
rect 8084 15206 8094 15258
rect 8118 15206 8148 15258
rect 8148 15206 8160 15258
rect 8160 15206 8174 15258
rect 8198 15206 8212 15258
rect 8212 15206 8224 15258
rect 8224 15206 8254 15258
rect 8278 15206 8288 15258
rect 8288 15206 8334 15258
rect 8038 15204 8094 15206
rect 8118 15204 8174 15206
rect 8198 15204 8254 15206
rect 8278 15204 8334 15206
rect 8038 14170 8094 14172
rect 8118 14170 8174 14172
rect 8198 14170 8254 14172
rect 8278 14170 8334 14172
rect 8038 14118 8084 14170
rect 8084 14118 8094 14170
rect 8118 14118 8148 14170
rect 8148 14118 8160 14170
rect 8160 14118 8174 14170
rect 8198 14118 8212 14170
rect 8212 14118 8224 14170
rect 8224 14118 8254 14170
rect 8278 14118 8288 14170
rect 8288 14118 8334 14170
rect 8038 14116 8094 14118
rect 8118 14116 8174 14118
rect 8198 14116 8254 14118
rect 8278 14116 8334 14118
rect 11580 29946 11636 29948
rect 11660 29946 11716 29948
rect 11740 29946 11796 29948
rect 11820 29946 11876 29948
rect 11580 29894 11626 29946
rect 11626 29894 11636 29946
rect 11660 29894 11690 29946
rect 11690 29894 11702 29946
rect 11702 29894 11716 29946
rect 11740 29894 11754 29946
rect 11754 29894 11766 29946
rect 11766 29894 11796 29946
rect 11820 29894 11830 29946
rect 11830 29894 11876 29946
rect 11580 29892 11636 29894
rect 11660 29892 11716 29894
rect 11740 29892 11796 29894
rect 11820 29892 11876 29894
rect 11058 28056 11114 28112
rect 11580 28858 11636 28860
rect 11660 28858 11716 28860
rect 11740 28858 11796 28860
rect 11820 28858 11876 28860
rect 11580 28806 11626 28858
rect 11626 28806 11636 28858
rect 11660 28806 11690 28858
rect 11690 28806 11702 28858
rect 11702 28806 11716 28858
rect 11740 28806 11754 28858
rect 11754 28806 11766 28858
rect 11766 28806 11796 28858
rect 11820 28806 11830 28858
rect 11830 28806 11876 28858
rect 11580 28804 11636 28806
rect 11660 28804 11716 28806
rect 11740 28804 11796 28806
rect 11820 28804 11876 28806
rect 12346 28056 12402 28112
rect 11580 27770 11636 27772
rect 11660 27770 11716 27772
rect 11740 27770 11796 27772
rect 11820 27770 11876 27772
rect 11580 27718 11626 27770
rect 11626 27718 11636 27770
rect 11660 27718 11690 27770
rect 11690 27718 11702 27770
rect 11702 27718 11716 27770
rect 11740 27718 11754 27770
rect 11754 27718 11766 27770
rect 11766 27718 11796 27770
rect 11820 27718 11830 27770
rect 11830 27718 11876 27770
rect 11580 27716 11636 27718
rect 11660 27716 11716 27718
rect 11740 27716 11796 27718
rect 11820 27716 11876 27718
rect 13634 28620 13690 28656
rect 13634 28600 13636 28620
rect 13636 28600 13688 28620
rect 13688 28600 13690 28620
rect 13634 28484 13690 28520
rect 13634 28464 13636 28484
rect 13636 28464 13688 28484
rect 13688 28464 13690 28484
rect 13358 27920 13414 27976
rect 11580 26682 11636 26684
rect 11660 26682 11716 26684
rect 11740 26682 11796 26684
rect 11820 26682 11876 26684
rect 11580 26630 11626 26682
rect 11626 26630 11636 26682
rect 11660 26630 11690 26682
rect 11690 26630 11702 26682
rect 11702 26630 11716 26682
rect 11740 26630 11754 26682
rect 11754 26630 11766 26682
rect 11766 26630 11796 26682
rect 11820 26630 11830 26682
rect 11830 26630 11876 26682
rect 11580 26628 11636 26630
rect 11660 26628 11716 26630
rect 11740 26628 11796 26630
rect 11820 26628 11876 26630
rect 11580 25594 11636 25596
rect 11660 25594 11716 25596
rect 11740 25594 11796 25596
rect 11820 25594 11876 25596
rect 11580 25542 11626 25594
rect 11626 25542 11636 25594
rect 11660 25542 11690 25594
rect 11690 25542 11702 25594
rect 11702 25542 11716 25594
rect 11740 25542 11754 25594
rect 11754 25542 11766 25594
rect 11766 25542 11796 25594
rect 11820 25542 11830 25594
rect 11830 25542 11876 25594
rect 11580 25540 11636 25542
rect 11660 25540 11716 25542
rect 11740 25540 11796 25542
rect 11820 25540 11876 25542
rect 9862 21392 9918 21448
rect 9862 20304 9918 20360
rect 10138 19352 10194 19408
rect 10598 22228 10654 22264
rect 10598 22208 10600 22228
rect 10600 22208 10652 22228
rect 10652 22208 10654 22228
rect 11580 24506 11636 24508
rect 11660 24506 11716 24508
rect 11740 24506 11796 24508
rect 11820 24506 11876 24508
rect 11580 24454 11626 24506
rect 11626 24454 11636 24506
rect 11660 24454 11690 24506
rect 11690 24454 11702 24506
rect 11702 24454 11716 24506
rect 11740 24454 11754 24506
rect 11754 24454 11766 24506
rect 11766 24454 11796 24506
rect 11820 24454 11830 24506
rect 11830 24454 11876 24506
rect 11580 24452 11636 24454
rect 11660 24452 11716 24454
rect 11740 24452 11796 24454
rect 11820 24452 11876 24454
rect 11580 23418 11636 23420
rect 11660 23418 11716 23420
rect 11740 23418 11796 23420
rect 11820 23418 11876 23420
rect 11580 23366 11626 23418
rect 11626 23366 11636 23418
rect 11660 23366 11690 23418
rect 11690 23366 11702 23418
rect 11702 23366 11716 23418
rect 11740 23366 11754 23418
rect 11754 23366 11766 23418
rect 11766 23366 11796 23418
rect 11820 23366 11830 23418
rect 11830 23366 11876 23418
rect 11580 23364 11636 23366
rect 11660 23364 11716 23366
rect 11740 23364 11796 23366
rect 11820 23364 11876 23366
rect 8038 13082 8094 13084
rect 8118 13082 8174 13084
rect 8198 13082 8254 13084
rect 8278 13082 8334 13084
rect 8038 13030 8084 13082
rect 8084 13030 8094 13082
rect 8118 13030 8148 13082
rect 8148 13030 8160 13082
rect 8160 13030 8174 13082
rect 8198 13030 8212 13082
rect 8212 13030 8224 13082
rect 8224 13030 8254 13082
rect 8278 13030 8288 13082
rect 8288 13030 8334 13082
rect 8038 13028 8094 13030
rect 8118 13028 8174 13030
rect 8198 13028 8254 13030
rect 8278 13028 8334 13030
rect 10414 19896 10470 19952
rect 10138 13912 10194 13968
rect 9678 13404 9680 13424
rect 9680 13404 9732 13424
rect 9732 13404 9734 13424
rect 9678 13368 9734 13404
rect 11580 22330 11636 22332
rect 11660 22330 11716 22332
rect 11740 22330 11796 22332
rect 11820 22330 11876 22332
rect 11580 22278 11626 22330
rect 11626 22278 11636 22330
rect 11660 22278 11690 22330
rect 11690 22278 11702 22330
rect 11702 22278 11716 22330
rect 11740 22278 11754 22330
rect 11754 22278 11766 22330
rect 11766 22278 11796 22330
rect 11820 22278 11830 22330
rect 11830 22278 11876 22330
rect 11580 22276 11636 22278
rect 11660 22276 11716 22278
rect 11740 22276 11796 22278
rect 11820 22276 11876 22278
rect 11580 21242 11636 21244
rect 11660 21242 11716 21244
rect 11740 21242 11796 21244
rect 11820 21242 11876 21244
rect 11580 21190 11626 21242
rect 11626 21190 11636 21242
rect 11660 21190 11690 21242
rect 11690 21190 11702 21242
rect 11702 21190 11716 21242
rect 11740 21190 11754 21242
rect 11754 21190 11766 21242
rect 11766 21190 11796 21242
rect 11820 21190 11830 21242
rect 11830 21190 11876 21242
rect 11580 21188 11636 21190
rect 11660 21188 11716 21190
rect 11740 21188 11796 21190
rect 11820 21188 11876 21190
rect 11242 20596 11298 20632
rect 11242 20576 11244 20596
rect 11244 20576 11296 20596
rect 11296 20576 11298 20596
rect 11580 20154 11636 20156
rect 11660 20154 11716 20156
rect 11740 20154 11796 20156
rect 11820 20154 11876 20156
rect 11580 20102 11626 20154
rect 11626 20102 11636 20154
rect 11660 20102 11690 20154
rect 11690 20102 11702 20154
rect 11702 20102 11716 20154
rect 11740 20102 11754 20154
rect 11754 20102 11766 20154
rect 11766 20102 11796 20154
rect 11820 20102 11830 20154
rect 11830 20102 11876 20154
rect 11580 20100 11636 20102
rect 11660 20100 11716 20102
rect 11740 20100 11796 20102
rect 11820 20100 11876 20102
rect 11580 19066 11636 19068
rect 11660 19066 11716 19068
rect 11740 19066 11796 19068
rect 11820 19066 11876 19068
rect 11580 19014 11626 19066
rect 11626 19014 11636 19066
rect 11660 19014 11690 19066
rect 11690 19014 11702 19066
rect 11702 19014 11716 19066
rect 11740 19014 11754 19066
rect 11754 19014 11766 19066
rect 11766 19014 11796 19066
rect 11820 19014 11830 19066
rect 11830 19014 11876 19066
rect 11580 19012 11636 19014
rect 11660 19012 11716 19014
rect 11740 19012 11796 19014
rect 11820 19012 11876 19014
rect 11580 17978 11636 17980
rect 11660 17978 11716 17980
rect 11740 17978 11796 17980
rect 11820 17978 11876 17980
rect 11580 17926 11626 17978
rect 11626 17926 11636 17978
rect 11660 17926 11690 17978
rect 11690 17926 11702 17978
rect 11702 17926 11716 17978
rect 11740 17926 11754 17978
rect 11754 17926 11766 17978
rect 11766 17926 11796 17978
rect 11820 17926 11830 17978
rect 11830 17926 11876 17978
rect 11580 17924 11636 17926
rect 11660 17924 11716 17926
rect 11740 17924 11796 17926
rect 11820 17924 11876 17926
rect 12070 19796 12072 19816
rect 12072 19796 12124 19816
rect 12124 19796 12126 19816
rect 12070 19760 12126 19796
rect 12622 20848 12678 20904
rect 10506 15544 10562 15600
rect 8038 11994 8094 11996
rect 8118 11994 8174 11996
rect 8198 11994 8254 11996
rect 8278 11994 8334 11996
rect 8038 11942 8084 11994
rect 8084 11942 8094 11994
rect 8118 11942 8148 11994
rect 8148 11942 8160 11994
rect 8160 11942 8174 11994
rect 8198 11942 8212 11994
rect 8212 11942 8224 11994
rect 8224 11942 8254 11994
rect 8278 11942 8288 11994
rect 8288 11942 8334 11994
rect 8038 11940 8094 11942
rect 8118 11940 8174 11942
rect 8198 11940 8254 11942
rect 8278 11940 8334 11942
rect 8038 10906 8094 10908
rect 8118 10906 8174 10908
rect 8198 10906 8254 10908
rect 8278 10906 8334 10908
rect 8038 10854 8084 10906
rect 8084 10854 8094 10906
rect 8118 10854 8148 10906
rect 8148 10854 8160 10906
rect 8160 10854 8174 10906
rect 8198 10854 8212 10906
rect 8212 10854 8224 10906
rect 8224 10854 8254 10906
rect 8278 10854 8288 10906
rect 8288 10854 8334 10906
rect 8038 10852 8094 10854
rect 8118 10852 8174 10854
rect 8198 10852 8254 10854
rect 8278 10852 8334 10854
rect 8038 9818 8094 9820
rect 8118 9818 8174 9820
rect 8198 9818 8254 9820
rect 8278 9818 8334 9820
rect 8038 9766 8084 9818
rect 8084 9766 8094 9818
rect 8118 9766 8148 9818
rect 8148 9766 8160 9818
rect 8160 9766 8174 9818
rect 8198 9766 8212 9818
rect 8212 9766 8224 9818
rect 8224 9766 8254 9818
rect 8278 9766 8288 9818
rect 8288 9766 8334 9818
rect 8038 9764 8094 9766
rect 8118 9764 8174 9766
rect 8198 9764 8254 9766
rect 8278 9764 8334 9766
rect 8850 9460 8852 9480
rect 8852 9460 8904 9480
rect 8904 9460 8906 9480
rect 8850 9424 8906 9460
rect 8038 8730 8094 8732
rect 8118 8730 8174 8732
rect 8198 8730 8254 8732
rect 8278 8730 8334 8732
rect 8038 8678 8084 8730
rect 8084 8678 8094 8730
rect 8118 8678 8148 8730
rect 8148 8678 8160 8730
rect 8160 8678 8174 8730
rect 8198 8678 8212 8730
rect 8212 8678 8224 8730
rect 8224 8678 8254 8730
rect 8278 8678 8288 8730
rect 8288 8678 8334 8730
rect 8038 8676 8094 8678
rect 8118 8676 8174 8678
rect 8198 8676 8254 8678
rect 8278 8676 8334 8678
rect 7746 6724 7802 6760
rect 7746 6704 7748 6724
rect 7748 6704 7800 6724
rect 7800 6704 7802 6724
rect 8038 7642 8094 7644
rect 8118 7642 8174 7644
rect 8198 7642 8254 7644
rect 8278 7642 8334 7644
rect 8038 7590 8084 7642
rect 8084 7590 8094 7642
rect 8118 7590 8148 7642
rect 8148 7590 8160 7642
rect 8160 7590 8174 7642
rect 8198 7590 8212 7642
rect 8212 7590 8224 7642
rect 8224 7590 8254 7642
rect 8278 7590 8288 7642
rect 8288 7590 8334 7642
rect 8038 7588 8094 7590
rect 8118 7588 8174 7590
rect 8198 7588 8254 7590
rect 8278 7588 8334 7590
rect 8038 6554 8094 6556
rect 8118 6554 8174 6556
rect 8198 6554 8254 6556
rect 8278 6554 8334 6556
rect 8038 6502 8084 6554
rect 8084 6502 8094 6554
rect 8118 6502 8148 6554
rect 8148 6502 8160 6554
rect 8160 6502 8174 6554
rect 8198 6502 8212 6554
rect 8212 6502 8224 6554
rect 8224 6502 8254 6554
rect 8278 6502 8288 6554
rect 8288 6502 8334 6554
rect 8038 6500 8094 6502
rect 8118 6500 8174 6502
rect 8198 6500 8254 6502
rect 8278 6500 8334 6502
rect 8038 5466 8094 5468
rect 8118 5466 8174 5468
rect 8198 5466 8254 5468
rect 8278 5466 8334 5468
rect 8038 5414 8084 5466
rect 8084 5414 8094 5466
rect 8118 5414 8148 5466
rect 8148 5414 8160 5466
rect 8160 5414 8174 5466
rect 8198 5414 8212 5466
rect 8212 5414 8224 5466
rect 8224 5414 8254 5466
rect 8278 5414 8288 5466
rect 8288 5414 8334 5466
rect 8038 5412 8094 5414
rect 8118 5412 8174 5414
rect 8198 5412 8254 5414
rect 8278 5412 8334 5414
rect 9034 8508 9036 8528
rect 9036 8508 9088 8528
rect 9088 8508 9090 8528
rect 9034 8472 9090 8508
rect 9770 9288 9826 9344
rect 10414 12144 10470 12200
rect 11580 16890 11636 16892
rect 11660 16890 11716 16892
rect 11740 16890 11796 16892
rect 11820 16890 11876 16892
rect 11580 16838 11626 16890
rect 11626 16838 11636 16890
rect 11660 16838 11690 16890
rect 11690 16838 11702 16890
rect 11702 16838 11716 16890
rect 11740 16838 11754 16890
rect 11754 16838 11766 16890
rect 11766 16838 11796 16890
rect 11820 16838 11830 16890
rect 11830 16838 11876 16890
rect 11580 16836 11636 16838
rect 11660 16836 11716 16838
rect 11740 16836 11796 16838
rect 11820 16836 11876 16838
rect 11580 15802 11636 15804
rect 11660 15802 11716 15804
rect 11740 15802 11796 15804
rect 11820 15802 11876 15804
rect 11580 15750 11626 15802
rect 11626 15750 11636 15802
rect 11660 15750 11690 15802
rect 11690 15750 11702 15802
rect 11702 15750 11716 15802
rect 11740 15750 11754 15802
rect 11754 15750 11766 15802
rect 11766 15750 11796 15802
rect 11820 15750 11830 15802
rect 11830 15750 11876 15802
rect 11580 15748 11636 15750
rect 11660 15748 11716 15750
rect 11740 15748 11796 15750
rect 11820 15748 11876 15750
rect 11580 14714 11636 14716
rect 11660 14714 11716 14716
rect 11740 14714 11796 14716
rect 11820 14714 11876 14716
rect 11580 14662 11626 14714
rect 11626 14662 11636 14714
rect 11660 14662 11690 14714
rect 11690 14662 11702 14714
rect 11702 14662 11716 14714
rect 11740 14662 11754 14714
rect 11754 14662 11766 14714
rect 11766 14662 11796 14714
rect 11820 14662 11830 14714
rect 11830 14662 11876 14714
rect 11580 14660 11636 14662
rect 11660 14660 11716 14662
rect 11740 14660 11796 14662
rect 11820 14660 11876 14662
rect 11580 13626 11636 13628
rect 11660 13626 11716 13628
rect 11740 13626 11796 13628
rect 11820 13626 11876 13628
rect 11580 13574 11626 13626
rect 11626 13574 11636 13626
rect 11660 13574 11690 13626
rect 11690 13574 11702 13626
rect 11702 13574 11716 13626
rect 11740 13574 11754 13626
rect 11754 13574 11766 13626
rect 11766 13574 11796 13626
rect 11820 13574 11830 13626
rect 11830 13574 11876 13626
rect 11580 13572 11636 13574
rect 11660 13572 11716 13574
rect 11740 13572 11796 13574
rect 11820 13572 11876 13574
rect 11518 13232 11574 13288
rect 11580 12538 11636 12540
rect 11660 12538 11716 12540
rect 11740 12538 11796 12540
rect 11820 12538 11876 12540
rect 11580 12486 11626 12538
rect 11626 12486 11636 12538
rect 11660 12486 11690 12538
rect 11690 12486 11702 12538
rect 11702 12486 11716 12538
rect 11740 12486 11754 12538
rect 11754 12486 11766 12538
rect 11766 12486 11796 12538
rect 11820 12486 11830 12538
rect 11830 12486 11876 12538
rect 11580 12484 11636 12486
rect 11660 12484 11716 12486
rect 11740 12484 11796 12486
rect 11820 12484 11876 12486
rect 13910 20576 13966 20632
rect 22204 30490 22260 30492
rect 22284 30490 22340 30492
rect 22364 30490 22420 30492
rect 22444 30490 22500 30492
rect 22204 30438 22250 30490
rect 22250 30438 22260 30490
rect 22284 30438 22314 30490
rect 22314 30438 22326 30490
rect 22326 30438 22340 30490
rect 22364 30438 22378 30490
rect 22378 30438 22390 30490
rect 22390 30438 22420 30490
rect 22444 30438 22454 30490
rect 22454 30438 22500 30490
rect 22204 30436 22260 30438
rect 22284 30436 22340 30438
rect 22364 30436 22420 30438
rect 22444 30436 22500 30438
rect 28906 30640 28962 30696
rect 15121 29402 15177 29404
rect 15201 29402 15257 29404
rect 15281 29402 15337 29404
rect 15361 29402 15417 29404
rect 15121 29350 15167 29402
rect 15167 29350 15177 29402
rect 15201 29350 15231 29402
rect 15231 29350 15243 29402
rect 15243 29350 15257 29402
rect 15281 29350 15295 29402
rect 15295 29350 15307 29402
rect 15307 29350 15337 29402
rect 15361 29350 15371 29402
rect 15371 29350 15417 29402
rect 15121 29348 15177 29350
rect 15201 29348 15257 29350
rect 15281 29348 15337 29350
rect 15361 29348 15417 29350
rect 15121 28314 15177 28316
rect 15201 28314 15257 28316
rect 15281 28314 15337 28316
rect 15361 28314 15417 28316
rect 15121 28262 15167 28314
rect 15167 28262 15177 28314
rect 15201 28262 15231 28314
rect 15231 28262 15243 28314
rect 15243 28262 15257 28314
rect 15281 28262 15295 28314
rect 15295 28262 15307 28314
rect 15307 28262 15337 28314
rect 15361 28262 15371 28314
rect 15371 28262 15417 28314
rect 15121 28260 15177 28262
rect 15201 28260 15257 28262
rect 15281 28260 15337 28262
rect 15361 28260 15417 28262
rect 15121 27226 15177 27228
rect 15201 27226 15257 27228
rect 15281 27226 15337 27228
rect 15361 27226 15417 27228
rect 15121 27174 15167 27226
rect 15167 27174 15177 27226
rect 15201 27174 15231 27226
rect 15231 27174 15243 27226
rect 15243 27174 15257 27226
rect 15281 27174 15295 27226
rect 15295 27174 15307 27226
rect 15307 27174 15337 27226
rect 15361 27174 15371 27226
rect 15371 27174 15417 27226
rect 15121 27172 15177 27174
rect 15201 27172 15257 27174
rect 15281 27172 15337 27174
rect 15361 27172 15417 27174
rect 15121 26138 15177 26140
rect 15201 26138 15257 26140
rect 15281 26138 15337 26140
rect 15361 26138 15417 26140
rect 15121 26086 15167 26138
rect 15167 26086 15177 26138
rect 15201 26086 15231 26138
rect 15231 26086 15243 26138
rect 15243 26086 15257 26138
rect 15281 26086 15295 26138
rect 15295 26086 15307 26138
rect 15307 26086 15337 26138
rect 15361 26086 15371 26138
rect 15371 26086 15417 26138
rect 15121 26084 15177 26086
rect 15201 26084 15257 26086
rect 15281 26084 15337 26086
rect 15361 26084 15417 26086
rect 18663 29946 18719 29948
rect 18743 29946 18799 29948
rect 18823 29946 18879 29948
rect 18903 29946 18959 29948
rect 18663 29894 18709 29946
rect 18709 29894 18719 29946
rect 18743 29894 18773 29946
rect 18773 29894 18785 29946
rect 18785 29894 18799 29946
rect 18823 29894 18837 29946
rect 18837 29894 18849 29946
rect 18849 29894 18879 29946
rect 18903 29894 18913 29946
rect 18913 29894 18959 29946
rect 18663 29892 18719 29894
rect 18743 29892 18799 29894
rect 18823 29892 18879 29894
rect 18903 29892 18959 29894
rect 17958 28464 18014 28520
rect 18663 28858 18719 28860
rect 18743 28858 18799 28860
rect 18823 28858 18879 28860
rect 18903 28858 18959 28860
rect 18663 28806 18709 28858
rect 18709 28806 18719 28858
rect 18743 28806 18773 28858
rect 18773 28806 18785 28858
rect 18785 28806 18799 28858
rect 18823 28806 18837 28858
rect 18837 28806 18849 28858
rect 18849 28806 18879 28858
rect 18903 28806 18913 28858
rect 18913 28806 18959 28858
rect 18663 28804 18719 28806
rect 18743 28804 18799 28806
rect 18823 28804 18879 28806
rect 18903 28804 18959 28806
rect 18663 27770 18719 27772
rect 18743 27770 18799 27772
rect 18823 27770 18879 27772
rect 18903 27770 18959 27772
rect 18663 27718 18709 27770
rect 18709 27718 18719 27770
rect 18743 27718 18773 27770
rect 18773 27718 18785 27770
rect 18785 27718 18799 27770
rect 18823 27718 18837 27770
rect 18837 27718 18849 27770
rect 18849 27718 18879 27770
rect 18903 27718 18913 27770
rect 18913 27718 18959 27770
rect 18663 27716 18719 27718
rect 18743 27716 18799 27718
rect 18823 27716 18879 27718
rect 18903 27716 18959 27718
rect 18663 26682 18719 26684
rect 18743 26682 18799 26684
rect 18823 26682 18879 26684
rect 18903 26682 18959 26684
rect 18663 26630 18709 26682
rect 18709 26630 18719 26682
rect 18743 26630 18773 26682
rect 18773 26630 18785 26682
rect 18785 26630 18799 26682
rect 18823 26630 18837 26682
rect 18837 26630 18849 26682
rect 18849 26630 18879 26682
rect 18903 26630 18913 26682
rect 18913 26630 18959 26682
rect 18663 26628 18719 26630
rect 18743 26628 18799 26630
rect 18823 26628 18879 26630
rect 18903 26628 18959 26630
rect 15121 25050 15177 25052
rect 15201 25050 15257 25052
rect 15281 25050 15337 25052
rect 15361 25050 15417 25052
rect 15121 24998 15167 25050
rect 15167 24998 15177 25050
rect 15201 24998 15231 25050
rect 15231 24998 15243 25050
rect 15243 24998 15257 25050
rect 15281 24998 15295 25050
rect 15295 24998 15307 25050
rect 15307 24998 15337 25050
rect 15361 24998 15371 25050
rect 15371 24998 15417 25050
rect 15121 24996 15177 24998
rect 15201 24996 15257 24998
rect 15281 24996 15337 24998
rect 15361 24996 15417 24998
rect 15121 23962 15177 23964
rect 15201 23962 15257 23964
rect 15281 23962 15337 23964
rect 15361 23962 15417 23964
rect 15121 23910 15167 23962
rect 15167 23910 15177 23962
rect 15201 23910 15231 23962
rect 15231 23910 15243 23962
rect 15243 23910 15257 23962
rect 15281 23910 15295 23962
rect 15295 23910 15307 23962
rect 15307 23910 15337 23962
rect 15361 23910 15371 23962
rect 15371 23910 15417 23962
rect 15121 23908 15177 23910
rect 15201 23908 15257 23910
rect 15281 23908 15337 23910
rect 15361 23908 15417 23910
rect 15121 22874 15177 22876
rect 15201 22874 15257 22876
rect 15281 22874 15337 22876
rect 15361 22874 15417 22876
rect 15121 22822 15167 22874
rect 15167 22822 15177 22874
rect 15201 22822 15231 22874
rect 15231 22822 15243 22874
rect 15243 22822 15257 22874
rect 15281 22822 15295 22874
rect 15295 22822 15307 22874
rect 15307 22822 15337 22874
rect 15361 22822 15371 22874
rect 15371 22822 15417 22874
rect 15121 22820 15177 22822
rect 15201 22820 15257 22822
rect 15281 22820 15337 22822
rect 15361 22820 15417 22822
rect 14278 19760 14334 19816
rect 15121 21786 15177 21788
rect 15201 21786 15257 21788
rect 15281 21786 15337 21788
rect 15361 21786 15417 21788
rect 15121 21734 15167 21786
rect 15167 21734 15177 21786
rect 15201 21734 15231 21786
rect 15231 21734 15243 21786
rect 15243 21734 15257 21786
rect 15281 21734 15295 21786
rect 15295 21734 15307 21786
rect 15307 21734 15337 21786
rect 15361 21734 15371 21786
rect 15371 21734 15417 21786
rect 15121 21732 15177 21734
rect 15201 21732 15257 21734
rect 15281 21732 15337 21734
rect 15361 21732 15417 21734
rect 15121 20698 15177 20700
rect 15201 20698 15257 20700
rect 15281 20698 15337 20700
rect 15361 20698 15417 20700
rect 15121 20646 15167 20698
rect 15167 20646 15177 20698
rect 15201 20646 15231 20698
rect 15231 20646 15243 20698
rect 15243 20646 15257 20698
rect 15281 20646 15295 20698
rect 15295 20646 15307 20698
rect 15307 20646 15337 20698
rect 15361 20646 15371 20698
rect 15371 20646 15417 20698
rect 15121 20644 15177 20646
rect 15201 20644 15257 20646
rect 15281 20644 15337 20646
rect 15361 20644 15417 20646
rect 15121 19610 15177 19612
rect 15201 19610 15257 19612
rect 15281 19610 15337 19612
rect 15361 19610 15417 19612
rect 15121 19558 15167 19610
rect 15167 19558 15177 19610
rect 15201 19558 15231 19610
rect 15231 19558 15243 19610
rect 15243 19558 15257 19610
rect 15281 19558 15295 19610
rect 15295 19558 15307 19610
rect 15307 19558 15337 19610
rect 15361 19558 15371 19610
rect 15371 19558 15417 19610
rect 15121 19556 15177 19558
rect 15201 19556 15257 19558
rect 15281 19556 15337 19558
rect 15361 19556 15417 19558
rect 14922 19352 14978 19408
rect 15934 20848 15990 20904
rect 12346 13912 12402 13968
rect 11580 11450 11636 11452
rect 11660 11450 11716 11452
rect 11740 11450 11796 11452
rect 11820 11450 11876 11452
rect 11580 11398 11626 11450
rect 11626 11398 11636 11450
rect 11660 11398 11690 11450
rect 11690 11398 11702 11450
rect 11702 11398 11716 11450
rect 11740 11398 11754 11450
rect 11754 11398 11766 11450
rect 11766 11398 11796 11450
rect 11820 11398 11830 11450
rect 11830 11398 11876 11450
rect 11580 11396 11636 11398
rect 11660 11396 11716 11398
rect 11740 11396 11796 11398
rect 11820 11396 11876 11398
rect 10322 9696 10378 9752
rect 10322 9288 10378 9344
rect 10874 9696 10930 9752
rect 11580 10362 11636 10364
rect 11660 10362 11716 10364
rect 11740 10362 11796 10364
rect 11820 10362 11876 10364
rect 11580 10310 11626 10362
rect 11626 10310 11636 10362
rect 11660 10310 11690 10362
rect 11690 10310 11702 10362
rect 11702 10310 11716 10362
rect 11740 10310 11754 10362
rect 11754 10310 11766 10362
rect 11766 10310 11796 10362
rect 11820 10310 11830 10362
rect 11830 10310 11876 10362
rect 11580 10308 11636 10310
rect 11660 10308 11716 10310
rect 11740 10308 11796 10310
rect 11820 10308 11876 10310
rect 11150 9696 11206 9752
rect 10506 8200 10562 8256
rect 11580 9274 11636 9276
rect 11660 9274 11716 9276
rect 11740 9274 11796 9276
rect 11820 9274 11876 9276
rect 11580 9222 11626 9274
rect 11626 9222 11636 9274
rect 11660 9222 11690 9274
rect 11690 9222 11702 9274
rect 11702 9222 11716 9274
rect 11740 9222 11754 9274
rect 11754 9222 11766 9274
rect 11766 9222 11796 9274
rect 11820 9222 11830 9274
rect 11830 9222 11876 9274
rect 11580 9220 11636 9222
rect 11660 9220 11716 9222
rect 11740 9220 11796 9222
rect 11820 9220 11876 9222
rect 13266 11056 13322 11112
rect 12254 9560 12310 9616
rect 11580 8186 11636 8188
rect 11660 8186 11716 8188
rect 11740 8186 11796 8188
rect 11820 8186 11876 8188
rect 11580 8134 11626 8186
rect 11626 8134 11636 8186
rect 11660 8134 11690 8186
rect 11690 8134 11702 8186
rect 11702 8134 11716 8186
rect 11740 8134 11754 8186
rect 11754 8134 11766 8186
rect 11766 8134 11796 8186
rect 11820 8134 11830 8186
rect 11830 8134 11876 8186
rect 11580 8132 11636 8134
rect 11660 8132 11716 8134
rect 11740 8132 11796 8134
rect 11820 8132 11876 8134
rect 11580 7098 11636 7100
rect 11660 7098 11716 7100
rect 11740 7098 11796 7100
rect 11820 7098 11876 7100
rect 11580 7046 11626 7098
rect 11626 7046 11636 7098
rect 11660 7046 11690 7098
rect 11690 7046 11702 7098
rect 11702 7046 11716 7098
rect 11740 7046 11754 7098
rect 11754 7046 11766 7098
rect 11766 7046 11796 7098
rect 11820 7046 11830 7098
rect 11830 7046 11876 7098
rect 11580 7044 11636 7046
rect 11660 7044 11716 7046
rect 11740 7044 11796 7046
rect 11820 7044 11876 7046
rect 10782 6704 10838 6760
rect 10966 6568 11022 6624
rect 11580 6010 11636 6012
rect 11660 6010 11716 6012
rect 11740 6010 11796 6012
rect 11820 6010 11876 6012
rect 11580 5958 11626 6010
rect 11626 5958 11636 6010
rect 11660 5958 11690 6010
rect 11690 5958 11702 6010
rect 11702 5958 11716 6010
rect 11740 5958 11754 6010
rect 11754 5958 11766 6010
rect 11766 5958 11796 6010
rect 11820 5958 11830 6010
rect 11830 5958 11876 6010
rect 11580 5956 11636 5958
rect 11660 5956 11716 5958
rect 11740 5956 11796 5958
rect 11820 5956 11876 5958
rect 13174 9596 13176 9616
rect 13176 9596 13228 9616
rect 13228 9596 13230 9616
rect 13174 9560 13230 9596
rect 14094 12144 14150 12200
rect 15121 18522 15177 18524
rect 15201 18522 15257 18524
rect 15281 18522 15337 18524
rect 15361 18522 15417 18524
rect 15121 18470 15167 18522
rect 15167 18470 15177 18522
rect 15201 18470 15231 18522
rect 15231 18470 15243 18522
rect 15243 18470 15257 18522
rect 15281 18470 15295 18522
rect 15295 18470 15307 18522
rect 15307 18470 15337 18522
rect 15361 18470 15371 18522
rect 15371 18470 15417 18522
rect 15121 18468 15177 18470
rect 15201 18468 15257 18470
rect 15281 18468 15337 18470
rect 15361 18468 15417 18470
rect 15198 17856 15254 17912
rect 15121 17434 15177 17436
rect 15201 17434 15257 17436
rect 15281 17434 15337 17436
rect 15361 17434 15417 17436
rect 15121 17382 15167 17434
rect 15167 17382 15177 17434
rect 15201 17382 15231 17434
rect 15231 17382 15243 17434
rect 15243 17382 15257 17434
rect 15281 17382 15295 17434
rect 15295 17382 15307 17434
rect 15307 17382 15337 17434
rect 15361 17382 15371 17434
rect 15371 17382 15417 17434
rect 15121 17380 15177 17382
rect 15201 17380 15257 17382
rect 15281 17380 15337 17382
rect 15361 17380 15417 17382
rect 14278 12280 14334 12336
rect 13910 6568 13966 6624
rect 14094 6704 14150 6760
rect 15121 16346 15177 16348
rect 15201 16346 15257 16348
rect 15281 16346 15337 16348
rect 15361 16346 15417 16348
rect 15121 16294 15167 16346
rect 15167 16294 15177 16346
rect 15201 16294 15231 16346
rect 15231 16294 15243 16346
rect 15243 16294 15257 16346
rect 15281 16294 15295 16346
rect 15295 16294 15307 16346
rect 15307 16294 15337 16346
rect 15361 16294 15371 16346
rect 15371 16294 15417 16346
rect 15121 16292 15177 16294
rect 15201 16292 15257 16294
rect 15281 16292 15337 16294
rect 15361 16292 15417 16294
rect 15121 15258 15177 15260
rect 15201 15258 15257 15260
rect 15281 15258 15337 15260
rect 15361 15258 15417 15260
rect 15121 15206 15167 15258
rect 15167 15206 15177 15258
rect 15201 15206 15231 15258
rect 15231 15206 15243 15258
rect 15243 15206 15257 15258
rect 15281 15206 15295 15258
rect 15295 15206 15307 15258
rect 15307 15206 15337 15258
rect 15361 15206 15371 15258
rect 15371 15206 15417 15258
rect 15121 15204 15177 15206
rect 15201 15204 15257 15206
rect 15281 15204 15337 15206
rect 15361 15204 15417 15206
rect 15121 14170 15177 14172
rect 15201 14170 15257 14172
rect 15281 14170 15337 14172
rect 15361 14170 15417 14172
rect 15121 14118 15167 14170
rect 15167 14118 15177 14170
rect 15201 14118 15231 14170
rect 15231 14118 15243 14170
rect 15243 14118 15257 14170
rect 15281 14118 15295 14170
rect 15295 14118 15307 14170
rect 15307 14118 15337 14170
rect 15361 14118 15371 14170
rect 15371 14118 15417 14170
rect 15121 14116 15177 14118
rect 15201 14116 15257 14118
rect 15281 14116 15337 14118
rect 15361 14116 15417 14118
rect 15121 13082 15177 13084
rect 15201 13082 15257 13084
rect 15281 13082 15337 13084
rect 15361 13082 15417 13084
rect 15121 13030 15167 13082
rect 15167 13030 15177 13082
rect 15201 13030 15231 13082
rect 15231 13030 15243 13082
rect 15243 13030 15257 13082
rect 15281 13030 15295 13082
rect 15295 13030 15307 13082
rect 15307 13030 15337 13082
rect 15361 13030 15371 13082
rect 15371 13030 15417 13082
rect 15121 13028 15177 13030
rect 15201 13028 15257 13030
rect 15281 13028 15337 13030
rect 15361 13028 15417 13030
rect 15121 11994 15177 11996
rect 15201 11994 15257 11996
rect 15281 11994 15337 11996
rect 15361 11994 15417 11996
rect 15121 11942 15167 11994
rect 15167 11942 15177 11994
rect 15201 11942 15231 11994
rect 15231 11942 15243 11994
rect 15243 11942 15257 11994
rect 15281 11942 15295 11994
rect 15295 11942 15307 11994
rect 15307 11942 15337 11994
rect 15361 11942 15371 11994
rect 15371 11942 15417 11994
rect 15121 11940 15177 11942
rect 15201 11940 15257 11942
rect 15281 11940 15337 11942
rect 15361 11940 15417 11942
rect 15121 10906 15177 10908
rect 15201 10906 15257 10908
rect 15281 10906 15337 10908
rect 15361 10906 15417 10908
rect 15121 10854 15167 10906
rect 15167 10854 15177 10906
rect 15201 10854 15231 10906
rect 15231 10854 15243 10906
rect 15243 10854 15257 10906
rect 15281 10854 15295 10906
rect 15295 10854 15307 10906
rect 15307 10854 15337 10906
rect 15361 10854 15371 10906
rect 15371 10854 15417 10906
rect 15121 10852 15177 10854
rect 15201 10852 15257 10854
rect 15281 10852 15337 10854
rect 15361 10852 15417 10854
rect 15121 9818 15177 9820
rect 15201 9818 15257 9820
rect 15281 9818 15337 9820
rect 15361 9818 15417 9820
rect 15121 9766 15167 9818
rect 15167 9766 15177 9818
rect 15201 9766 15231 9818
rect 15231 9766 15243 9818
rect 15243 9766 15257 9818
rect 15281 9766 15295 9818
rect 15295 9766 15307 9818
rect 15307 9766 15337 9818
rect 15361 9766 15371 9818
rect 15371 9766 15417 9818
rect 15121 9764 15177 9766
rect 15201 9764 15257 9766
rect 15281 9764 15337 9766
rect 15361 9764 15417 9766
rect 15121 8730 15177 8732
rect 15201 8730 15257 8732
rect 15281 8730 15337 8732
rect 15361 8730 15417 8732
rect 15121 8678 15167 8730
rect 15167 8678 15177 8730
rect 15201 8678 15231 8730
rect 15231 8678 15243 8730
rect 15243 8678 15257 8730
rect 15281 8678 15295 8730
rect 15295 8678 15307 8730
rect 15307 8678 15337 8730
rect 15361 8678 15371 8730
rect 15371 8678 15417 8730
rect 15121 8676 15177 8678
rect 15201 8676 15257 8678
rect 15281 8676 15337 8678
rect 15361 8676 15417 8678
rect 15121 7642 15177 7644
rect 15201 7642 15257 7644
rect 15281 7642 15337 7644
rect 15361 7642 15417 7644
rect 15121 7590 15167 7642
rect 15167 7590 15177 7642
rect 15201 7590 15231 7642
rect 15231 7590 15243 7642
rect 15243 7590 15257 7642
rect 15281 7590 15295 7642
rect 15295 7590 15307 7642
rect 15307 7590 15337 7642
rect 15361 7590 15371 7642
rect 15371 7590 15417 7642
rect 15121 7588 15177 7590
rect 15201 7588 15257 7590
rect 15281 7588 15337 7590
rect 15361 7588 15417 7590
rect 15121 6554 15177 6556
rect 15201 6554 15257 6556
rect 15281 6554 15337 6556
rect 15361 6554 15417 6556
rect 15121 6502 15167 6554
rect 15167 6502 15177 6554
rect 15201 6502 15231 6554
rect 15231 6502 15243 6554
rect 15243 6502 15257 6554
rect 15281 6502 15295 6554
rect 15295 6502 15307 6554
rect 15307 6502 15337 6554
rect 15361 6502 15371 6554
rect 15371 6502 15417 6554
rect 15121 6500 15177 6502
rect 15201 6500 15257 6502
rect 15281 6500 15337 6502
rect 15361 6500 15417 6502
rect 15121 5466 15177 5468
rect 15201 5466 15257 5468
rect 15281 5466 15337 5468
rect 15361 5466 15417 5468
rect 15121 5414 15167 5466
rect 15167 5414 15177 5466
rect 15201 5414 15231 5466
rect 15231 5414 15243 5466
rect 15243 5414 15257 5466
rect 15281 5414 15295 5466
rect 15295 5414 15307 5466
rect 15307 5414 15337 5466
rect 15361 5414 15371 5466
rect 15371 5414 15417 5466
rect 15121 5412 15177 5414
rect 15201 5412 15257 5414
rect 15281 5412 15337 5414
rect 15361 5412 15417 5414
rect 11580 4922 11636 4924
rect 11660 4922 11716 4924
rect 11740 4922 11796 4924
rect 11820 4922 11876 4924
rect 11580 4870 11626 4922
rect 11626 4870 11636 4922
rect 11660 4870 11690 4922
rect 11690 4870 11702 4922
rect 11702 4870 11716 4922
rect 11740 4870 11754 4922
rect 11754 4870 11766 4922
rect 11766 4870 11796 4922
rect 11820 4870 11830 4922
rect 11830 4870 11876 4922
rect 11580 4868 11636 4870
rect 11660 4868 11716 4870
rect 11740 4868 11796 4870
rect 11820 4868 11876 4870
rect 8038 4378 8094 4380
rect 8118 4378 8174 4380
rect 8198 4378 8254 4380
rect 8278 4378 8334 4380
rect 8038 4326 8084 4378
rect 8084 4326 8094 4378
rect 8118 4326 8148 4378
rect 8148 4326 8160 4378
rect 8160 4326 8174 4378
rect 8198 4326 8212 4378
rect 8212 4326 8224 4378
rect 8224 4326 8254 4378
rect 8278 4326 8288 4378
rect 8288 4326 8334 4378
rect 8038 4324 8094 4326
rect 8118 4324 8174 4326
rect 8198 4324 8254 4326
rect 8278 4324 8334 4326
rect 4497 3834 4553 3836
rect 4577 3834 4633 3836
rect 4657 3834 4713 3836
rect 4737 3834 4793 3836
rect 4497 3782 4543 3834
rect 4543 3782 4553 3834
rect 4577 3782 4607 3834
rect 4607 3782 4619 3834
rect 4619 3782 4633 3834
rect 4657 3782 4671 3834
rect 4671 3782 4683 3834
rect 4683 3782 4713 3834
rect 4737 3782 4747 3834
rect 4747 3782 4793 3834
rect 4497 3780 4553 3782
rect 4577 3780 4633 3782
rect 4657 3780 4713 3782
rect 4737 3780 4793 3782
rect 11580 3834 11636 3836
rect 11660 3834 11716 3836
rect 11740 3834 11796 3836
rect 11820 3834 11876 3836
rect 11580 3782 11626 3834
rect 11626 3782 11636 3834
rect 11660 3782 11690 3834
rect 11690 3782 11702 3834
rect 11702 3782 11716 3834
rect 11740 3782 11754 3834
rect 11754 3782 11766 3834
rect 11766 3782 11796 3834
rect 11820 3782 11830 3834
rect 11830 3782 11876 3834
rect 11580 3780 11636 3782
rect 11660 3780 11716 3782
rect 11740 3780 11796 3782
rect 11820 3780 11876 3782
rect 938 3440 994 3496
rect 8038 3290 8094 3292
rect 8118 3290 8174 3292
rect 8198 3290 8254 3292
rect 8278 3290 8334 3292
rect 8038 3238 8084 3290
rect 8084 3238 8094 3290
rect 8118 3238 8148 3290
rect 8148 3238 8160 3290
rect 8160 3238 8174 3290
rect 8198 3238 8212 3290
rect 8212 3238 8224 3290
rect 8224 3238 8254 3290
rect 8278 3238 8288 3290
rect 8288 3238 8334 3290
rect 8038 3236 8094 3238
rect 8118 3236 8174 3238
rect 8198 3236 8254 3238
rect 8278 3236 8334 3238
rect 4497 2746 4553 2748
rect 4577 2746 4633 2748
rect 4657 2746 4713 2748
rect 4737 2746 4793 2748
rect 4497 2694 4543 2746
rect 4543 2694 4553 2746
rect 4577 2694 4607 2746
rect 4607 2694 4619 2746
rect 4619 2694 4633 2746
rect 4657 2694 4671 2746
rect 4671 2694 4683 2746
rect 4683 2694 4713 2746
rect 4737 2694 4747 2746
rect 4747 2694 4793 2746
rect 4497 2692 4553 2694
rect 4577 2692 4633 2694
rect 4657 2692 4713 2694
rect 4737 2692 4793 2694
rect 11580 2746 11636 2748
rect 11660 2746 11716 2748
rect 11740 2746 11796 2748
rect 11820 2746 11876 2748
rect 11580 2694 11626 2746
rect 11626 2694 11636 2746
rect 11660 2694 11690 2746
rect 11690 2694 11702 2746
rect 11702 2694 11716 2746
rect 11740 2694 11754 2746
rect 11754 2694 11766 2746
rect 11766 2694 11796 2746
rect 11820 2694 11830 2746
rect 11830 2694 11876 2746
rect 11580 2692 11636 2694
rect 11660 2692 11716 2694
rect 11740 2692 11796 2694
rect 11820 2692 11876 2694
rect 13174 3460 13230 3496
rect 13174 3440 13176 3460
rect 13176 3440 13228 3460
rect 13228 3440 13230 3460
rect 15121 4378 15177 4380
rect 15201 4378 15257 4380
rect 15281 4378 15337 4380
rect 15361 4378 15417 4380
rect 15121 4326 15167 4378
rect 15167 4326 15177 4378
rect 15201 4326 15231 4378
rect 15231 4326 15243 4378
rect 15243 4326 15257 4378
rect 15281 4326 15295 4378
rect 15295 4326 15307 4378
rect 15307 4326 15337 4378
rect 15361 4326 15371 4378
rect 15371 4326 15417 4378
rect 15121 4324 15177 4326
rect 15201 4324 15257 4326
rect 15281 4324 15337 4326
rect 15361 4324 15417 4326
rect 16302 20712 16358 20768
rect 16302 15136 16358 15192
rect 19338 28056 19394 28112
rect 22204 29402 22260 29404
rect 22284 29402 22340 29404
rect 22364 29402 22420 29404
rect 22444 29402 22500 29404
rect 22204 29350 22250 29402
rect 22250 29350 22260 29402
rect 22284 29350 22314 29402
rect 22314 29350 22326 29402
rect 22326 29350 22340 29402
rect 22364 29350 22378 29402
rect 22378 29350 22390 29402
rect 22390 29350 22420 29402
rect 22444 29350 22454 29402
rect 22454 29350 22500 29402
rect 22204 29348 22260 29350
rect 22284 29348 22340 29350
rect 22364 29348 22420 29350
rect 22444 29348 22500 29350
rect 18663 25594 18719 25596
rect 18743 25594 18799 25596
rect 18823 25594 18879 25596
rect 18903 25594 18959 25596
rect 18663 25542 18709 25594
rect 18709 25542 18719 25594
rect 18743 25542 18773 25594
rect 18773 25542 18785 25594
rect 18785 25542 18799 25594
rect 18823 25542 18837 25594
rect 18837 25542 18849 25594
rect 18849 25542 18879 25594
rect 18903 25542 18913 25594
rect 18913 25542 18959 25594
rect 18663 25540 18719 25542
rect 18743 25540 18799 25542
rect 18823 25540 18879 25542
rect 18903 25540 18959 25542
rect 18663 24506 18719 24508
rect 18743 24506 18799 24508
rect 18823 24506 18879 24508
rect 18903 24506 18959 24508
rect 18663 24454 18709 24506
rect 18709 24454 18719 24506
rect 18743 24454 18773 24506
rect 18773 24454 18785 24506
rect 18785 24454 18799 24506
rect 18823 24454 18837 24506
rect 18837 24454 18849 24506
rect 18849 24454 18879 24506
rect 18903 24454 18913 24506
rect 18913 24454 18959 24506
rect 18663 24452 18719 24454
rect 18743 24452 18799 24454
rect 18823 24452 18879 24454
rect 18903 24452 18959 24454
rect 18663 23418 18719 23420
rect 18743 23418 18799 23420
rect 18823 23418 18879 23420
rect 18903 23418 18959 23420
rect 18663 23366 18709 23418
rect 18709 23366 18719 23418
rect 18743 23366 18773 23418
rect 18773 23366 18785 23418
rect 18785 23366 18799 23418
rect 18823 23366 18837 23418
rect 18837 23366 18849 23418
rect 18849 23366 18879 23418
rect 18903 23366 18913 23418
rect 18913 23366 18959 23418
rect 18663 23364 18719 23366
rect 18743 23364 18799 23366
rect 18823 23364 18879 23366
rect 18903 23364 18959 23366
rect 18663 22330 18719 22332
rect 18743 22330 18799 22332
rect 18823 22330 18879 22332
rect 18903 22330 18959 22332
rect 18663 22278 18709 22330
rect 18709 22278 18719 22330
rect 18743 22278 18773 22330
rect 18773 22278 18785 22330
rect 18785 22278 18799 22330
rect 18823 22278 18837 22330
rect 18837 22278 18849 22330
rect 18849 22278 18879 22330
rect 18903 22278 18913 22330
rect 18913 22278 18959 22330
rect 18663 22276 18719 22278
rect 18743 22276 18799 22278
rect 18823 22276 18879 22278
rect 18903 22276 18959 22278
rect 22006 28600 22062 28656
rect 21270 27956 21272 27976
rect 21272 27956 21324 27976
rect 21324 27956 21326 27976
rect 21270 27920 21326 27956
rect 22204 28314 22260 28316
rect 22284 28314 22340 28316
rect 22364 28314 22420 28316
rect 22444 28314 22500 28316
rect 22204 28262 22250 28314
rect 22250 28262 22260 28314
rect 22284 28262 22314 28314
rect 22314 28262 22326 28314
rect 22326 28262 22340 28314
rect 22364 28262 22378 28314
rect 22378 28262 22390 28314
rect 22390 28262 22420 28314
rect 22444 28262 22454 28314
rect 22454 28262 22500 28314
rect 22204 28260 22260 28262
rect 22284 28260 22340 28262
rect 22364 28260 22420 28262
rect 22444 28260 22500 28262
rect 22204 27226 22260 27228
rect 22284 27226 22340 27228
rect 22364 27226 22420 27228
rect 22444 27226 22500 27228
rect 22204 27174 22250 27226
rect 22250 27174 22260 27226
rect 22284 27174 22314 27226
rect 22314 27174 22326 27226
rect 22326 27174 22340 27226
rect 22364 27174 22378 27226
rect 22378 27174 22390 27226
rect 22390 27174 22420 27226
rect 22444 27174 22454 27226
rect 22454 27174 22500 27226
rect 22204 27172 22260 27174
rect 22284 27172 22340 27174
rect 22364 27172 22420 27174
rect 22444 27172 22500 27174
rect 22204 26138 22260 26140
rect 22284 26138 22340 26140
rect 22364 26138 22420 26140
rect 22444 26138 22500 26140
rect 22204 26086 22250 26138
rect 22250 26086 22260 26138
rect 22284 26086 22314 26138
rect 22314 26086 22326 26138
rect 22326 26086 22340 26138
rect 22364 26086 22378 26138
rect 22378 26086 22390 26138
rect 22390 26086 22420 26138
rect 22444 26086 22454 26138
rect 22454 26086 22500 26138
rect 22204 26084 22260 26086
rect 22284 26084 22340 26086
rect 22364 26084 22420 26086
rect 22444 26084 22500 26086
rect 22204 25050 22260 25052
rect 22284 25050 22340 25052
rect 22364 25050 22420 25052
rect 22444 25050 22500 25052
rect 22204 24998 22250 25050
rect 22250 24998 22260 25050
rect 22284 24998 22314 25050
rect 22314 24998 22326 25050
rect 22326 24998 22340 25050
rect 22364 24998 22378 25050
rect 22378 24998 22390 25050
rect 22390 24998 22420 25050
rect 22444 24998 22454 25050
rect 22454 24998 22500 25050
rect 22204 24996 22260 24998
rect 22284 24996 22340 24998
rect 22364 24996 22420 24998
rect 22444 24996 22500 24998
rect 17682 21936 17738 21992
rect 16946 19896 17002 19952
rect 18663 21242 18719 21244
rect 18743 21242 18799 21244
rect 18823 21242 18879 21244
rect 18903 21242 18959 21244
rect 18663 21190 18709 21242
rect 18709 21190 18719 21242
rect 18743 21190 18773 21242
rect 18773 21190 18785 21242
rect 18785 21190 18799 21242
rect 18823 21190 18837 21242
rect 18837 21190 18849 21242
rect 18849 21190 18879 21242
rect 18903 21190 18913 21242
rect 18913 21190 18959 21242
rect 18663 21188 18719 21190
rect 18743 21188 18799 21190
rect 18823 21188 18879 21190
rect 18903 21188 18959 21190
rect 18663 20154 18719 20156
rect 18743 20154 18799 20156
rect 18823 20154 18879 20156
rect 18903 20154 18959 20156
rect 18663 20102 18709 20154
rect 18709 20102 18719 20154
rect 18743 20102 18773 20154
rect 18773 20102 18785 20154
rect 18785 20102 18799 20154
rect 18823 20102 18837 20154
rect 18837 20102 18849 20154
rect 18849 20102 18879 20154
rect 18903 20102 18913 20154
rect 18913 20102 18959 20154
rect 18663 20100 18719 20102
rect 18743 20100 18799 20102
rect 18823 20100 18879 20102
rect 18903 20100 18959 20102
rect 18663 19066 18719 19068
rect 18743 19066 18799 19068
rect 18823 19066 18879 19068
rect 18903 19066 18959 19068
rect 18663 19014 18709 19066
rect 18709 19014 18719 19066
rect 18743 19014 18773 19066
rect 18773 19014 18785 19066
rect 18785 19014 18799 19066
rect 18823 19014 18837 19066
rect 18837 19014 18849 19066
rect 18849 19014 18879 19066
rect 18903 19014 18913 19066
rect 18913 19014 18959 19066
rect 18663 19012 18719 19014
rect 18743 19012 18799 19014
rect 18823 19012 18879 19014
rect 18903 19012 18959 19014
rect 18418 17856 18474 17912
rect 18663 17978 18719 17980
rect 18743 17978 18799 17980
rect 18823 17978 18879 17980
rect 18903 17978 18959 17980
rect 18663 17926 18709 17978
rect 18709 17926 18719 17978
rect 18743 17926 18773 17978
rect 18773 17926 18785 17978
rect 18785 17926 18799 17978
rect 18823 17926 18837 17978
rect 18837 17926 18849 17978
rect 18849 17926 18879 17978
rect 18903 17926 18913 17978
rect 18913 17926 18959 17978
rect 18663 17924 18719 17926
rect 18743 17924 18799 17926
rect 18823 17924 18879 17926
rect 18903 17924 18959 17926
rect 22204 23962 22260 23964
rect 22284 23962 22340 23964
rect 22364 23962 22420 23964
rect 22444 23962 22500 23964
rect 22204 23910 22250 23962
rect 22250 23910 22260 23962
rect 22284 23910 22314 23962
rect 22314 23910 22326 23962
rect 22326 23910 22340 23962
rect 22364 23910 22378 23962
rect 22378 23910 22390 23962
rect 22390 23910 22420 23962
rect 22444 23910 22454 23962
rect 22454 23910 22500 23962
rect 22204 23908 22260 23910
rect 22284 23908 22340 23910
rect 22364 23908 22420 23910
rect 22444 23908 22500 23910
rect 21178 23044 21234 23080
rect 21178 23024 21180 23044
rect 21180 23024 21232 23044
rect 21232 23024 21234 23044
rect 20350 22108 20352 22128
rect 20352 22108 20404 22128
rect 20404 22108 20406 22128
rect 20350 22072 20406 22108
rect 22204 22874 22260 22876
rect 22284 22874 22340 22876
rect 22364 22874 22420 22876
rect 22444 22874 22500 22876
rect 22204 22822 22250 22874
rect 22250 22822 22260 22874
rect 22284 22822 22314 22874
rect 22314 22822 22326 22874
rect 22326 22822 22340 22874
rect 22364 22822 22378 22874
rect 22378 22822 22390 22874
rect 22390 22822 22420 22874
rect 22444 22822 22454 22874
rect 22454 22822 22500 22874
rect 22204 22820 22260 22822
rect 22284 22820 22340 22822
rect 22364 22820 22420 22822
rect 22444 22820 22500 22822
rect 18663 16890 18719 16892
rect 18743 16890 18799 16892
rect 18823 16890 18879 16892
rect 18903 16890 18959 16892
rect 18663 16838 18709 16890
rect 18709 16838 18719 16890
rect 18743 16838 18773 16890
rect 18773 16838 18785 16890
rect 18785 16838 18799 16890
rect 18823 16838 18837 16890
rect 18837 16838 18849 16890
rect 18849 16838 18879 16890
rect 18903 16838 18913 16890
rect 18913 16838 18959 16890
rect 18663 16836 18719 16838
rect 18743 16836 18799 16838
rect 18823 16836 18879 16838
rect 18903 16836 18959 16838
rect 18663 15802 18719 15804
rect 18743 15802 18799 15804
rect 18823 15802 18879 15804
rect 18903 15802 18959 15804
rect 18663 15750 18709 15802
rect 18709 15750 18719 15802
rect 18743 15750 18773 15802
rect 18773 15750 18785 15802
rect 18785 15750 18799 15802
rect 18823 15750 18837 15802
rect 18837 15750 18849 15802
rect 18849 15750 18879 15802
rect 18903 15750 18913 15802
rect 18913 15750 18959 15802
rect 18663 15748 18719 15750
rect 18743 15748 18799 15750
rect 18823 15748 18879 15750
rect 18903 15748 18959 15750
rect 17958 15564 18014 15600
rect 17958 15544 17960 15564
rect 17960 15544 18012 15564
rect 18012 15544 18014 15564
rect 16670 12280 16726 12336
rect 16026 9560 16082 9616
rect 17038 9580 17094 9616
rect 18663 14714 18719 14716
rect 18743 14714 18799 14716
rect 18823 14714 18879 14716
rect 18903 14714 18959 14716
rect 18663 14662 18709 14714
rect 18709 14662 18719 14714
rect 18743 14662 18773 14714
rect 18773 14662 18785 14714
rect 18785 14662 18799 14714
rect 18823 14662 18837 14714
rect 18837 14662 18849 14714
rect 18849 14662 18879 14714
rect 18903 14662 18913 14714
rect 18913 14662 18959 14714
rect 18663 14660 18719 14662
rect 18743 14660 18799 14662
rect 18823 14660 18879 14662
rect 18903 14660 18959 14662
rect 17038 9560 17040 9580
rect 17040 9560 17092 9580
rect 17092 9560 17094 9580
rect 17130 9444 17186 9480
rect 17130 9424 17132 9444
rect 17132 9424 17184 9444
rect 17184 9424 17186 9444
rect 19430 17584 19486 17640
rect 20258 17720 20314 17776
rect 19062 13776 19118 13832
rect 18663 13626 18719 13628
rect 18743 13626 18799 13628
rect 18823 13626 18879 13628
rect 18903 13626 18959 13628
rect 18663 13574 18709 13626
rect 18709 13574 18719 13626
rect 18743 13574 18773 13626
rect 18773 13574 18785 13626
rect 18785 13574 18799 13626
rect 18823 13574 18837 13626
rect 18837 13574 18849 13626
rect 18849 13574 18879 13626
rect 18903 13574 18913 13626
rect 18913 13574 18959 13626
rect 18663 13572 18719 13574
rect 18743 13572 18799 13574
rect 18823 13572 18879 13574
rect 18903 13572 18959 13574
rect 18663 12538 18719 12540
rect 18743 12538 18799 12540
rect 18823 12538 18879 12540
rect 18903 12538 18959 12540
rect 18663 12486 18709 12538
rect 18709 12486 18719 12538
rect 18743 12486 18773 12538
rect 18773 12486 18785 12538
rect 18785 12486 18799 12538
rect 18823 12486 18837 12538
rect 18837 12486 18849 12538
rect 18849 12486 18879 12538
rect 18903 12486 18913 12538
rect 18913 12486 18959 12538
rect 18663 12484 18719 12486
rect 18743 12484 18799 12486
rect 18823 12484 18879 12486
rect 18903 12484 18959 12486
rect 19154 12280 19210 12336
rect 18663 11450 18719 11452
rect 18743 11450 18799 11452
rect 18823 11450 18879 11452
rect 18903 11450 18959 11452
rect 18663 11398 18709 11450
rect 18709 11398 18719 11450
rect 18743 11398 18773 11450
rect 18773 11398 18785 11450
rect 18785 11398 18799 11450
rect 18823 11398 18837 11450
rect 18837 11398 18849 11450
rect 18849 11398 18879 11450
rect 18903 11398 18913 11450
rect 18913 11398 18959 11450
rect 18663 11396 18719 11398
rect 18743 11396 18799 11398
rect 18823 11396 18879 11398
rect 18903 11396 18959 11398
rect 18694 11092 18696 11112
rect 18696 11092 18748 11112
rect 18748 11092 18750 11112
rect 18694 11056 18750 11092
rect 17406 7928 17462 7984
rect 17222 7384 17278 7440
rect 16210 4936 16266 4992
rect 15198 3440 15254 3496
rect 15121 3290 15177 3292
rect 15201 3290 15257 3292
rect 15281 3290 15337 3292
rect 15361 3290 15417 3292
rect 15121 3238 15167 3290
rect 15167 3238 15177 3290
rect 15201 3238 15231 3290
rect 15231 3238 15243 3290
rect 15243 3238 15257 3290
rect 15281 3238 15295 3290
rect 15295 3238 15307 3290
rect 15307 3238 15337 3290
rect 15361 3238 15371 3290
rect 15371 3238 15417 3290
rect 15121 3236 15177 3238
rect 15201 3236 15257 3238
rect 15281 3236 15337 3238
rect 15361 3236 15417 3238
rect 17866 7404 17922 7440
rect 18663 10362 18719 10364
rect 18743 10362 18799 10364
rect 18823 10362 18879 10364
rect 18903 10362 18959 10364
rect 18663 10310 18709 10362
rect 18709 10310 18719 10362
rect 18743 10310 18773 10362
rect 18773 10310 18785 10362
rect 18785 10310 18799 10362
rect 18823 10310 18837 10362
rect 18837 10310 18849 10362
rect 18849 10310 18879 10362
rect 18903 10310 18913 10362
rect 18913 10310 18959 10362
rect 18663 10308 18719 10310
rect 18743 10308 18799 10310
rect 18823 10308 18879 10310
rect 18903 10308 18959 10310
rect 18663 9274 18719 9276
rect 18743 9274 18799 9276
rect 18823 9274 18879 9276
rect 18903 9274 18959 9276
rect 18663 9222 18709 9274
rect 18709 9222 18719 9274
rect 18743 9222 18773 9274
rect 18773 9222 18785 9274
rect 18785 9222 18799 9274
rect 18823 9222 18837 9274
rect 18837 9222 18849 9274
rect 18849 9222 18879 9274
rect 18903 9222 18913 9274
rect 18913 9222 18959 9274
rect 18663 9220 18719 9222
rect 18743 9220 18799 9222
rect 18823 9220 18879 9222
rect 18903 9220 18959 9222
rect 20166 13776 20222 13832
rect 22204 21786 22260 21788
rect 22284 21786 22340 21788
rect 22364 21786 22420 21788
rect 22444 21786 22500 21788
rect 22204 21734 22250 21786
rect 22250 21734 22260 21786
rect 22284 21734 22314 21786
rect 22314 21734 22326 21786
rect 22326 21734 22340 21786
rect 22364 21734 22378 21786
rect 22378 21734 22390 21786
rect 22390 21734 22420 21786
rect 22444 21734 22454 21786
rect 22454 21734 22500 21786
rect 22204 21732 22260 21734
rect 22284 21732 22340 21734
rect 22364 21732 22420 21734
rect 22444 21732 22500 21734
rect 21822 21528 21878 21584
rect 22190 21120 22246 21176
rect 22204 20698 22260 20700
rect 22284 20698 22340 20700
rect 22364 20698 22420 20700
rect 22444 20698 22500 20700
rect 22204 20646 22250 20698
rect 22250 20646 22260 20698
rect 22284 20646 22314 20698
rect 22314 20646 22326 20698
rect 22326 20646 22340 20698
rect 22364 20646 22378 20698
rect 22378 20646 22390 20698
rect 22390 20646 22420 20698
rect 22444 20646 22454 20698
rect 22454 20646 22500 20698
rect 22204 20644 22260 20646
rect 22284 20644 22340 20646
rect 22364 20644 22420 20646
rect 22444 20644 22500 20646
rect 22204 19610 22260 19612
rect 22284 19610 22340 19612
rect 22364 19610 22420 19612
rect 22444 19610 22500 19612
rect 22204 19558 22250 19610
rect 22250 19558 22260 19610
rect 22284 19558 22314 19610
rect 22314 19558 22326 19610
rect 22326 19558 22340 19610
rect 22364 19558 22378 19610
rect 22378 19558 22390 19610
rect 22390 19558 22420 19610
rect 22444 19558 22454 19610
rect 22454 19558 22500 19610
rect 22204 19556 22260 19558
rect 22284 19556 22340 19558
rect 22364 19556 22420 19558
rect 22444 19556 22500 19558
rect 22204 18522 22260 18524
rect 22284 18522 22340 18524
rect 22364 18522 22420 18524
rect 22444 18522 22500 18524
rect 22204 18470 22250 18522
rect 22250 18470 22260 18522
rect 22284 18470 22314 18522
rect 22314 18470 22326 18522
rect 22326 18470 22340 18522
rect 22364 18470 22378 18522
rect 22378 18470 22390 18522
rect 22390 18470 22420 18522
rect 22444 18470 22454 18522
rect 22454 18470 22500 18522
rect 22204 18468 22260 18470
rect 22284 18468 22340 18470
rect 22364 18468 22420 18470
rect 22444 18468 22500 18470
rect 22926 21120 22982 21176
rect 23478 21120 23534 21176
rect 24398 22480 24454 22536
rect 22204 17434 22260 17436
rect 22284 17434 22340 17436
rect 22364 17434 22420 17436
rect 22444 17434 22500 17436
rect 22204 17382 22250 17434
rect 22250 17382 22260 17434
rect 22284 17382 22314 17434
rect 22314 17382 22326 17434
rect 22326 17382 22340 17434
rect 22364 17382 22378 17434
rect 22378 17382 22390 17434
rect 22390 17382 22420 17434
rect 22444 17382 22454 17434
rect 22454 17382 22500 17434
rect 22204 17380 22260 17382
rect 22284 17380 22340 17382
rect 22364 17380 22420 17382
rect 22444 17380 22500 17382
rect 22204 16346 22260 16348
rect 22284 16346 22340 16348
rect 22364 16346 22420 16348
rect 22444 16346 22500 16348
rect 22204 16294 22250 16346
rect 22250 16294 22260 16346
rect 22284 16294 22314 16346
rect 22314 16294 22326 16346
rect 22326 16294 22340 16346
rect 22364 16294 22378 16346
rect 22378 16294 22390 16346
rect 22390 16294 22420 16346
rect 22444 16294 22454 16346
rect 22454 16294 22500 16346
rect 22204 16292 22260 16294
rect 22284 16292 22340 16294
rect 22364 16292 22420 16294
rect 22444 16292 22500 16294
rect 22204 15258 22260 15260
rect 22284 15258 22340 15260
rect 22364 15258 22420 15260
rect 22444 15258 22500 15260
rect 22204 15206 22250 15258
rect 22250 15206 22260 15258
rect 22284 15206 22314 15258
rect 22314 15206 22326 15258
rect 22326 15206 22340 15258
rect 22364 15206 22378 15258
rect 22378 15206 22390 15258
rect 22390 15206 22420 15258
rect 22444 15206 22454 15258
rect 22454 15206 22500 15258
rect 22204 15204 22260 15206
rect 22284 15204 22340 15206
rect 22364 15204 22420 15206
rect 22444 15204 22500 15206
rect 19890 10104 19946 10160
rect 21546 11092 21548 11112
rect 21548 11092 21600 11112
rect 21600 11092 21602 11112
rect 21546 11056 21602 11092
rect 22204 14170 22260 14172
rect 22284 14170 22340 14172
rect 22364 14170 22420 14172
rect 22444 14170 22500 14172
rect 22204 14118 22250 14170
rect 22250 14118 22260 14170
rect 22284 14118 22314 14170
rect 22314 14118 22326 14170
rect 22326 14118 22340 14170
rect 22364 14118 22378 14170
rect 22378 14118 22390 14170
rect 22390 14118 22420 14170
rect 22444 14118 22454 14170
rect 22454 14118 22500 14170
rect 22204 14116 22260 14118
rect 22284 14116 22340 14118
rect 22364 14116 22420 14118
rect 22444 14116 22500 14118
rect 22204 13082 22260 13084
rect 22284 13082 22340 13084
rect 22364 13082 22420 13084
rect 22444 13082 22500 13084
rect 22204 13030 22250 13082
rect 22250 13030 22260 13082
rect 22284 13030 22314 13082
rect 22314 13030 22326 13082
rect 22326 13030 22340 13082
rect 22364 13030 22378 13082
rect 22378 13030 22390 13082
rect 22390 13030 22420 13082
rect 22444 13030 22454 13082
rect 22454 13030 22500 13082
rect 22204 13028 22260 13030
rect 22284 13028 22340 13030
rect 22364 13028 22420 13030
rect 22444 13028 22500 13030
rect 22204 11994 22260 11996
rect 22284 11994 22340 11996
rect 22364 11994 22420 11996
rect 22444 11994 22500 11996
rect 22204 11942 22250 11994
rect 22250 11942 22260 11994
rect 22284 11942 22314 11994
rect 22314 11942 22326 11994
rect 22326 11942 22340 11994
rect 22364 11942 22378 11994
rect 22378 11942 22390 11994
rect 22390 11942 22420 11994
rect 22444 11942 22454 11994
rect 22454 11942 22500 11994
rect 22204 11940 22260 11942
rect 22284 11940 22340 11942
rect 22364 11940 22420 11942
rect 22444 11940 22500 11942
rect 22204 10906 22260 10908
rect 22284 10906 22340 10908
rect 22364 10906 22420 10908
rect 22444 10906 22500 10908
rect 22204 10854 22250 10906
rect 22250 10854 22260 10906
rect 22284 10854 22314 10906
rect 22314 10854 22326 10906
rect 22326 10854 22340 10906
rect 22364 10854 22378 10906
rect 22378 10854 22390 10906
rect 22390 10854 22420 10906
rect 22444 10854 22454 10906
rect 22454 10854 22500 10906
rect 22204 10852 22260 10854
rect 22284 10852 22340 10854
rect 22364 10852 22420 10854
rect 22444 10852 22500 10854
rect 22834 12280 22890 12336
rect 22650 10104 22706 10160
rect 22204 9818 22260 9820
rect 22284 9818 22340 9820
rect 22364 9818 22420 9820
rect 22444 9818 22500 9820
rect 22204 9766 22250 9818
rect 22250 9766 22260 9818
rect 22284 9766 22314 9818
rect 22314 9766 22326 9818
rect 22326 9766 22340 9818
rect 22364 9766 22378 9818
rect 22378 9766 22390 9818
rect 22390 9766 22420 9818
rect 22444 9766 22454 9818
rect 22454 9766 22500 9818
rect 22204 9764 22260 9766
rect 22284 9764 22340 9766
rect 22364 9764 22420 9766
rect 22444 9764 22500 9766
rect 18663 8186 18719 8188
rect 18743 8186 18799 8188
rect 18823 8186 18879 8188
rect 18903 8186 18959 8188
rect 18663 8134 18709 8186
rect 18709 8134 18719 8186
rect 18743 8134 18773 8186
rect 18773 8134 18785 8186
rect 18785 8134 18799 8186
rect 18823 8134 18837 8186
rect 18837 8134 18849 8186
rect 18849 8134 18879 8186
rect 18903 8134 18913 8186
rect 18913 8134 18959 8186
rect 18663 8132 18719 8134
rect 18743 8132 18799 8134
rect 18823 8132 18879 8134
rect 18903 8132 18959 8134
rect 17866 7384 17868 7404
rect 17868 7384 17920 7404
rect 17920 7384 17922 7404
rect 17038 5072 17094 5128
rect 18663 7098 18719 7100
rect 18743 7098 18799 7100
rect 18823 7098 18879 7100
rect 18903 7098 18959 7100
rect 18663 7046 18709 7098
rect 18709 7046 18719 7098
rect 18743 7046 18773 7098
rect 18773 7046 18785 7098
rect 18785 7046 18799 7098
rect 18823 7046 18837 7098
rect 18837 7046 18849 7098
rect 18849 7046 18879 7098
rect 18903 7046 18913 7098
rect 18913 7046 18959 7098
rect 18663 7044 18719 7046
rect 18743 7044 18799 7046
rect 18823 7044 18879 7046
rect 18903 7044 18959 7046
rect 22204 8730 22260 8732
rect 22284 8730 22340 8732
rect 22364 8730 22420 8732
rect 22444 8730 22500 8732
rect 22204 8678 22250 8730
rect 22250 8678 22260 8730
rect 22284 8678 22314 8730
rect 22314 8678 22326 8730
rect 22326 8678 22340 8730
rect 22364 8678 22378 8730
rect 22378 8678 22390 8730
rect 22390 8678 22420 8730
rect 22444 8678 22454 8730
rect 22454 8678 22500 8730
rect 22204 8676 22260 8678
rect 22284 8676 22340 8678
rect 22364 8676 22420 8678
rect 22444 8676 22500 8678
rect 20074 6704 20130 6760
rect 22204 7642 22260 7644
rect 22284 7642 22340 7644
rect 22364 7642 22420 7644
rect 22444 7642 22500 7644
rect 22204 7590 22250 7642
rect 22250 7590 22260 7642
rect 22284 7590 22314 7642
rect 22314 7590 22326 7642
rect 22326 7590 22340 7642
rect 22364 7590 22378 7642
rect 22378 7590 22390 7642
rect 22390 7590 22420 7642
rect 22444 7590 22454 7642
rect 22454 7590 22500 7642
rect 22204 7588 22260 7590
rect 22284 7588 22340 7590
rect 22364 7588 22420 7590
rect 22444 7588 22500 7590
rect 22834 7928 22890 7984
rect 22204 6554 22260 6556
rect 22284 6554 22340 6556
rect 22364 6554 22420 6556
rect 22444 6554 22500 6556
rect 22204 6502 22250 6554
rect 22250 6502 22260 6554
rect 22284 6502 22314 6554
rect 22314 6502 22326 6554
rect 22326 6502 22340 6554
rect 22364 6502 22378 6554
rect 22378 6502 22390 6554
rect 22390 6502 22420 6554
rect 22444 6502 22454 6554
rect 22454 6502 22500 6554
rect 22204 6500 22260 6502
rect 22284 6500 22340 6502
rect 22364 6500 22420 6502
rect 22444 6500 22500 6502
rect 20258 6316 20314 6352
rect 20258 6296 20260 6316
rect 20260 6296 20312 6316
rect 20312 6296 20314 6316
rect 18663 6010 18719 6012
rect 18743 6010 18799 6012
rect 18823 6010 18879 6012
rect 18903 6010 18959 6012
rect 18663 5958 18709 6010
rect 18709 5958 18719 6010
rect 18743 5958 18773 6010
rect 18773 5958 18785 6010
rect 18785 5958 18799 6010
rect 18823 5958 18837 6010
rect 18837 5958 18849 6010
rect 18849 5958 18879 6010
rect 18903 5958 18913 6010
rect 18913 5958 18959 6010
rect 18663 5956 18719 5958
rect 18743 5956 18799 5958
rect 18823 5956 18879 5958
rect 18903 5956 18959 5958
rect 18234 5072 18290 5128
rect 18326 4936 18382 4992
rect 18663 4922 18719 4924
rect 18743 4922 18799 4924
rect 18823 4922 18879 4924
rect 18903 4922 18959 4924
rect 18663 4870 18709 4922
rect 18709 4870 18719 4922
rect 18743 4870 18773 4922
rect 18773 4870 18785 4922
rect 18785 4870 18799 4922
rect 18823 4870 18837 4922
rect 18837 4870 18849 4922
rect 18849 4870 18879 4922
rect 18903 4870 18913 4922
rect 18913 4870 18959 4922
rect 18663 4868 18719 4870
rect 18743 4868 18799 4870
rect 18823 4868 18879 4870
rect 18903 4868 18959 4870
rect 18663 3834 18719 3836
rect 18743 3834 18799 3836
rect 18823 3834 18879 3836
rect 18903 3834 18959 3836
rect 18663 3782 18709 3834
rect 18709 3782 18719 3834
rect 18743 3782 18773 3834
rect 18773 3782 18785 3834
rect 18785 3782 18799 3834
rect 18823 3782 18837 3834
rect 18837 3782 18849 3834
rect 18849 3782 18879 3834
rect 18903 3782 18913 3834
rect 18913 3782 18959 3834
rect 18663 3780 18719 3782
rect 18743 3780 18799 3782
rect 18823 3780 18879 3782
rect 18903 3780 18959 3782
rect 18663 2746 18719 2748
rect 18743 2746 18799 2748
rect 18823 2746 18879 2748
rect 18903 2746 18959 2748
rect 18663 2694 18709 2746
rect 18709 2694 18719 2746
rect 18743 2694 18773 2746
rect 18773 2694 18785 2746
rect 18785 2694 18799 2746
rect 18823 2694 18837 2746
rect 18837 2694 18849 2746
rect 18849 2694 18879 2746
rect 18903 2694 18913 2746
rect 18913 2694 18959 2746
rect 18663 2692 18719 2694
rect 18743 2692 18799 2694
rect 18823 2692 18879 2694
rect 18903 2692 18959 2694
rect 22204 5466 22260 5468
rect 22284 5466 22340 5468
rect 22364 5466 22420 5468
rect 22444 5466 22500 5468
rect 22204 5414 22250 5466
rect 22250 5414 22260 5466
rect 22284 5414 22314 5466
rect 22314 5414 22326 5466
rect 22326 5414 22340 5466
rect 22364 5414 22378 5466
rect 22378 5414 22390 5466
rect 22390 5414 22420 5466
rect 22444 5414 22454 5466
rect 22454 5414 22500 5466
rect 22204 5412 22260 5414
rect 22284 5412 22340 5414
rect 22364 5412 22420 5414
rect 22444 5412 22500 5414
rect 22204 4378 22260 4380
rect 22284 4378 22340 4380
rect 22364 4378 22420 4380
rect 22444 4378 22500 4380
rect 22204 4326 22250 4378
rect 22250 4326 22260 4378
rect 22284 4326 22314 4378
rect 22314 4326 22326 4378
rect 22326 4326 22340 4378
rect 22364 4326 22378 4378
rect 22378 4326 22390 4378
rect 22390 4326 22420 4378
rect 22444 4326 22454 4378
rect 22454 4326 22500 4378
rect 22204 4324 22260 4326
rect 22284 4324 22340 4326
rect 22364 4324 22420 4326
rect 22444 4324 22500 4326
rect 25746 29946 25802 29948
rect 25826 29946 25882 29948
rect 25906 29946 25962 29948
rect 25986 29946 26042 29948
rect 25746 29894 25792 29946
rect 25792 29894 25802 29946
rect 25826 29894 25856 29946
rect 25856 29894 25868 29946
rect 25868 29894 25882 29946
rect 25906 29894 25920 29946
rect 25920 29894 25932 29946
rect 25932 29894 25962 29946
rect 25986 29894 25996 29946
rect 25996 29894 26042 29946
rect 25746 29892 25802 29894
rect 25826 29892 25882 29894
rect 25906 29892 25962 29894
rect 25986 29892 26042 29894
rect 29287 30490 29343 30492
rect 29367 30490 29423 30492
rect 29447 30490 29503 30492
rect 29527 30490 29583 30492
rect 29287 30438 29333 30490
rect 29333 30438 29343 30490
rect 29367 30438 29397 30490
rect 29397 30438 29409 30490
rect 29409 30438 29423 30490
rect 29447 30438 29461 30490
rect 29461 30438 29473 30490
rect 29473 30438 29503 30490
rect 29527 30438 29537 30490
rect 29537 30438 29583 30490
rect 29287 30436 29343 30438
rect 29367 30436 29423 30438
rect 29447 30436 29503 30438
rect 29527 30436 29583 30438
rect 29287 29402 29343 29404
rect 29367 29402 29423 29404
rect 29447 29402 29503 29404
rect 29527 29402 29583 29404
rect 29287 29350 29333 29402
rect 29333 29350 29343 29402
rect 29367 29350 29397 29402
rect 29397 29350 29409 29402
rect 29409 29350 29423 29402
rect 29447 29350 29461 29402
rect 29461 29350 29473 29402
rect 29473 29350 29503 29402
rect 29527 29350 29537 29402
rect 29537 29350 29583 29402
rect 29287 29348 29343 29350
rect 29367 29348 29423 29350
rect 29447 29348 29503 29350
rect 29527 29348 29583 29350
rect 28722 29008 28778 29064
rect 25746 28858 25802 28860
rect 25826 28858 25882 28860
rect 25906 28858 25962 28860
rect 25986 28858 26042 28860
rect 25746 28806 25792 28858
rect 25792 28806 25802 28858
rect 25826 28806 25856 28858
rect 25856 28806 25868 28858
rect 25868 28806 25882 28858
rect 25906 28806 25920 28858
rect 25920 28806 25932 28858
rect 25932 28806 25962 28858
rect 25986 28806 25996 28858
rect 25996 28806 26042 28858
rect 25746 28804 25802 28806
rect 25826 28804 25882 28806
rect 25906 28804 25962 28806
rect 25986 28804 26042 28806
rect 29287 28314 29343 28316
rect 29367 28314 29423 28316
rect 29447 28314 29503 28316
rect 29527 28314 29583 28316
rect 29287 28262 29333 28314
rect 29333 28262 29343 28314
rect 29367 28262 29397 28314
rect 29397 28262 29409 28314
rect 29409 28262 29423 28314
rect 29447 28262 29461 28314
rect 29461 28262 29473 28314
rect 29473 28262 29503 28314
rect 29527 28262 29537 28314
rect 29537 28262 29583 28314
rect 29287 28260 29343 28262
rect 29367 28260 29423 28262
rect 29447 28260 29503 28262
rect 29527 28260 29583 28262
rect 25746 27770 25802 27772
rect 25826 27770 25882 27772
rect 25906 27770 25962 27772
rect 25986 27770 26042 27772
rect 25746 27718 25792 27770
rect 25792 27718 25802 27770
rect 25826 27718 25856 27770
rect 25856 27718 25868 27770
rect 25868 27718 25882 27770
rect 25906 27718 25920 27770
rect 25920 27718 25932 27770
rect 25932 27718 25962 27770
rect 25986 27718 25996 27770
rect 25996 27718 26042 27770
rect 25746 27716 25802 27718
rect 25826 27716 25882 27718
rect 25906 27716 25962 27718
rect 25986 27716 26042 27718
rect 29287 27226 29343 27228
rect 29367 27226 29423 27228
rect 29447 27226 29503 27228
rect 29527 27226 29583 27228
rect 29287 27174 29333 27226
rect 29333 27174 29343 27226
rect 29367 27174 29397 27226
rect 29397 27174 29409 27226
rect 29409 27174 29423 27226
rect 29447 27174 29461 27226
rect 29461 27174 29473 27226
rect 29473 27174 29503 27226
rect 29527 27174 29537 27226
rect 29537 27174 29583 27226
rect 29287 27172 29343 27174
rect 29367 27172 29423 27174
rect 29447 27172 29503 27174
rect 29527 27172 29583 27174
rect 25746 26682 25802 26684
rect 25826 26682 25882 26684
rect 25906 26682 25962 26684
rect 25986 26682 26042 26684
rect 25746 26630 25792 26682
rect 25792 26630 25802 26682
rect 25826 26630 25856 26682
rect 25856 26630 25868 26682
rect 25868 26630 25882 26682
rect 25906 26630 25920 26682
rect 25920 26630 25932 26682
rect 25932 26630 25962 26682
rect 25986 26630 25996 26682
rect 25996 26630 26042 26682
rect 25746 26628 25802 26630
rect 25826 26628 25882 26630
rect 25906 26628 25962 26630
rect 25986 26628 26042 26630
rect 25746 25594 25802 25596
rect 25826 25594 25882 25596
rect 25906 25594 25962 25596
rect 25986 25594 26042 25596
rect 25746 25542 25792 25594
rect 25792 25542 25802 25594
rect 25826 25542 25856 25594
rect 25856 25542 25868 25594
rect 25868 25542 25882 25594
rect 25906 25542 25920 25594
rect 25920 25542 25932 25594
rect 25932 25542 25962 25594
rect 25986 25542 25996 25594
rect 25996 25542 26042 25594
rect 25746 25540 25802 25542
rect 25826 25540 25882 25542
rect 25906 25540 25962 25542
rect 25986 25540 26042 25542
rect 25746 24506 25802 24508
rect 25826 24506 25882 24508
rect 25906 24506 25962 24508
rect 25986 24506 26042 24508
rect 25746 24454 25792 24506
rect 25792 24454 25802 24506
rect 25826 24454 25856 24506
rect 25856 24454 25868 24506
rect 25868 24454 25882 24506
rect 25906 24454 25920 24506
rect 25920 24454 25932 24506
rect 25932 24454 25962 24506
rect 25986 24454 25996 24506
rect 25996 24454 26042 24506
rect 25746 24452 25802 24454
rect 25826 24452 25882 24454
rect 25906 24452 25962 24454
rect 25986 24452 26042 24454
rect 25746 23418 25802 23420
rect 25826 23418 25882 23420
rect 25906 23418 25962 23420
rect 25986 23418 26042 23420
rect 25746 23366 25792 23418
rect 25792 23366 25802 23418
rect 25826 23366 25856 23418
rect 25856 23366 25868 23418
rect 25868 23366 25882 23418
rect 25906 23366 25920 23418
rect 25920 23366 25932 23418
rect 25932 23366 25962 23418
rect 25986 23366 25996 23418
rect 25996 23366 26042 23418
rect 25746 23364 25802 23366
rect 25826 23364 25882 23366
rect 25906 23364 25962 23366
rect 25986 23364 26042 23366
rect 24674 22072 24730 22128
rect 25746 22330 25802 22332
rect 25826 22330 25882 22332
rect 25906 22330 25962 22332
rect 25986 22330 26042 22332
rect 25746 22278 25792 22330
rect 25792 22278 25802 22330
rect 25826 22278 25856 22330
rect 25856 22278 25868 22330
rect 25868 22278 25882 22330
rect 25906 22278 25920 22330
rect 25920 22278 25932 22330
rect 25932 22278 25962 22330
rect 25986 22278 25996 22330
rect 25996 22278 26042 22330
rect 25746 22276 25802 22278
rect 25826 22276 25882 22278
rect 25906 22276 25962 22278
rect 25986 22276 26042 22278
rect 25318 21548 25374 21584
rect 26146 21936 26202 21992
rect 25318 21528 25320 21548
rect 25320 21528 25372 21548
rect 25372 21528 25374 21548
rect 25746 21242 25802 21244
rect 25826 21242 25882 21244
rect 25906 21242 25962 21244
rect 25986 21242 26042 21244
rect 25746 21190 25792 21242
rect 25792 21190 25802 21242
rect 25826 21190 25856 21242
rect 25856 21190 25868 21242
rect 25868 21190 25882 21242
rect 25906 21190 25920 21242
rect 25920 21190 25932 21242
rect 25932 21190 25962 21242
rect 25986 21190 25996 21242
rect 25996 21190 26042 21242
rect 25746 21188 25802 21190
rect 25826 21188 25882 21190
rect 25906 21188 25962 21190
rect 25986 21188 26042 21190
rect 25594 21120 25650 21176
rect 27066 21412 27122 21448
rect 27066 21392 27068 21412
rect 27068 21392 27120 21412
rect 27120 21392 27122 21412
rect 25746 20154 25802 20156
rect 25826 20154 25882 20156
rect 25906 20154 25962 20156
rect 25986 20154 26042 20156
rect 25746 20102 25792 20154
rect 25792 20102 25802 20154
rect 25826 20102 25856 20154
rect 25856 20102 25868 20154
rect 25868 20102 25882 20154
rect 25906 20102 25920 20154
rect 25920 20102 25932 20154
rect 25932 20102 25962 20154
rect 25986 20102 25996 20154
rect 25996 20102 26042 20154
rect 25746 20100 25802 20102
rect 25826 20100 25882 20102
rect 25906 20100 25962 20102
rect 25986 20100 26042 20102
rect 25746 19066 25802 19068
rect 25826 19066 25882 19068
rect 25906 19066 25962 19068
rect 25986 19066 26042 19068
rect 25746 19014 25792 19066
rect 25792 19014 25802 19066
rect 25826 19014 25856 19066
rect 25856 19014 25868 19066
rect 25868 19014 25882 19066
rect 25906 19014 25920 19066
rect 25920 19014 25932 19066
rect 25932 19014 25962 19066
rect 25986 19014 25996 19066
rect 25996 19014 26042 19066
rect 25746 19012 25802 19014
rect 25826 19012 25882 19014
rect 25906 19012 25962 19014
rect 25986 19012 26042 19014
rect 25746 17978 25802 17980
rect 25826 17978 25882 17980
rect 25906 17978 25962 17980
rect 25986 17978 26042 17980
rect 25746 17926 25792 17978
rect 25792 17926 25802 17978
rect 25826 17926 25856 17978
rect 25856 17926 25868 17978
rect 25868 17926 25882 17978
rect 25906 17926 25920 17978
rect 25920 17926 25932 17978
rect 25932 17926 25962 17978
rect 25986 17926 25996 17978
rect 25996 17926 26042 17978
rect 25746 17924 25802 17926
rect 25826 17924 25882 17926
rect 25906 17924 25962 17926
rect 25986 17924 26042 17926
rect 26146 17720 26202 17776
rect 26054 17196 26110 17232
rect 26054 17176 26056 17196
rect 26056 17176 26108 17196
rect 26108 17176 26110 17196
rect 25746 16890 25802 16892
rect 25826 16890 25882 16892
rect 25906 16890 25962 16892
rect 25986 16890 26042 16892
rect 25746 16838 25792 16890
rect 25792 16838 25802 16890
rect 25826 16838 25856 16890
rect 25856 16838 25868 16890
rect 25868 16838 25882 16890
rect 25906 16838 25920 16890
rect 25920 16838 25932 16890
rect 25932 16838 25962 16890
rect 25986 16838 25996 16890
rect 25996 16838 26042 16890
rect 25746 16836 25802 16838
rect 25826 16836 25882 16838
rect 25906 16836 25962 16838
rect 25986 16836 26042 16838
rect 26054 16396 26056 16416
rect 26056 16396 26108 16416
rect 26108 16396 26110 16416
rect 26054 16360 26110 16396
rect 25134 15408 25190 15464
rect 25746 15802 25802 15804
rect 25826 15802 25882 15804
rect 25906 15802 25962 15804
rect 25986 15802 26042 15804
rect 25746 15750 25792 15802
rect 25792 15750 25802 15802
rect 25826 15750 25856 15802
rect 25856 15750 25868 15802
rect 25868 15750 25882 15802
rect 25906 15750 25920 15802
rect 25920 15750 25932 15802
rect 25932 15750 25962 15802
rect 25986 15750 25996 15802
rect 25996 15750 26042 15802
rect 25746 15748 25802 15750
rect 25826 15748 25882 15750
rect 25906 15748 25962 15750
rect 25986 15748 26042 15750
rect 26698 17584 26754 17640
rect 26514 15408 26570 15464
rect 25746 14714 25802 14716
rect 25826 14714 25882 14716
rect 25906 14714 25962 14716
rect 25986 14714 26042 14716
rect 25746 14662 25792 14714
rect 25792 14662 25802 14714
rect 25826 14662 25856 14714
rect 25856 14662 25868 14714
rect 25868 14662 25882 14714
rect 25906 14662 25920 14714
rect 25920 14662 25932 14714
rect 25932 14662 25962 14714
rect 25986 14662 25996 14714
rect 25996 14662 26042 14714
rect 25746 14660 25802 14662
rect 25826 14660 25882 14662
rect 25906 14660 25962 14662
rect 25986 14660 26042 14662
rect 27526 17604 27582 17640
rect 27526 17584 27528 17604
rect 27528 17584 27580 17604
rect 27580 17584 27582 17604
rect 27250 17196 27306 17232
rect 27250 17176 27252 17196
rect 27252 17176 27304 17196
rect 27304 17176 27306 17196
rect 27710 17176 27766 17232
rect 27986 16396 27988 16416
rect 27988 16396 28040 16416
rect 28040 16396 28042 16416
rect 27986 16360 28042 16396
rect 25746 13626 25802 13628
rect 25826 13626 25882 13628
rect 25906 13626 25962 13628
rect 25986 13626 26042 13628
rect 25746 13574 25792 13626
rect 25792 13574 25802 13626
rect 25826 13574 25856 13626
rect 25856 13574 25868 13626
rect 25868 13574 25882 13626
rect 25906 13574 25920 13626
rect 25920 13574 25932 13626
rect 25932 13574 25962 13626
rect 25986 13574 25996 13626
rect 25996 13574 26042 13626
rect 25746 13572 25802 13574
rect 25826 13572 25882 13574
rect 25906 13572 25962 13574
rect 25986 13572 26042 13574
rect 25746 12538 25802 12540
rect 25826 12538 25882 12540
rect 25906 12538 25962 12540
rect 25986 12538 26042 12540
rect 25746 12486 25792 12538
rect 25792 12486 25802 12538
rect 25826 12486 25856 12538
rect 25856 12486 25868 12538
rect 25868 12486 25882 12538
rect 25906 12486 25920 12538
rect 25920 12486 25932 12538
rect 25932 12486 25962 12538
rect 25986 12486 25996 12538
rect 25996 12486 26042 12538
rect 25746 12484 25802 12486
rect 25826 12484 25882 12486
rect 25906 12484 25962 12486
rect 25986 12484 26042 12486
rect 24398 11056 24454 11112
rect 24306 5480 24362 5536
rect 25746 11450 25802 11452
rect 25826 11450 25882 11452
rect 25906 11450 25962 11452
rect 25986 11450 26042 11452
rect 25746 11398 25792 11450
rect 25792 11398 25802 11450
rect 25826 11398 25856 11450
rect 25856 11398 25868 11450
rect 25868 11398 25882 11450
rect 25906 11398 25920 11450
rect 25920 11398 25932 11450
rect 25932 11398 25962 11450
rect 25986 11398 25996 11450
rect 25996 11398 26042 11450
rect 25746 11396 25802 11398
rect 25826 11396 25882 11398
rect 25906 11396 25962 11398
rect 25986 11396 26042 11398
rect 25746 10362 25802 10364
rect 25826 10362 25882 10364
rect 25906 10362 25962 10364
rect 25986 10362 26042 10364
rect 25746 10310 25792 10362
rect 25792 10310 25802 10362
rect 25826 10310 25856 10362
rect 25856 10310 25868 10362
rect 25868 10310 25882 10362
rect 25906 10310 25920 10362
rect 25920 10310 25932 10362
rect 25932 10310 25962 10362
rect 25986 10310 25996 10362
rect 25996 10310 26042 10362
rect 25746 10308 25802 10310
rect 25826 10308 25882 10310
rect 25906 10308 25962 10310
rect 25986 10308 26042 10310
rect 25746 9274 25802 9276
rect 25826 9274 25882 9276
rect 25906 9274 25962 9276
rect 25986 9274 26042 9276
rect 25746 9222 25792 9274
rect 25792 9222 25802 9274
rect 25826 9222 25856 9274
rect 25856 9222 25868 9274
rect 25868 9222 25882 9274
rect 25906 9222 25920 9274
rect 25920 9222 25932 9274
rect 25932 9222 25962 9274
rect 25986 9222 25996 9274
rect 25996 9222 26042 9274
rect 25746 9220 25802 9222
rect 25826 9220 25882 9222
rect 25906 9220 25962 9222
rect 25986 9220 26042 9222
rect 26146 8492 26202 8528
rect 26146 8472 26148 8492
rect 26148 8472 26200 8492
rect 26200 8472 26202 8492
rect 25746 8186 25802 8188
rect 25826 8186 25882 8188
rect 25906 8186 25962 8188
rect 25986 8186 26042 8188
rect 25746 8134 25792 8186
rect 25792 8134 25802 8186
rect 25826 8134 25856 8186
rect 25856 8134 25868 8186
rect 25868 8134 25882 8186
rect 25906 8134 25920 8186
rect 25920 8134 25932 8186
rect 25932 8134 25962 8186
rect 25986 8134 25996 8186
rect 25996 8134 26042 8186
rect 25746 8132 25802 8134
rect 25826 8132 25882 8134
rect 25906 8132 25962 8134
rect 25986 8132 26042 8134
rect 25746 7098 25802 7100
rect 25826 7098 25882 7100
rect 25906 7098 25962 7100
rect 25986 7098 26042 7100
rect 25746 7046 25792 7098
rect 25792 7046 25802 7098
rect 25826 7046 25856 7098
rect 25856 7046 25868 7098
rect 25868 7046 25882 7098
rect 25906 7046 25920 7098
rect 25920 7046 25932 7098
rect 25932 7046 25962 7098
rect 25986 7046 25996 7098
rect 25996 7046 26042 7098
rect 25746 7044 25802 7046
rect 25826 7044 25882 7046
rect 25906 7044 25962 7046
rect 25986 7044 26042 7046
rect 25746 6010 25802 6012
rect 25826 6010 25882 6012
rect 25906 6010 25962 6012
rect 25986 6010 26042 6012
rect 25746 5958 25792 6010
rect 25792 5958 25802 6010
rect 25826 5958 25856 6010
rect 25856 5958 25868 6010
rect 25868 5958 25882 6010
rect 25906 5958 25920 6010
rect 25920 5958 25932 6010
rect 25932 5958 25962 6010
rect 25986 5958 25996 6010
rect 25996 5958 26042 6010
rect 25746 5956 25802 5958
rect 25826 5956 25882 5958
rect 25906 5956 25962 5958
rect 25986 5956 26042 5958
rect 25746 4922 25802 4924
rect 25826 4922 25882 4924
rect 25906 4922 25962 4924
rect 25986 4922 26042 4924
rect 25746 4870 25792 4922
rect 25792 4870 25802 4922
rect 25826 4870 25856 4922
rect 25856 4870 25868 4922
rect 25868 4870 25882 4922
rect 25906 4870 25920 4922
rect 25920 4870 25932 4922
rect 25932 4870 25962 4922
rect 25986 4870 25996 4922
rect 25996 4870 26042 4922
rect 25746 4868 25802 4870
rect 25826 4868 25882 4870
rect 25906 4868 25962 4870
rect 25986 4868 26042 4870
rect 24214 3984 24270 4040
rect 25746 3834 25802 3836
rect 25826 3834 25882 3836
rect 25906 3834 25962 3836
rect 25986 3834 26042 3836
rect 25746 3782 25792 3834
rect 25792 3782 25802 3834
rect 25826 3782 25856 3834
rect 25856 3782 25868 3834
rect 25868 3782 25882 3834
rect 25906 3782 25920 3834
rect 25920 3782 25932 3834
rect 25932 3782 25962 3834
rect 25986 3782 25996 3834
rect 25996 3782 26042 3834
rect 25746 3780 25802 3782
rect 25826 3780 25882 3782
rect 25906 3780 25962 3782
rect 25986 3780 26042 3782
rect 22204 3290 22260 3292
rect 22284 3290 22340 3292
rect 22364 3290 22420 3292
rect 22444 3290 22500 3292
rect 22204 3238 22250 3290
rect 22250 3238 22260 3290
rect 22284 3238 22314 3290
rect 22314 3238 22326 3290
rect 22326 3238 22340 3290
rect 22364 3238 22378 3290
rect 22378 3238 22390 3290
rect 22390 3238 22420 3290
rect 22444 3238 22454 3290
rect 22454 3238 22500 3290
rect 22204 3236 22260 3238
rect 22284 3236 22340 3238
rect 22364 3236 22420 3238
rect 22444 3236 22500 3238
rect 27802 8472 27858 8528
rect 28998 26560 29054 26616
rect 29287 26138 29343 26140
rect 29367 26138 29423 26140
rect 29447 26138 29503 26140
rect 29527 26138 29583 26140
rect 29287 26086 29333 26138
rect 29333 26086 29343 26138
rect 29367 26086 29397 26138
rect 29397 26086 29409 26138
rect 29409 26086 29423 26138
rect 29447 26086 29461 26138
rect 29461 26086 29473 26138
rect 29473 26086 29503 26138
rect 29527 26086 29537 26138
rect 29537 26086 29583 26138
rect 29287 26084 29343 26086
rect 29367 26084 29423 26086
rect 29447 26084 29503 26086
rect 29527 26084 29583 26086
rect 29287 25050 29343 25052
rect 29367 25050 29423 25052
rect 29447 25050 29503 25052
rect 29527 25050 29583 25052
rect 29287 24998 29333 25050
rect 29333 24998 29343 25050
rect 29367 24998 29397 25050
rect 29397 24998 29409 25050
rect 29409 24998 29423 25050
rect 29447 24998 29461 25050
rect 29461 24998 29473 25050
rect 29473 24998 29503 25050
rect 29527 24998 29537 25050
rect 29537 24998 29583 25050
rect 29287 24996 29343 24998
rect 29367 24996 29423 24998
rect 29447 24996 29503 24998
rect 29527 24996 29583 24998
rect 29287 23962 29343 23964
rect 29367 23962 29423 23964
rect 29447 23962 29503 23964
rect 29527 23962 29583 23964
rect 29287 23910 29333 23962
rect 29333 23910 29343 23962
rect 29367 23910 29397 23962
rect 29397 23910 29409 23962
rect 29409 23910 29423 23962
rect 29447 23910 29461 23962
rect 29461 23910 29473 23962
rect 29473 23910 29503 23962
rect 29527 23910 29537 23962
rect 29537 23910 29583 23962
rect 29287 23908 29343 23910
rect 29367 23908 29423 23910
rect 29447 23908 29503 23910
rect 29527 23908 29583 23910
rect 29287 22874 29343 22876
rect 29367 22874 29423 22876
rect 29447 22874 29503 22876
rect 29527 22874 29583 22876
rect 29287 22822 29333 22874
rect 29333 22822 29343 22874
rect 29367 22822 29397 22874
rect 29397 22822 29409 22874
rect 29409 22822 29423 22874
rect 29447 22822 29461 22874
rect 29461 22822 29473 22874
rect 29473 22822 29503 22874
rect 29527 22822 29537 22874
rect 29537 22822 29583 22874
rect 29287 22820 29343 22822
rect 29367 22820 29423 22822
rect 29447 22820 29503 22822
rect 29527 22820 29583 22822
rect 28998 22500 29054 22536
rect 28998 22480 29000 22500
rect 29000 22480 29052 22500
rect 29052 22480 29054 22500
rect 29287 21786 29343 21788
rect 29367 21786 29423 21788
rect 29447 21786 29503 21788
rect 29527 21786 29583 21788
rect 29287 21734 29333 21786
rect 29333 21734 29343 21786
rect 29367 21734 29397 21786
rect 29397 21734 29409 21786
rect 29409 21734 29423 21786
rect 29447 21734 29461 21786
rect 29461 21734 29473 21786
rect 29473 21734 29503 21786
rect 29527 21734 29537 21786
rect 29537 21734 29583 21786
rect 29287 21732 29343 21734
rect 29367 21732 29423 21734
rect 29447 21732 29503 21734
rect 29527 21732 29583 21734
rect 29287 20698 29343 20700
rect 29367 20698 29423 20700
rect 29447 20698 29503 20700
rect 29527 20698 29583 20700
rect 29287 20646 29333 20698
rect 29333 20646 29343 20698
rect 29367 20646 29397 20698
rect 29397 20646 29409 20698
rect 29409 20646 29423 20698
rect 29447 20646 29461 20698
rect 29461 20646 29473 20698
rect 29473 20646 29503 20698
rect 29527 20646 29537 20698
rect 29537 20646 29583 20698
rect 29287 20644 29343 20646
rect 29367 20644 29423 20646
rect 29447 20644 29503 20646
rect 29527 20644 29583 20646
rect 25746 2746 25802 2748
rect 25826 2746 25882 2748
rect 25906 2746 25962 2748
rect 25986 2746 26042 2748
rect 25746 2694 25792 2746
rect 25792 2694 25802 2746
rect 25826 2694 25856 2746
rect 25856 2694 25868 2746
rect 25868 2694 25882 2746
rect 25906 2694 25920 2746
rect 25920 2694 25932 2746
rect 25932 2694 25962 2746
rect 25986 2694 25996 2746
rect 25996 2694 26042 2746
rect 25746 2692 25802 2694
rect 25826 2692 25882 2694
rect 25906 2692 25962 2694
rect 25986 2692 26042 2694
rect 29287 19610 29343 19612
rect 29367 19610 29423 19612
rect 29447 19610 29503 19612
rect 29527 19610 29583 19612
rect 29287 19558 29333 19610
rect 29333 19558 29343 19610
rect 29367 19558 29397 19610
rect 29397 19558 29409 19610
rect 29409 19558 29423 19610
rect 29447 19558 29461 19610
rect 29461 19558 29473 19610
rect 29473 19558 29503 19610
rect 29527 19558 29537 19610
rect 29537 19558 29583 19610
rect 29287 19556 29343 19558
rect 29367 19556 29423 19558
rect 29447 19556 29503 19558
rect 29527 19556 29583 19558
rect 29458 18672 29514 18728
rect 29287 18522 29343 18524
rect 29367 18522 29423 18524
rect 29447 18522 29503 18524
rect 29527 18522 29583 18524
rect 29287 18470 29333 18522
rect 29333 18470 29343 18522
rect 29367 18470 29397 18522
rect 29397 18470 29409 18522
rect 29409 18470 29423 18522
rect 29447 18470 29461 18522
rect 29461 18470 29473 18522
rect 29473 18470 29503 18522
rect 29527 18470 29537 18522
rect 29537 18470 29583 18522
rect 29287 18468 29343 18470
rect 29367 18468 29423 18470
rect 29447 18468 29503 18470
rect 29527 18468 29583 18470
rect 29287 17434 29343 17436
rect 29367 17434 29423 17436
rect 29447 17434 29503 17436
rect 29527 17434 29583 17436
rect 29287 17382 29333 17434
rect 29333 17382 29343 17434
rect 29367 17382 29397 17434
rect 29397 17382 29409 17434
rect 29409 17382 29423 17434
rect 29447 17382 29461 17434
rect 29461 17382 29473 17434
rect 29473 17382 29503 17434
rect 29527 17382 29537 17434
rect 29537 17382 29583 17434
rect 29287 17380 29343 17382
rect 29367 17380 29423 17382
rect 29447 17380 29503 17382
rect 29527 17380 29583 17382
rect 29287 16346 29343 16348
rect 29367 16346 29423 16348
rect 29447 16346 29503 16348
rect 29527 16346 29583 16348
rect 29287 16294 29333 16346
rect 29333 16294 29343 16346
rect 29367 16294 29397 16346
rect 29397 16294 29409 16346
rect 29409 16294 29423 16346
rect 29447 16294 29461 16346
rect 29461 16294 29473 16346
rect 29473 16294 29503 16346
rect 29527 16294 29537 16346
rect 29537 16294 29583 16346
rect 29287 16292 29343 16294
rect 29367 16292 29423 16294
rect 29447 16292 29503 16294
rect 29527 16292 29583 16294
rect 29287 15258 29343 15260
rect 29367 15258 29423 15260
rect 29447 15258 29503 15260
rect 29527 15258 29583 15260
rect 29287 15206 29333 15258
rect 29333 15206 29343 15258
rect 29367 15206 29397 15258
rect 29397 15206 29409 15258
rect 29409 15206 29423 15258
rect 29447 15206 29461 15258
rect 29461 15206 29473 15258
rect 29473 15206 29503 15258
rect 29527 15206 29537 15258
rect 29537 15206 29583 15258
rect 29287 15204 29343 15206
rect 29367 15204 29423 15206
rect 29447 15204 29503 15206
rect 29527 15204 29583 15206
rect 28998 14320 29054 14376
rect 29287 14170 29343 14172
rect 29367 14170 29423 14172
rect 29447 14170 29503 14172
rect 29527 14170 29583 14172
rect 29287 14118 29333 14170
rect 29333 14118 29343 14170
rect 29367 14118 29397 14170
rect 29397 14118 29409 14170
rect 29409 14118 29423 14170
rect 29447 14118 29461 14170
rect 29461 14118 29473 14170
rect 29473 14118 29503 14170
rect 29527 14118 29537 14170
rect 29537 14118 29583 14170
rect 29287 14116 29343 14118
rect 29367 14116 29423 14118
rect 29447 14116 29503 14118
rect 29527 14116 29583 14118
rect 29287 13082 29343 13084
rect 29367 13082 29423 13084
rect 29447 13082 29503 13084
rect 29527 13082 29583 13084
rect 29287 13030 29333 13082
rect 29333 13030 29343 13082
rect 29367 13030 29397 13082
rect 29397 13030 29409 13082
rect 29409 13030 29423 13082
rect 29447 13030 29461 13082
rect 29461 13030 29473 13082
rect 29473 13030 29503 13082
rect 29527 13030 29537 13082
rect 29537 13030 29583 13082
rect 29287 13028 29343 13030
rect 29367 13028 29423 13030
rect 29447 13028 29503 13030
rect 29527 13028 29583 13030
rect 29287 11994 29343 11996
rect 29367 11994 29423 11996
rect 29447 11994 29503 11996
rect 29527 11994 29583 11996
rect 29287 11942 29333 11994
rect 29333 11942 29343 11994
rect 29367 11942 29397 11994
rect 29397 11942 29409 11994
rect 29409 11942 29423 11994
rect 29447 11942 29461 11994
rect 29461 11942 29473 11994
rect 29473 11942 29503 11994
rect 29527 11942 29537 11994
rect 29537 11942 29583 11994
rect 29287 11940 29343 11942
rect 29367 11940 29423 11942
rect 29447 11940 29503 11942
rect 29527 11940 29583 11942
rect 29090 11076 29146 11112
rect 29090 11056 29092 11076
rect 29092 11056 29144 11076
rect 29144 11056 29146 11076
rect 29287 10906 29343 10908
rect 29367 10906 29423 10908
rect 29447 10906 29503 10908
rect 29527 10906 29583 10908
rect 29287 10854 29333 10906
rect 29333 10854 29343 10906
rect 29367 10854 29397 10906
rect 29397 10854 29409 10906
rect 29409 10854 29423 10906
rect 29447 10854 29461 10906
rect 29461 10854 29473 10906
rect 29473 10854 29503 10906
rect 29527 10854 29537 10906
rect 29537 10854 29583 10906
rect 29287 10852 29343 10854
rect 29367 10852 29423 10854
rect 29447 10852 29503 10854
rect 29527 10852 29583 10854
rect 29287 9818 29343 9820
rect 29367 9818 29423 9820
rect 29447 9818 29503 9820
rect 29527 9818 29583 9820
rect 29287 9766 29333 9818
rect 29333 9766 29343 9818
rect 29367 9766 29397 9818
rect 29397 9766 29409 9818
rect 29409 9766 29423 9818
rect 29447 9766 29461 9818
rect 29461 9766 29473 9818
rect 29473 9766 29503 9818
rect 29527 9766 29537 9818
rect 29537 9766 29583 9818
rect 29287 9764 29343 9766
rect 29367 9764 29423 9766
rect 29447 9764 29503 9766
rect 29527 9764 29583 9766
rect 29287 8730 29343 8732
rect 29367 8730 29423 8732
rect 29447 8730 29503 8732
rect 29527 8730 29583 8732
rect 29287 8678 29333 8730
rect 29333 8678 29343 8730
rect 29367 8678 29397 8730
rect 29397 8678 29409 8730
rect 29409 8678 29423 8730
rect 29447 8678 29461 8730
rect 29461 8678 29473 8730
rect 29473 8678 29503 8730
rect 29527 8678 29537 8730
rect 29537 8678 29583 8730
rect 29287 8676 29343 8678
rect 29367 8676 29423 8678
rect 29447 8676 29503 8678
rect 29527 8676 29583 8678
rect 29287 7642 29343 7644
rect 29367 7642 29423 7644
rect 29447 7642 29503 7644
rect 29527 7642 29583 7644
rect 29287 7590 29333 7642
rect 29333 7590 29343 7642
rect 29367 7590 29397 7642
rect 29397 7590 29409 7642
rect 29409 7590 29423 7642
rect 29447 7590 29461 7642
rect 29461 7590 29473 7642
rect 29473 7590 29503 7642
rect 29527 7590 29537 7642
rect 29537 7590 29583 7642
rect 29287 7588 29343 7590
rect 29367 7588 29423 7590
rect 29447 7588 29503 7590
rect 29527 7588 29583 7590
rect 29090 6840 29146 6896
rect 29287 6554 29343 6556
rect 29367 6554 29423 6556
rect 29447 6554 29503 6556
rect 29527 6554 29583 6556
rect 29287 6502 29333 6554
rect 29333 6502 29343 6554
rect 29367 6502 29397 6554
rect 29397 6502 29409 6554
rect 29409 6502 29423 6554
rect 29447 6502 29461 6554
rect 29461 6502 29473 6554
rect 29473 6502 29503 6554
rect 29527 6502 29537 6554
rect 29537 6502 29583 6554
rect 29287 6500 29343 6502
rect 29367 6500 29423 6502
rect 29447 6500 29503 6502
rect 29527 6500 29583 6502
rect 29287 5466 29343 5468
rect 29367 5466 29423 5468
rect 29447 5466 29503 5468
rect 29527 5466 29583 5468
rect 29287 5414 29333 5466
rect 29333 5414 29343 5466
rect 29367 5414 29397 5466
rect 29397 5414 29409 5466
rect 29409 5414 29423 5466
rect 29447 5414 29461 5466
rect 29461 5414 29473 5466
rect 29473 5414 29503 5466
rect 29527 5414 29537 5466
rect 29537 5414 29583 5466
rect 29287 5412 29343 5414
rect 29367 5412 29423 5414
rect 29447 5412 29503 5414
rect 29527 5412 29583 5414
rect 29287 4378 29343 4380
rect 29367 4378 29423 4380
rect 29447 4378 29503 4380
rect 29527 4378 29583 4380
rect 29287 4326 29333 4378
rect 29333 4326 29343 4378
rect 29367 4326 29397 4378
rect 29397 4326 29409 4378
rect 29409 4326 29423 4378
rect 29447 4326 29461 4378
rect 29461 4326 29473 4378
rect 29473 4326 29503 4378
rect 29527 4326 29537 4378
rect 29537 4326 29583 4378
rect 29287 4324 29343 4326
rect 29367 4324 29423 4326
rect 29447 4324 29503 4326
rect 29527 4324 29583 4326
rect 29287 3290 29343 3292
rect 29367 3290 29423 3292
rect 29447 3290 29503 3292
rect 29527 3290 29583 3292
rect 29287 3238 29333 3290
rect 29333 3238 29343 3290
rect 29367 3238 29397 3290
rect 29397 3238 29409 3290
rect 29409 3238 29423 3290
rect 29447 3238 29461 3290
rect 29461 3238 29473 3290
rect 29473 3238 29503 3290
rect 29527 3238 29537 3290
rect 29537 3238 29583 3290
rect 29287 3236 29343 3238
rect 29367 3236 29423 3238
rect 29447 3236 29503 3238
rect 29527 3236 29583 3238
rect 28998 2796 29000 2816
rect 29000 2796 29052 2816
rect 29052 2796 29054 2816
rect 28998 2760 29054 2796
rect 8038 2202 8094 2204
rect 8118 2202 8174 2204
rect 8198 2202 8254 2204
rect 8278 2202 8334 2204
rect 8038 2150 8084 2202
rect 8084 2150 8094 2202
rect 8118 2150 8148 2202
rect 8148 2150 8160 2202
rect 8160 2150 8174 2202
rect 8198 2150 8212 2202
rect 8212 2150 8224 2202
rect 8224 2150 8254 2202
rect 8278 2150 8288 2202
rect 8288 2150 8334 2202
rect 8038 2148 8094 2150
rect 8118 2148 8174 2150
rect 8198 2148 8254 2150
rect 8278 2148 8334 2150
rect 15121 2202 15177 2204
rect 15201 2202 15257 2204
rect 15281 2202 15337 2204
rect 15361 2202 15417 2204
rect 15121 2150 15167 2202
rect 15167 2150 15177 2202
rect 15201 2150 15231 2202
rect 15231 2150 15243 2202
rect 15243 2150 15257 2202
rect 15281 2150 15295 2202
rect 15295 2150 15307 2202
rect 15307 2150 15337 2202
rect 15361 2150 15371 2202
rect 15371 2150 15417 2202
rect 15121 2148 15177 2150
rect 15201 2148 15257 2150
rect 15281 2148 15337 2150
rect 15361 2148 15417 2150
rect 22204 2202 22260 2204
rect 22284 2202 22340 2204
rect 22364 2202 22420 2204
rect 22444 2202 22500 2204
rect 22204 2150 22250 2202
rect 22250 2150 22260 2202
rect 22284 2150 22314 2202
rect 22314 2150 22326 2202
rect 22326 2150 22340 2202
rect 22364 2150 22378 2202
rect 22378 2150 22390 2202
rect 22390 2150 22420 2202
rect 22444 2150 22454 2202
rect 22454 2150 22500 2202
rect 22204 2148 22260 2150
rect 22284 2148 22340 2150
rect 22364 2148 22420 2150
rect 22444 2148 22500 2150
rect 29287 2202 29343 2204
rect 29367 2202 29423 2204
rect 29447 2202 29503 2204
rect 29527 2202 29583 2204
rect 29287 2150 29333 2202
rect 29333 2150 29343 2202
rect 29367 2150 29397 2202
rect 29397 2150 29409 2202
rect 29409 2150 29423 2202
rect 29447 2150 29461 2202
rect 29461 2150 29473 2202
rect 29473 2150 29503 2202
rect 29527 2150 29537 2202
rect 29537 2150 29583 2202
rect 29287 2148 29343 2150
rect 29367 2148 29423 2150
rect 29447 2148 29503 2150
rect 29527 2148 29583 2150
<< metal3 >>
rect 0 31378 800 31408
rect 0 31288 858 31378
rect 798 30970 858 31288
rect 1577 30970 1643 30973
rect 798 30968 1643 30970
rect 798 30912 1582 30968
rect 1638 30912 1643 30968
rect 798 30910 1643 30912
rect 1577 30907 1643 30910
rect 28901 30698 28967 30701
rect 29781 30698 30581 30728
rect 28901 30696 30581 30698
rect 28901 30640 28906 30696
rect 28962 30640 30581 30696
rect 28901 30638 30581 30640
rect 28901 30635 28967 30638
rect 29781 30608 30581 30638
rect 8028 30496 8344 30497
rect 8028 30432 8034 30496
rect 8098 30432 8114 30496
rect 8178 30432 8194 30496
rect 8258 30432 8274 30496
rect 8338 30432 8344 30496
rect 8028 30431 8344 30432
rect 15111 30496 15427 30497
rect 15111 30432 15117 30496
rect 15181 30432 15197 30496
rect 15261 30432 15277 30496
rect 15341 30432 15357 30496
rect 15421 30432 15427 30496
rect 15111 30431 15427 30432
rect 22194 30496 22510 30497
rect 22194 30432 22200 30496
rect 22264 30432 22280 30496
rect 22344 30432 22360 30496
rect 22424 30432 22440 30496
rect 22504 30432 22510 30496
rect 22194 30431 22510 30432
rect 29277 30496 29593 30497
rect 29277 30432 29283 30496
rect 29347 30432 29363 30496
rect 29427 30432 29443 30496
rect 29507 30432 29523 30496
rect 29587 30432 29593 30496
rect 29277 30431 29593 30432
rect 4487 29952 4803 29953
rect 4487 29888 4493 29952
rect 4557 29888 4573 29952
rect 4637 29888 4653 29952
rect 4717 29888 4733 29952
rect 4797 29888 4803 29952
rect 4487 29887 4803 29888
rect 11570 29952 11886 29953
rect 11570 29888 11576 29952
rect 11640 29888 11656 29952
rect 11720 29888 11736 29952
rect 11800 29888 11816 29952
rect 11880 29888 11886 29952
rect 11570 29887 11886 29888
rect 18653 29952 18969 29953
rect 18653 29888 18659 29952
rect 18723 29888 18739 29952
rect 18803 29888 18819 29952
rect 18883 29888 18899 29952
rect 18963 29888 18969 29952
rect 18653 29887 18969 29888
rect 25736 29952 26052 29953
rect 25736 29888 25742 29952
rect 25806 29888 25822 29952
rect 25886 29888 25902 29952
rect 25966 29888 25982 29952
rect 26046 29888 26052 29952
rect 25736 29887 26052 29888
rect 8028 29408 8344 29409
rect 8028 29344 8034 29408
rect 8098 29344 8114 29408
rect 8178 29344 8194 29408
rect 8258 29344 8274 29408
rect 8338 29344 8344 29408
rect 8028 29343 8344 29344
rect 15111 29408 15427 29409
rect 15111 29344 15117 29408
rect 15181 29344 15197 29408
rect 15261 29344 15277 29408
rect 15341 29344 15357 29408
rect 15421 29344 15427 29408
rect 15111 29343 15427 29344
rect 22194 29408 22510 29409
rect 22194 29344 22200 29408
rect 22264 29344 22280 29408
rect 22344 29344 22360 29408
rect 22424 29344 22440 29408
rect 22504 29344 22510 29408
rect 22194 29343 22510 29344
rect 29277 29408 29593 29409
rect 29277 29344 29283 29408
rect 29347 29344 29363 29408
rect 29427 29344 29443 29408
rect 29507 29344 29523 29408
rect 29587 29344 29593 29408
rect 29277 29343 29593 29344
rect 28717 29068 28783 29069
rect 28717 29064 28764 29068
rect 28828 29066 28834 29068
rect 28717 29008 28722 29064
rect 28717 29004 28764 29008
rect 28828 29006 28874 29066
rect 28828 29004 28834 29006
rect 28717 29003 28783 29004
rect 4487 28864 4803 28865
rect 4487 28800 4493 28864
rect 4557 28800 4573 28864
rect 4637 28800 4653 28864
rect 4717 28800 4733 28864
rect 4797 28800 4803 28864
rect 4487 28799 4803 28800
rect 11570 28864 11886 28865
rect 11570 28800 11576 28864
rect 11640 28800 11656 28864
rect 11720 28800 11736 28864
rect 11800 28800 11816 28864
rect 11880 28800 11886 28864
rect 11570 28799 11886 28800
rect 18653 28864 18969 28865
rect 18653 28800 18659 28864
rect 18723 28800 18739 28864
rect 18803 28800 18819 28864
rect 18883 28800 18899 28864
rect 18963 28800 18969 28864
rect 18653 28799 18969 28800
rect 25736 28864 26052 28865
rect 25736 28800 25742 28864
rect 25806 28800 25822 28864
rect 25886 28800 25902 28864
rect 25966 28800 25982 28864
rect 26046 28800 26052 28864
rect 25736 28799 26052 28800
rect 13629 28658 13695 28661
rect 22001 28658 22067 28661
rect 13629 28656 22067 28658
rect 13629 28600 13634 28656
rect 13690 28600 22006 28656
rect 22062 28600 22067 28656
rect 13629 28598 22067 28600
rect 13629 28595 13695 28598
rect 22001 28595 22067 28598
rect 13629 28522 13695 28525
rect 17953 28522 18019 28525
rect 13629 28520 18019 28522
rect 13629 28464 13634 28520
rect 13690 28464 17958 28520
rect 18014 28464 18019 28520
rect 13629 28462 18019 28464
rect 13629 28459 13695 28462
rect 17953 28459 18019 28462
rect 8028 28320 8344 28321
rect 8028 28256 8034 28320
rect 8098 28256 8114 28320
rect 8178 28256 8194 28320
rect 8258 28256 8274 28320
rect 8338 28256 8344 28320
rect 8028 28255 8344 28256
rect 15111 28320 15427 28321
rect 15111 28256 15117 28320
rect 15181 28256 15197 28320
rect 15261 28256 15277 28320
rect 15341 28256 15357 28320
rect 15421 28256 15427 28320
rect 15111 28255 15427 28256
rect 22194 28320 22510 28321
rect 22194 28256 22200 28320
rect 22264 28256 22280 28320
rect 22344 28256 22360 28320
rect 22424 28256 22440 28320
rect 22504 28256 22510 28320
rect 22194 28255 22510 28256
rect 29277 28320 29593 28321
rect 29277 28256 29283 28320
rect 29347 28256 29363 28320
rect 29427 28256 29443 28320
rect 29507 28256 29523 28320
rect 29587 28256 29593 28320
rect 29277 28255 29593 28256
rect 11053 28114 11119 28117
rect 12341 28114 12407 28117
rect 19333 28114 19399 28117
rect 11053 28112 19399 28114
rect 11053 28056 11058 28112
rect 11114 28056 12346 28112
rect 12402 28056 19338 28112
rect 19394 28056 19399 28112
rect 11053 28054 19399 28056
rect 11053 28051 11119 28054
rect 12341 28051 12407 28054
rect 19333 28051 19399 28054
rect 13353 27978 13419 27981
rect 21265 27978 21331 27981
rect 13353 27976 21331 27978
rect 13353 27920 13358 27976
rect 13414 27920 21270 27976
rect 21326 27920 21331 27976
rect 13353 27918 21331 27920
rect 13353 27915 13419 27918
rect 21265 27915 21331 27918
rect 4487 27776 4803 27777
rect 4487 27712 4493 27776
rect 4557 27712 4573 27776
rect 4637 27712 4653 27776
rect 4717 27712 4733 27776
rect 4797 27712 4803 27776
rect 4487 27711 4803 27712
rect 11570 27776 11886 27777
rect 11570 27712 11576 27776
rect 11640 27712 11656 27776
rect 11720 27712 11736 27776
rect 11800 27712 11816 27776
rect 11880 27712 11886 27776
rect 11570 27711 11886 27712
rect 18653 27776 18969 27777
rect 18653 27712 18659 27776
rect 18723 27712 18739 27776
rect 18803 27712 18819 27776
rect 18883 27712 18899 27776
rect 18963 27712 18969 27776
rect 18653 27711 18969 27712
rect 25736 27776 26052 27777
rect 25736 27712 25742 27776
rect 25806 27712 25822 27776
rect 25886 27712 25902 27776
rect 25966 27712 25982 27776
rect 26046 27712 26052 27776
rect 25736 27711 26052 27712
rect 0 27298 800 27328
rect 933 27298 999 27301
rect 0 27296 999 27298
rect 0 27240 938 27296
rect 994 27240 999 27296
rect 0 27238 999 27240
rect 0 27208 800 27238
rect 933 27235 999 27238
rect 8028 27232 8344 27233
rect 8028 27168 8034 27232
rect 8098 27168 8114 27232
rect 8178 27168 8194 27232
rect 8258 27168 8274 27232
rect 8338 27168 8344 27232
rect 8028 27167 8344 27168
rect 15111 27232 15427 27233
rect 15111 27168 15117 27232
rect 15181 27168 15197 27232
rect 15261 27168 15277 27232
rect 15341 27168 15357 27232
rect 15421 27168 15427 27232
rect 15111 27167 15427 27168
rect 22194 27232 22510 27233
rect 22194 27168 22200 27232
rect 22264 27168 22280 27232
rect 22344 27168 22360 27232
rect 22424 27168 22440 27232
rect 22504 27168 22510 27232
rect 22194 27167 22510 27168
rect 29277 27232 29593 27233
rect 29277 27168 29283 27232
rect 29347 27168 29363 27232
rect 29427 27168 29443 27232
rect 29507 27168 29523 27232
rect 29587 27168 29593 27232
rect 29277 27167 29593 27168
rect 4487 26688 4803 26689
rect 4487 26624 4493 26688
rect 4557 26624 4573 26688
rect 4637 26624 4653 26688
rect 4717 26624 4733 26688
rect 4797 26624 4803 26688
rect 4487 26623 4803 26624
rect 11570 26688 11886 26689
rect 11570 26624 11576 26688
rect 11640 26624 11656 26688
rect 11720 26624 11736 26688
rect 11800 26624 11816 26688
rect 11880 26624 11886 26688
rect 11570 26623 11886 26624
rect 18653 26688 18969 26689
rect 18653 26624 18659 26688
rect 18723 26624 18739 26688
rect 18803 26624 18819 26688
rect 18883 26624 18899 26688
rect 18963 26624 18969 26688
rect 18653 26623 18969 26624
rect 25736 26688 26052 26689
rect 25736 26624 25742 26688
rect 25806 26624 25822 26688
rect 25886 26624 25902 26688
rect 25966 26624 25982 26688
rect 26046 26624 26052 26688
rect 25736 26623 26052 26624
rect 28993 26618 29059 26621
rect 29781 26618 30581 26648
rect 28993 26616 30581 26618
rect 28993 26560 28998 26616
rect 29054 26560 30581 26616
rect 28993 26558 30581 26560
rect 28993 26555 29059 26558
rect 29781 26528 30581 26558
rect 8028 26144 8344 26145
rect 8028 26080 8034 26144
rect 8098 26080 8114 26144
rect 8178 26080 8194 26144
rect 8258 26080 8274 26144
rect 8338 26080 8344 26144
rect 8028 26079 8344 26080
rect 15111 26144 15427 26145
rect 15111 26080 15117 26144
rect 15181 26080 15197 26144
rect 15261 26080 15277 26144
rect 15341 26080 15357 26144
rect 15421 26080 15427 26144
rect 15111 26079 15427 26080
rect 22194 26144 22510 26145
rect 22194 26080 22200 26144
rect 22264 26080 22280 26144
rect 22344 26080 22360 26144
rect 22424 26080 22440 26144
rect 22504 26080 22510 26144
rect 22194 26079 22510 26080
rect 29277 26144 29593 26145
rect 29277 26080 29283 26144
rect 29347 26080 29363 26144
rect 29427 26080 29443 26144
rect 29507 26080 29523 26144
rect 29587 26080 29593 26144
rect 29277 26079 29593 26080
rect 4487 25600 4803 25601
rect 4487 25536 4493 25600
rect 4557 25536 4573 25600
rect 4637 25536 4653 25600
rect 4717 25536 4733 25600
rect 4797 25536 4803 25600
rect 4487 25535 4803 25536
rect 11570 25600 11886 25601
rect 11570 25536 11576 25600
rect 11640 25536 11656 25600
rect 11720 25536 11736 25600
rect 11800 25536 11816 25600
rect 11880 25536 11886 25600
rect 11570 25535 11886 25536
rect 18653 25600 18969 25601
rect 18653 25536 18659 25600
rect 18723 25536 18739 25600
rect 18803 25536 18819 25600
rect 18883 25536 18899 25600
rect 18963 25536 18969 25600
rect 18653 25535 18969 25536
rect 25736 25600 26052 25601
rect 25736 25536 25742 25600
rect 25806 25536 25822 25600
rect 25886 25536 25902 25600
rect 25966 25536 25982 25600
rect 26046 25536 26052 25600
rect 25736 25535 26052 25536
rect 8028 25056 8344 25057
rect 8028 24992 8034 25056
rect 8098 24992 8114 25056
rect 8178 24992 8194 25056
rect 8258 24992 8274 25056
rect 8338 24992 8344 25056
rect 8028 24991 8344 24992
rect 15111 25056 15427 25057
rect 15111 24992 15117 25056
rect 15181 24992 15197 25056
rect 15261 24992 15277 25056
rect 15341 24992 15357 25056
rect 15421 24992 15427 25056
rect 15111 24991 15427 24992
rect 22194 25056 22510 25057
rect 22194 24992 22200 25056
rect 22264 24992 22280 25056
rect 22344 24992 22360 25056
rect 22424 24992 22440 25056
rect 22504 24992 22510 25056
rect 22194 24991 22510 24992
rect 29277 25056 29593 25057
rect 29277 24992 29283 25056
rect 29347 24992 29363 25056
rect 29427 24992 29443 25056
rect 29507 24992 29523 25056
rect 29587 24992 29593 25056
rect 29277 24991 29593 24992
rect 4487 24512 4803 24513
rect 4487 24448 4493 24512
rect 4557 24448 4573 24512
rect 4637 24448 4653 24512
rect 4717 24448 4733 24512
rect 4797 24448 4803 24512
rect 4487 24447 4803 24448
rect 11570 24512 11886 24513
rect 11570 24448 11576 24512
rect 11640 24448 11656 24512
rect 11720 24448 11736 24512
rect 11800 24448 11816 24512
rect 11880 24448 11886 24512
rect 11570 24447 11886 24448
rect 18653 24512 18969 24513
rect 18653 24448 18659 24512
rect 18723 24448 18739 24512
rect 18803 24448 18819 24512
rect 18883 24448 18899 24512
rect 18963 24448 18969 24512
rect 18653 24447 18969 24448
rect 25736 24512 26052 24513
rect 25736 24448 25742 24512
rect 25806 24448 25822 24512
rect 25886 24448 25902 24512
rect 25966 24448 25982 24512
rect 26046 24448 26052 24512
rect 25736 24447 26052 24448
rect 8028 23968 8344 23969
rect 8028 23904 8034 23968
rect 8098 23904 8114 23968
rect 8178 23904 8194 23968
rect 8258 23904 8274 23968
rect 8338 23904 8344 23968
rect 8028 23903 8344 23904
rect 15111 23968 15427 23969
rect 15111 23904 15117 23968
rect 15181 23904 15197 23968
rect 15261 23904 15277 23968
rect 15341 23904 15357 23968
rect 15421 23904 15427 23968
rect 15111 23903 15427 23904
rect 22194 23968 22510 23969
rect 22194 23904 22200 23968
rect 22264 23904 22280 23968
rect 22344 23904 22360 23968
rect 22424 23904 22440 23968
rect 22504 23904 22510 23968
rect 22194 23903 22510 23904
rect 29277 23968 29593 23969
rect 29277 23904 29283 23968
rect 29347 23904 29363 23968
rect 29427 23904 29443 23968
rect 29507 23904 29523 23968
rect 29587 23904 29593 23968
rect 29277 23903 29593 23904
rect 1577 23490 1643 23493
rect 798 23488 1643 23490
rect 798 23432 1582 23488
rect 1638 23432 1643 23488
rect 798 23430 1643 23432
rect 798 23248 858 23430
rect 1577 23427 1643 23430
rect 4487 23424 4803 23425
rect 4487 23360 4493 23424
rect 4557 23360 4573 23424
rect 4637 23360 4653 23424
rect 4717 23360 4733 23424
rect 4797 23360 4803 23424
rect 4487 23359 4803 23360
rect 11570 23424 11886 23425
rect 11570 23360 11576 23424
rect 11640 23360 11656 23424
rect 11720 23360 11736 23424
rect 11800 23360 11816 23424
rect 11880 23360 11886 23424
rect 11570 23359 11886 23360
rect 18653 23424 18969 23425
rect 18653 23360 18659 23424
rect 18723 23360 18739 23424
rect 18803 23360 18819 23424
rect 18883 23360 18899 23424
rect 18963 23360 18969 23424
rect 18653 23359 18969 23360
rect 25736 23424 26052 23425
rect 25736 23360 25742 23424
rect 25806 23360 25822 23424
rect 25886 23360 25902 23424
rect 25966 23360 25982 23424
rect 26046 23360 26052 23424
rect 25736 23359 26052 23360
rect 0 23158 858 23248
rect 0 23128 800 23158
rect 1485 23082 1551 23085
rect 21173 23082 21239 23085
rect 1485 23080 21239 23082
rect 1485 23024 1490 23080
rect 1546 23024 21178 23080
rect 21234 23024 21239 23080
rect 1485 23022 21239 23024
rect 1485 23019 1551 23022
rect 21173 23019 21239 23022
rect 8028 22880 8344 22881
rect 8028 22816 8034 22880
rect 8098 22816 8114 22880
rect 8178 22816 8194 22880
rect 8258 22816 8274 22880
rect 8338 22816 8344 22880
rect 8028 22815 8344 22816
rect 15111 22880 15427 22881
rect 15111 22816 15117 22880
rect 15181 22816 15197 22880
rect 15261 22816 15277 22880
rect 15341 22816 15357 22880
rect 15421 22816 15427 22880
rect 15111 22815 15427 22816
rect 22194 22880 22510 22881
rect 22194 22816 22200 22880
rect 22264 22816 22280 22880
rect 22344 22816 22360 22880
rect 22424 22816 22440 22880
rect 22504 22816 22510 22880
rect 22194 22815 22510 22816
rect 29277 22880 29593 22881
rect 29277 22816 29283 22880
rect 29347 22816 29363 22880
rect 29427 22816 29443 22880
rect 29507 22816 29523 22880
rect 29587 22816 29593 22880
rect 29277 22815 29593 22816
rect 24393 22540 24459 22541
rect 24342 22476 24348 22540
rect 24412 22538 24459 22540
rect 28993 22538 29059 22541
rect 29781 22538 30581 22568
rect 24412 22536 24504 22538
rect 24454 22480 24504 22536
rect 24412 22478 24504 22480
rect 28993 22536 30581 22538
rect 28993 22480 28998 22536
rect 29054 22480 30581 22536
rect 28993 22478 30581 22480
rect 24412 22476 24459 22478
rect 24393 22475 24459 22476
rect 28993 22475 29059 22478
rect 29781 22448 30581 22478
rect 4487 22336 4803 22337
rect 4487 22272 4493 22336
rect 4557 22272 4573 22336
rect 4637 22272 4653 22336
rect 4717 22272 4733 22336
rect 4797 22272 4803 22336
rect 4487 22271 4803 22272
rect 11570 22336 11886 22337
rect 11570 22272 11576 22336
rect 11640 22272 11656 22336
rect 11720 22272 11736 22336
rect 11800 22272 11816 22336
rect 11880 22272 11886 22336
rect 11570 22271 11886 22272
rect 18653 22336 18969 22337
rect 18653 22272 18659 22336
rect 18723 22272 18739 22336
rect 18803 22272 18819 22336
rect 18883 22272 18899 22336
rect 18963 22272 18969 22336
rect 18653 22271 18969 22272
rect 25736 22336 26052 22337
rect 25736 22272 25742 22336
rect 25806 22272 25822 22336
rect 25886 22272 25902 22336
rect 25966 22272 25982 22336
rect 26046 22272 26052 22336
rect 25736 22271 26052 22272
rect 8109 22266 8175 22269
rect 10593 22266 10659 22269
rect 8109 22264 10659 22266
rect 8109 22208 8114 22264
rect 8170 22208 10598 22264
rect 10654 22208 10659 22264
rect 8109 22206 10659 22208
rect 8109 22203 8175 22206
rect 10593 22203 10659 22206
rect 20345 22130 20411 22133
rect 24669 22130 24735 22133
rect 20345 22128 24735 22130
rect 20345 22072 20350 22128
rect 20406 22072 24674 22128
rect 24730 22072 24735 22128
rect 20345 22070 24735 22072
rect 20345 22067 20411 22070
rect 24669 22067 24735 22070
rect 5441 21994 5507 21997
rect 7281 21994 7347 21997
rect 5441 21992 7347 21994
rect 5441 21936 5446 21992
rect 5502 21936 7286 21992
rect 7342 21936 7347 21992
rect 5441 21934 7347 21936
rect 5441 21931 5507 21934
rect 7281 21931 7347 21934
rect 17677 21994 17743 21997
rect 26141 21994 26207 21997
rect 17677 21992 26207 21994
rect 17677 21936 17682 21992
rect 17738 21936 26146 21992
rect 26202 21936 26207 21992
rect 17677 21934 26207 21936
rect 17677 21931 17743 21934
rect 26141 21931 26207 21934
rect 8028 21792 8344 21793
rect 8028 21728 8034 21792
rect 8098 21728 8114 21792
rect 8178 21728 8194 21792
rect 8258 21728 8274 21792
rect 8338 21728 8344 21792
rect 8028 21727 8344 21728
rect 15111 21792 15427 21793
rect 15111 21728 15117 21792
rect 15181 21728 15197 21792
rect 15261 21728 15277 21792
rect 15341 21728 15357 21792
rect 15421 21728 15427 21792
rect 15111 21727 15427 21728
rect 22194 21792 22510 21793
rect 22194 21728 22200 21792
rect 22264 21728 22280 21792
rect 22344 21728 22360 21792
rect 22424 21728 22440 21792
rect 22504 21728 22510 21792
rect 22194 21727 22510 21728
rect 29277 21792 29593 21793
rect 29277 21728 29283 21792
rect 29347 21728 29363 21792
rect 29427 21728 29443 21792
rect 29507 21728 29523 21792
rect 29587 21728 29593 21792
rect 29277 21727 29593 21728
rect 4153 21586 4219 21589
rect 6913 21586 6979 21589
rect 4153 21584 6979 21586
rect 4153 21528 4158 21584
rect 4214 21528 6918 21584
rect 6974 21528 6979 21584
rect 4153 21526 6979 21528
rect 4153 21523 4219 21526
rect 6913 21523 6979 21526
rect 21817 21586 21883 21589
rect 25313 21586 25379 21589
rect 21817 21584 25379 21586
rect 21817 21528 21822 21584
rect 21878 21528 25318 21584
rect 25374 21528 25379 21584
rect 21817 21526 25379 21528
rect 21817 21523 21883 21526
rect 25313 21523 25379 21526
rect 5809 21450 5875 21453
rect 8385 21450 8451 21453
rect 5809 21448 8451 21450
rect 5809 21392 5814 21448
rect 5870 21392 8390 21448
rect 8446 21392 8451 21448
rect 5809 21390 8451 21392
rect 5809 21387 5875 21390
rect 8385 21387 8451 21390
rect 9857 21450 9923 21453
rect 27061 21450 27127 21453
rect 9857 21448 27127 21450
rect 9857 21392 9862 21448
rect 9918 21392 27066 21448
rect 27122 21392 27127 21448
rect 9857 21390 27127 21392
rect 9857 21387 9923 21390
rect 27061 21387 27127 21390
rect 5901 21314 5967 21317
rect 8569 21314 8635 21317
rect 5901 21312 8635 21314
rect 5901 21256 5906 21312
rect 5962 21256 8574 21312
rect 8630 21256 8635 21312
rect 5901 21254 8635 21256
rect 5901 21251 5967 21254
rect 8569 21251 8635 21254
rect 4487 21248 4803 21249
rect 4487 21184 4493 21248
rect 4557 21184 4573 21248
rect 4637 21184 4653 21248
rect 4717 21184 4733 21248
rect 4797 21184 4803 21248
rect 4487 21183 4803 21184
rect 11570 21248 11886 21249
rect 11570 21184 11576 21248
rect 11640 21184 11656 21248
rect 11720 21184 11736 21248
rect 11800 21184 11816 21248
rect 11880 21184 11886 21248
rect 11570 21183 11886 21184
rect 18653 21248 18969 21249
rect 18653 21184 18659 21248
rect 18723 21184 18739 21248
rect 18803 21184 18819 21248
rect 18883 21184 18899 21248
rect 18963 21184 18969 21248
rect 18653 21183 18969 21184
rect 25736 21248 26052 21249
rect 25736 21184 25742 21248
rect 25806 21184 25822 21248
rect 25886 21184 25902 21248
rect 25966 21184 25982 21248
rect 26046 21184 26052 21248
rect 25736 21183 26052 21184
rect 22185 21178 22251 21181
rect 22921 21178 22987 21181
rect 22185 21176 22987 21178
rect 22185 21120 22190 21176
rect 22246 21120 22926 21176
rect 22982 21120 22987 21176
rect 22185 21118 22987 21120
rect 22185 21115 22251 21118
rect 22921 21115 22987 21118
rect 23473 21178 23539 21181
rect 25589 21178 25655 21181
rect 23473 21176 25655 21178
rect 23473 21120 23478 21176
rect 23534 21120 25594 21176
rect 25650 21120 25655 21176
rect 23473 21118 25655 21120
rect 23473 21115 23539 21118
rect 25589 21115 25655 21118
rect 12617 20906 12683 20909
rect 15929 20906 15995 20909
rect 12617 20904 15995 20906
rect 12617 20848 12622 20904
rect 12678 20848 15934 20904
rect 15990 20848 15995 20904
rect 12617 20846 15995 20848
rect 12617 20843 12683 20846
rect 15929 20843 15995 20846
rect 16297 20772 16363 20773
rect 16246 20708 16252 20772
rect 16316 20770 16363 20772
rect 16316 20768 16408 20770
rect 16358 20712 16408 20768
rect 16316 20710 16408 20712
rect 16316 20708 16363 20710
rect 16297 20707 16363 20708
rect 8028 20704 8344 20705
rect 8028 20640 8034 20704
rect 8098 20640 8114 20704
rect 8178 20640 8194 20704
rect 8258 20640 8274 20704
rect 8338 20640 8344 20704
rect 8028 20639 8344 20640
rect 15111 20704 15427 20705
rect 15111 20640 15117 20704
rect 15181 20640 15197 20704
rect 15261 20640 15277 20704
rect 15341 20640 15357 20704
rect 15421 20640 15427 20704
rect 15111 20639 15427 20640
rect 22194 20704 22510 20705
rect 22194 20640 22200 20704
rect 22264 20640 22280 20704
rect 22344 20640 22360 20704
rect 22424 20640 22440 20704
rect 22504 20640 22510 20704
rect 22194 20639 22510 20640
rect 29277 20704 29593 20705
rect 29277 20640 29283 20704
rect 29347 20640 29363 20704
rect 29427 20640 29443 20704
rect 29507 20640 29523 20704
rect 29587 20640 29593 20704
rect 29277 20639 29593 20640
rect 11237 20634 11303 20637
rect 13905 20634 13971 20637
rect 11237 20632 13971 20634
rect 11237 20576 11242 20632
rect 11298 20576 13910 20632
rect 13966 20576 13971 20632
rect 11237 20574 13971 20576
rect 11237 20571 11303 20574
rect 13905 20571 13971 20574
rect 4889 20362 4955 20365
rect 9857 20362 9923 20365
rect 4889 20360 9923 20362
rect 4889 20304 4894 20360
rect 4950 20304 9862 20360
rect 9918 20304 9923 20360
rect 4889 20302 9923 20304
rect 4889 20299 4955 20302
rect 9857 20299 9923 20302
rect 4487 20160 4803 20161
rect 4487 20096 4493 20160
rect 4557 20096 4573 20160
rect 4637 20096 4653 20160
rect 4717 20096 4733 20160
rect 4797 20096 4803 20160
rect 4487 20095 4803 20096
rect 11570 20160 11886 20161
rect 11570 20096 11576 20160
rect 11640 20096 11656 20160
rect 11720 20096 11736 20160
rect 11800 20096 11816 20160
rect 11880 20096 11886 20160
rect 11570 20095 11886 20096
rect 18653 20160 18969 20161
rect 18653 20096 18659 20160
rect 18723 20096 18739 20160
rect 18803 20096 18819 20160
rect 18883 20096 18899 20160
rect 18963 20096 18969 20160
rect 18653 20095 18969 20096
rect 25736 20160 26052 20161
rect 25736 20096 25742 20160
rect 25806 20096 25822 20160
rect 25886 20096 25902 20160
rect 25966 20096 25982 20160
rect 26046 20096 26052 20160
rect 25736 20095 26052 20096
rect 10409 19954 10475 19957
rect 16941 19954 17007 19957
rect 10409 19952 17007 19954
rect 10409 19896 10414 19952
rect 10470 19896 16946 19952
rect 17002 19896 17007 19952
rect 10409 19894 17007 19896
rect 10409 19891 10475 19894
rect 16941 19891 17007 19894
rect 0 19818 800 19848
rect 12065 19818 12131 19821
rect 14273 19818 14339 19821
rect 0 19728 858 19818
rect 12065 19816 14339 19818
rect 12065 19760 12070 19816
rect 12126 19760 14278 19816
rect 14334 19760 14339 19816
rect 12065 19758 14339 19760
rect 12065 19755 12131 19758
rect 14273 19755 14339 19758
rect 798 19546 858 19728
rect 8028 19616 8344 19617
rect 8028 19552 8034 19616
rect 8098 19552 8114 19616
rect 8178 19552 8194 19616
rect 8258 19552 8274 19616
rect 8338 19552 8344 19616
rect 8028 19551 8344 19552
rect 15111 19616 15427 19617
rect 15111 19552 15117 19616
rect 15181 19552 15197 19616
rect 15261 19552 15277 19616
rect 15341 19552 15357 19616
rect 15421 19552 15427 19616
rect 15111 19551 15427 19552
rect 22194 19616 22510 19617
rect 22194 19552 22200 19616
rect 22264 19552 22280 19616
rect 22344 19552 22360 19616
rect 22424 19552 22440 19616
rect 22504 19552 22510 19616
rect 22194 19551 22510 19552
rect 29277 19616 29593 19617
rect 29277 19552 29283 19616
rect 29347 19552 29363 19616
rect 29427 19552 29443 19616
rect 29507 19552 29523 19616
rect 29587 19552 29593 19616
rect 29277 19551 29593 19552
rect 1577 19546 1643 19549
rect 798 19544 1643 19546
rect 798 19488 1582 19544
rect 1638 19488 1643 19544
rect 798 19486 1643 19488
rect 1577 19483 1643 19486
rect 10133 19412 10199 19413
rect 10133 19410 10180 19412
rect 10088 19408 10180 19410
rect 10244 19410 10250 19412
rect 14917 19410 14983 19413
rect 10244 19408 14983 19410
rect 10088 19352 10138 19408
rect 10244 19352 14922 19408
rect 14978 19352 14983 19408
rect 10088 19350 10180 19352
rect 10133 19348 10180 19350
rect 10244 19350 14983 19352
rect 10244 19348 10250 19350
rect 10133 19347 10199 19348
rect 14917 19347 14983 19350
rect 4487 19072 4803 19073
rect 4487 19008 4493 19072
rect 4557 19008 4573 19072
rect 4637 19008 4653 19072
rect 4717 19008 4733 19072
rect 4797 19008 4803 19072
rect 4487 19007 4803 19008
rect 11570 19072 11886 19073
rect 11570 19008 11576 19072
rect 11640 19008 11656 19072
rect 11720 19008 11736 19072
rect 11800 19008 11816 19072
rect 11880 19008 11886 19072
rect 11570 19007 11886 19008
rect 18653 19072 18969 19073
rect 18653 19008 18659 19072
rect 18723 19008 18739 19072
rect 18803 19008 18819 19072
rect 18883 19008 18899 19072
rect 18963 19008 18969 19072
rect 18653 19007 18969 19008
rect 25736 19072 26052 19073
rect 25736 19008 25742 19072
rect 25806 19008 25822 19072
rect 25886 19008 25902 19072
rect 25966 19008 25982 19072
rect 26046 19008 26052 19072
rect 25736 19007 26052 19008
rect 29453 18730 29519 18733
rect 29453 18728 29930 18730
rect 29453 18672 29458 18728
rect 29514 18672 29930 18728
rect 29453 18670 29930 18672
rect 29453 18667 29519 18670
rect 8028 18528 8344 18529
rect 8028 18464 8034 18528
rect 8098 18464 8114 18528
rect 8178 18464 8194 18528
rect 8258 18464 8274 18528
rect 8338 18464 8344 18528
rect 8028 18463 8344 18464
rect 15111 18528 15427 18529
rect 15111 18464 15117 18528
rect 15181 18464 15197 18528
rect 15261 18464 15277 18528
rect 15341 18464 15357 18528
rect 15421 18464 15427 18528
rect 15111 18463 15427 18464
rect 22194 18528 22510 18529
rect 22194 18464 22200 18528
rect 22264 18464 22280 18528
rect 22344 18464 22360 18528
rect 22424 18464 22440 18528
rect 22504 18464 22510 18528
rect 22194 18463 22510 18464
rect 29277 18528 29593 18529
rect 29277 18464 29283 18528
rect 29347 18464 29363 18528
rect 29427 18464 29443 18528
rect 29507 18464 29523 18528
rect 29587 18464 29593 18528
rect 29870 18488 29930 18670
rect 29277 18463 29593 18464
rect 29781 18368 30581 18488
rect 4487 17984 4803 17985
rect 4487 17920 4493 17984
rect 4557 17920 4573 17984
rect 4637 17920 4653 17984
rect 4717 17920 4733 17984
rect 4797 17920 4803 17984
rect 4487 17919 4803 17920
rect 11570 17984 11886 17985
rect 11570 17920 11576 17984
rect 11640 17920 11656 17984
rect 11720 17920 11736 17984
rect 11800 17920 11816 17984
rect 11880 17920 11886 17984
rect 11570 17919 11886 17920
rect 18653 17984 18969 17985
rect 18653 17920 18659 17984
rect 18723 17920 18739 17984
rect 18803 17920 18819 17984
rect 18883 17920 18899 17984
rect 18963 17920 18969 17984
rect 18653 17919 18969 17920
rect 25736 17984 26052 17985
rect 25736 17920 25742 17984
rect 25806 17920 25822 17984
rect 25886 17920 25902 17984
rect 25966 17920 25982 17984
rect 26046 17920 26052 17984
rect 25736 17919 26052 17920
rect 15193 17914 15259 17917
rect 18413 17914 18479 17917
rect 15193 17912 18479 17914
rect 15193 17856 15198 17912
rect 15254 17856 18418 17912
rect 18474 17856 18479 17912
rect 15193 17854 18479 17856
rect 15193 17851 15259 17854
rect 18413 17851 18479 17854
rect 20253 17778 20319 17781
rect 26141 17778 26207 17781
rect 20253 17776 26207 17778
rect 20253 17720 20258 17776
rect 20314 17720 26146 17776
rect 26202 17720 26207 17776
rect 20253 17718 26207 17720
rect 20253 17715 20319 17718
rect 26141 17715 26207 17718
rect 7097 17642 7163 17645
rect 19425 17642 19491 17645
rect 7097 17640 19491 17642
rect 7097 17584 7102 17640
rect 7158 17584 19430 17640
rect 19486 17584 19491 17640
rect 7097 17582 19491 17584
rect 7097 17579 7163 17582
rect 19425 17579 19491 17582
rect 26693 17642 26759 17645
rect 27521 17642 27587 17645
rect 26693 17640 27587 17642
rect 26693 17584 26698 17640
rect 26754 17584 27526 17640
rect 27582 17584 27587 17640
rect 26693 17582 27587 17584
rect 26693 17579 26759 17582
rect 27521 17579 27587 17582
rect 8028 17440 8344 17441
rect 8028 17376 8034 17440
rect 8098 17376 8114 17440
rect 8178 17376 8194 17440
rect 8258 17376 8274 17440
rect 8338 17376 8344 17440
rect 8028 17375 8344 17376
rect 15111 17440 15427 17441
rect 15111 17376 15117 17440
rect 15181 17376 15197 17440
rect 15261 17376 15277 17440
rect 15341 17376 15357 17440
rect 15421 17376 15427 17440
rect 15111 17375 15427 17376
rect 22194 17440 22510 17441
rect 22194 17376 22200 17440
rect 22264 17376 22280 17440
rect 22344 17376 22360 17440
rect 22424 17376 22440 17440
rect 22504 17376 22510 17440
rect 22194 17375 22510 17376
rect 29277 17440 29593 17441
rect 29277 17376 29283 17440
rect 29347 17376 29363 17440
rect 29427 17376 29443 17440
rect 29507 17376 29523 17440
rect 29587 17376 29593 17440
rect 29277 17375 29593 17376
rect 26049 17234 26115 17237
rect 27245 17234 27311 17237
rect 27705 17236 27771 17237
rect 26049 17232 27311 17234
rect 26049 17176 26054 17232
rect 26110 17176 27250 17232
rect 27306 17176 27311 17232
rect 26049 17174 27311 17176
rect 26049 17171 26115 17174
rect 27245 17171 27311 17174
rect 27654 17172 27660 17236
rect 27724 17234 27771 17236
rect 27724 17232 27816 17234
rect 27766 17176 27816 17232
rect 27724 17174 27816 17176
rect 27724 17172 27771 17174
rect 27705 17171 27771 17172
rect 4613 17098 4679 17101
rect 5257 17098 5323 17101
rect 4613 17096 5323 17098
rect 4613 17040 4618 17096
rect 4674 17040 5262 17096
rect 5318 17040 5323 17096
rect 4613 17038 5323 17040
rect 4613 17035 4679 17038
rect 5257 17035 5323 17038
rect 4487 16896 4803 16897
rect 4487 16832 4493 16896
rect 4557 16832 4573 16896
rect 4637 16832 4653 16896
rect 4717 16832 4733 16896
rect 4797 16832 4803 16896
rect 4487 16831 4803 16832
rect 11570 16896 11886 16897
rect 11570 16832 11576 16896
rect 11640 16832 11656 16896
rect 11720 16832 11736 16896
rect 11800 16832 11816 16896
rect 11880 16832 11886 16896
rect 11570 16831 11886 16832
rect 18653 16896 18969 16897
rect 18653 16832 18659 16896
rect 18723 16832 18739 16896
rect 18803 16832 18819 16896
rect 18883 16832 18899 16896
rect 18963 16832 18969 16896
rect 18653 16831 18969 16832
rect 25736 16896 26052 16897
rect 25736 16832 25742 16896
rect 25806 16832 25822 16896
rect 25886 16832 25902 16896
rect 25966 16832 25982 16896
rect 26046 16832 26052 16896
rect 25736 16831 26052 16832
rect 26049 16418 26115 16421
rect 27981 16418 28047 16421
rect 26049 16416 28047 16418
rect 26049 16360 26054 16416
rect 26110 16360 27986 16416
rect 28042 16360 28047 16416
rect 26049 16358 28047 16360
rect 26049 16355 26115 16358
rect 27981 16355 28047 16358
rect 8028 16352 8344 16353
rect 8028 16288 8034 16352
rect 8098 16288 8114 16352
rect 8178 16288 8194 16352
rect 8258 16288 8274 16352
rect 8338 16288 8344 16352
rect 8028 16287 8344 16288
rect 15111 16352 15427 16353
rect 15111 16288 15117 16352
rect 15181 16288 15197 16352
rect 15261 16288 15277 16352
rect 15341 16288 15357 16352
rect 15421 16288 15427 16352
rect 15111 16287 15427 16288
rect 22194 16352 22510 16353
rect 22194 16288 22200 16352
rect 22264 16288 22280 16352
rect 22344 16288 22360 16352
rect 22424 16288 22440 16352
rect 22504 16288 22510 16352
rect 22194 16287 22510 16288
rect 29277 16352 29593 16353
rect 29277 16288 29283 16352
rect 29347 16288 29363 16352
rect 29427 16288 29443 16352
rect 29507 16288 29523 16352
rect 29587 16288 29593 16352
rect 29277 16287 29593 16288
rect 4487 15808 4803 15809
rect 0 15738 800 15768
rect 4487 15744 4493 15808
rect 4557 15744 4573 15808
rect 4637 15744 4653 15808
rect 4717 15744 4733 15808
rect 4797 15744 4803 15808
rect 4487 15743 4803 15744
rect 11570 15808 11886 15809
rect 11570 15744 11576 15808
rect 11640 15744 11656 15808
rect 11720 15744 11736 15808
rect 11800 15744 11816 15808
rect 11880 15744 11886 15808
rect 11570 15743 11886 15744
rect 18653 15808 18969 15809
rect 18653 15744 18659 15808
rect 18723 15744 18739 15808
rect 18803 15744 18819 15808
rect 18883 15744 18899 15808
rect 18963 15744 18969 15808
rect 18653 15743 18969 15744
rect 25736 15808 26052 15809
rect 25736 15744 25742 15808
rect 25806 15744 25822 15808
rect 25886 15744 25902 15808
rect 25966 15744 25982 15808
rect 26046 15744 26052 15808
rect 25736 15743 26052 15744
rect 933 15738 999 15741
rect 0 15736 999 15738
rect 0 15680 938 15736
rect 994 15680 999 15736
rect 0 15678 999 15680
rect 0 15648 800 15678
rect 933 15675 999 15678
rect 10501 15602 10567 15605
rect 17953 15602 18019 15605
rect 10501 15600 18019 15602
rect 10501 15544 10506 15600
rect 10562 15544 17958 15600
rect 18014 15544 18019 15600
rect 10501 15542 18019 15544
rect 10501 15539 10567 15542
rect 17953 15539 18019 15542
rect 4061 15466 4127 15469
rect 6637 15466 6703 15469
rect 4061 15464 6703 15466
rect 4061 15408 4066 15464
rect 4122 15408 6642 15464
rect 6698 15408 6703 15464
rect 4061 15406 6703 15408
rect 4061 15403 4127 15406
rect 6637 15403 6703 15406
rect 25129 15466 25195 15469
rect 26509 15466 26575 15469
rect 25129 15464 26575 15466
rect 25129 15408 25134 15464
rect 25190 15408 26514 15464
rect 26570 15408 26575 15464
rect 25129 15406 26575 15408
rect 25129 15403 25195 15406
rect 26509 15403 26575 15406
rect 8028 15264 8344 15265
rect 8028 15200 8034 15264
rect 8098 15200 8114 15264
rect 8178 15200 8194 15264
rect 8258 15200 8274 15264
rect 8338 15200 8344 15264
rect 8028 15199 8344 15200
rect 15111 15264 15427 15265
rect 15111 15200 15117 15264
rect 15181 15200 15197 15264
rect 15261 15200 15277 15264
rect 15341 15200 15357 15264
rect 15421 15200 15427 15264
rect 15111 15199 15427 15200
rect 22194 15264 22510 15265
rect 22194 15200 22200 15264
rect 22264 15200 22280 15264
rect 22344 15200 22360 15264
rect 22424 15200 22440 15264
rect 22504 15200 22510 15264
rect 22194 15199 22510 15200
rect 29277 15264 29593 15265
rect 29277 15200 29283 15264
rect 29347 15200 29363 15264
rect 29427 15200 29443 15264
rect 29507 15200 29523 15264
rect 29587 15200 29593 15264
rect 29277 15199 29593 15200
rect 16297 15196 16363 15197
rect 16246 15194 16252 15196
rect 16206 15134 16252 15194
rect 16316 15192 16363 15196
rect 16358 15136 16363 15192
rect 16246 15132 16252 15134
rect 16316 15132 16363 15136
rect 16297 15131 16363 15132
rect 4487 14720 4803 14721
rect 4487 14656 4493 14720
rect 4557 14656 4573 14720
rect 4637 14656 4653 14720
rect 4717 14656 4733 14720
rect 4797 14656 4803 14720
rect 4487 14655 4803 14656
rect 11570 14720 11886 14721
rect 11570 14656 11576 14720
rect 11640 14656 11656 14720
rect 11720 14656 11736 14720
rect 11800 14656 11816 14720
rect 11880 14656 11886 14720
rect 11570 14655 11886 14656
rect 18653 14720 18969 14721
rect 18653 14656 18659 14720
rect 18723 14656 18739 14720
rect 18803 14656 18819 14720
rect 18883 14656 18899 14720
rect 18963 14656 18969 14720
rect 18653 14655 18969 14656
rect 25736 14720 26052 14721
rect 25736 14656 25742 14720
rect 25806 14656 25822 14720
rect 25886 14656 25902 14720
rect 25966 14656 25982 14720
rect 26046 14656 26052 14720
rect 25736 14655 26052 14656
rect 28993 14378 29059 14381
rect 29781 14378 30581 14408
rect 28993 14376 30581 14378
rect 28993 14320 28998 14376
rect 29054 14320 30581 14376
rect 28993 14318 30581 14320
rect 28993 14315 29059 14318
rect 29781 14288 30581 14318
rect 8028 14176 8344 14177
rect 8028 14112 8034 14176
rect 8098 14112 8114 14176
rect 8178 14112 8194 14176
rect 8258 14112 8274 14176
rect 8338 14112 8344 14176
rect 8028 14111 8344 14112
rect 15111 14176 15427 14177
rect 15111 14112 15117 14176
rect 15181 14112 15197 14176
rect 15261 14112 15277 14176
rect 15341 14112 15357 14176
rect 15421 14112 15427 14176
rect 15111 14111 15427 14112
rect 22194 14176 22510 14177
rect 22194 14112 22200 14176
rect 22264 14112 22280 14176
rect 22344 14112 22360 14176
rect 22424 14112 22440 14176
rect 22504 14112 22510 14176
rect 22194 14111 22510 14112
rect 29277 14176 29593 14177
rect 29277 14112 29283 14176
rect 29347 14112 29363 14176
rect 29427 14112 29443 14176
rect 29507 14112 29523 14176
rect 29587 14112 29593 14176
rect 29277 14111 29593 14112
rect 10133 13970 10199 13973
rect 12341 13970 12407 13973
rect 10133 13968 12407 13970
rect 10133 13912 10138 13968
rect 10194 13912 12346 13968
rect 12402 13912 12407 13968
rect 10133 13910 12407 13912
rect 10133 13907 10199 13910
rect 12341 13907 12407 13910
rect 19057 13834 19123 13837
rect 20161 13834 20227 13837
rect 19057 13832 20227 13834
rect 19057 13776 19062 13832
rect 19118 13776 20166 13832
rect 20222 13776 20227 13832
rect 19057 13774 20227 13776
rect 19057 13771 19123 13774
rect 20161 13771 20227 13774
rect 4487 13632 4803 13633
rect 4487 13568 4493 13632
rect 4557 13568 4573 13632
rect 4637 13568 4653 13632
rect 4717 13568 4733 13632
rect 4797 13568 4803 13632
rect 4487 13567 4803 13568
rect 11570 13632 11886 13633
rect 11570 13568 11576 13632
rect 11640 13568 11656 13632
rect 11720 13568 11736 13632
rect 11800 13568 11816 13632
rect 11880 13568 11886 13632
rect 11570 13567 11886 13568
rect 18653 13632 18969 13633
rect 18653 13568 18659 13632
rect 18723 13568 18739 13632
rect 18803 13568 18819 13632
rect 18883 13568 18899 13632
rect 18963 13568 18969 13632
rect 18653 13567 18969 13568
rect 25736 13632 26052 13633
rect 25736 13568 25742 13632
rect 25806 13568 25822 13632
rect 25886 13568 25902 13632
rect 25966 13568 25982 13632
rect 26046 13568 26052 13632
rect 25736 13567 26052 13568
rect 9673 13426 9739 13429
rect 9673 13424 10610 13426
rect 9673 13368 9678 13424
rect 9734 13368 10610 13424
rect 9673 13366 10610 13368
rect 9673 13363 9739 13366
rect 10550 13292 10610 13366
rect 10542 13228 10548 13292
rect 10612 13290 10618 13292
rect 11513 13290 11579 13293
rect 10612 13288 11579 13290
rect 10612 13232 11518 13288
rect 11574 13232 11579 13288
rect 10612 13230 11579 13232
rect 10612 13228 10618 13230
rect 11513 13227 11579 13230
rect 8028 13088 8344 13089
rect 8028 13024 8034 13088
rect 8098 13024 8114 13088
rect 8178 13024 8194 13088
rect 8258 13024 8274 13088
rect 8338 13024 8344 13088
rect 8028 13023 8344 13024
rect 15111 13088 15427 13089
rect 15111 13024 15117 13088
rect 15181 13024 15197 13088
rect 15261 13024 15277 13088
rect 15341 13024 15357 13088
rect 15421 13024 15427 13088
rect 15111 13023 15427 13024
rect 22194 13088 22510 13089
rect 22194 13024 22200 13088
rect 22264 13024 22280 13088
rect 22344 13024 22360 13088
rect 22424 13024 22440 13088
rect 22504 13024 22510 13088
rect 22194 13023 22510 13024
rect 29277 13088 29593 13089
rect 29277 13024 29283 13088
rect 29347 13024 29363 13088
rect 29427 13024 29443 13088
rect 29507 13024 29523 13088
rect 29587 13024 29593 13088
rect 29277 13023 29593 13024
rect 4487 12544 4803 12545
rect 4487 12480 4493 12544
rect 4557 12480 4573 12544
rect 4637 12480 4653 12544
rect 4717 12480 4733 12544
rect 4797 12480 4803 12544
rect 4487 12479 4803 12480
rect 11570 12544 11886 12545
rect 11570 12480 11576 12544
rect 11640 12480 11656 12544
rect 11720 12480 11736 12544
rect 11800 12480 11816 12544
rect 11880 12480 11886 12544
rect 11570 12479 11886 12480
rect 18653 12544 18969 12545
rect 18653 12480 18659 12544
rect 18723 12480 18739 12544
rect 18803 12480 18819 12544
rect 18883 12480 18899 12544
rect 18963 12480 18969 12544
rect 18653 12479 18969 12480
rect 25736 12544 26052 12545
rect 25736 12480 25742 12544
rect 25806 12480 25822 12544
rect 25886 12480 25902 12544
rect 25966 12480 25982 12544
rect 26046 12480 26052 12544
rect 25736 12479 26052 12480
rect 3049 12338 3115 12341
rect 14273 12338 14339 12341
rect 16665 12338 16731 12341
rect 19149 12338 19215 12341
rect 22829 12338 22895 12341
rect 3049 12336 16731 12338
rect 3049 12280 3054 12336
rect 3110 12280 14278 12336
rect 14334 12280 16670 12336
rect 16726 12280 16731 12336
rect 3049 12278 16731 12280
rect 3049 12275 3115 12278
rect 14273 12275 14339 12278
rect 16665 12275 16731 12278
rect 16806 12336 22895 12338
rect 16806 12280 19154 12336
rect 19210 12280 22834 12336
rect 22890 12280 22895 12336
rect 16806 12278 22895 12280
rect 3785 12202 3851 12205
rect 5165 12202 5231 12205
rect 10409 12202 10475 12205
rect 3785 12200 10475 12202
rect 3785 12144 3790 12200
rect 3846 12144 5170 12200
rect 5226 12144 10414 12200
rect 10470 12144 10475 12200
rect 3785 12142 10475 12144
rect 3785 12139 3851 12142
rect 5165 12139 5231 12142
rect 10409 12139 10475 12142
rect 14089 12202 14155 12205
rect 16806 12202 16866 12278
rect 19149 12275 19215 12278
rect 22829 12275 22895 12278
rect 14089 12200 16866 12202
rect 14089 12144 14094 12200
rect 14150 12144 16866 12200
rect 14089 12142 16866 12144
rect 14089 12139 14155 12142
rect 8028 12000 8344 12001
rect 8028 11936 8034 12000
rect 8098 11936 8114 12000
rect 8178 11936 8194 12000
rect 8258 11936 8274 12000
rect 8338 11936 8344 12000
rect 8028 11935 8344 11936
rect 15111 12000 15427 12001
rect 15111 11936 15117 12000
rect 15181 11936 15197 12000
rect 15261 11936 15277 12000
rect 15341 11936 15357 12000
rect 15421 11936 15427 12000
rect 15111 11935 15427 11936
rect 22194 12000 22510 12001
rect 22194 11936 22200 12000
rect 22264 11936 22280 12000
rect 22344 11936 22360 12000
rect 22424 11936 22440 12000
rect 22504 11936 22510 12000
rect 22194 11935 22510 11936
rect 29277 12000 29593 12001
rect 29277 11936 29283 12000
rect 29347 11936 29363 12000
rect 29427 11936 29443 12000
rect 29507 11936 29523 12000
rect 29587 11936 29593 12000
rect 29277 11935 29593 11936
rect 2221 11794 2287 11797
rect 27654 11794 27660 11796
rect 2221 11792 27660 11794
rect 2221 11736 2226 11792
rect 2282 11736 27660 11792
rect 2221 11734 27660 11736
rect 2221 11731 2287 11734
rect 27654 11732 27660 11734
rect 27724 11732 27730 11796
rect 0 11658 800 11688
rect 933 11658 999 11661
rect 0 11656 999 11658
rect 0 11600 938 11656
rect 994 11600 999 11656
rect 0 11598 999 11600
rect 0 11568 800 11598
rect 933 11595 999 11598
rect 4487 11456 4803 11457
rect 4487 11392 4493 11456
rect 4557 11392 4573 11456
rect 4637 11392 4653 11456
rect 4717 11392 4733 11456
rect 4797 11392 4803 11456
rect 4487 11391 4803 11392
rect 11570 11456 11886 11457
rect 11570 11392 11576 11456
rect 11640 11392 11656 11456
rect 11720 11392 11736 11456
rect 11800 11392 11816 11456
rect 11880 11392 11886 11456
rect 11570 11391 11886 11392
rect 18653 11456 18969 11457
rect 18653 11392 18659 11456
rect 18723 11392 18739 11456
rect 18803 11392 18819 11456
rect 18883 11392 18899 11456
rect 18963 11392 18969 11456
rect 18653 11391 18969 11392
rect 25736 11456 26052 11457
rect 25736 11392 25742 11456
rect 25806 11392 25822 11456
rect 25886 11392 25902 11456
rect 25966 11392 25982 11456
rect 26046 11392 26052 11456
rect 25736 11391 26052 11392
rect 13261 11114 13327 11117
rect 18689 11114 18755 11117
rect 13261 11112 18755 11114
rect 13261 11056 13266 11112
rect 13322 11056 18694 11112
rect 18750 11056 18755 11112
rect 13261 11054 18755 11056
rect 13261 11051 13327 11054
rect 18689 11051 18755 11054
rect 21541 11114 21607 11117
rect 24393 11114 24459 11117
rect 21541 11112 24459 11114
rect 21541 11056 21546 11112
rect 21602 11056 24398 11112
rect 24454 11056 24459 11112
rect 21541 11054 24459 11056
rect 21541 11051 21607 11054
rect 24393 11051 24459 11054
rect 29085 11114 29151 11117
rect 29085 11112 29746 11114
rect 29085 11056 29090 11112
rect 29146 11056 29746 11112
rect 29085 11054 29746 11056
rect 29085 11051 29151 11054
rect 29686 11012 29746 11054
rect 29686 11008 29930 11012
rect 29686 10952 30581 11008
rect 8028 10912 8344 10913
rect 8028 10848 8034 10912
rect 8098 10848 8114 10912
rect 8178 10848 8194 10912
rect 8258 10848 8274 10912
rect 8338 10848 8344 10912
rect 8028 10847 8344 10848
rect 15111 10912 15427 10913
rect 15111 10848 15117 10912
rect 15181 10848 15197 10912
rect 15261 10848 15277 10912
rect 15341 10848 15357 10912
rect 15421 10848 15427 10912
rect 15111 10847 15427 10848
rect 22194 10912 22510 10913
rect 22194 10848 22200 10912
rect 22264 10848 22280 10912
rect 22344 10848 22360 10912
rect 22424 10848 22440 10912
rect 22504 10848 22510 10912
rect 22194 10847 22510 10848
rect 29277 10912 29593 10913
rect 29277 10848 29283 10912
rect 29347 10848 29363 10912
rect 29427 10848 29443 10912
rect 29507 10848 29523 10912
rect 29587 10848 29593 10912
rect 29781 10888 30581 10952
rect 29277 10847 29593 10848
rect 4487 10368 4803 10369
rect 4487 10304 4493 10368
rect 4557 10304 4573 10368
rect 4637 10304 4653 10368
rect 4717 10304 4733 10368
rect 4797 10304 4803 10368
rect 4487 10303 4803 10304
rect 11570 10368 11886 10369
rect 11570 10304 11576 10368
rect 11640 10304 11656 10368
rect 11720 10304 11736 10368
rect 11800 10304 11816 10368
rect 11880 10304 11886 10368
rect 11570 10303 11886 10304
rect 18653 10368 18969 10369
rect 18653 10304 18659 10368
rect 18723 10304 18739 10368
rect 18803 10304 18819 10368
rect 18883 10304 18899 10368
rect 18963 10304 18969 10368
rect 18653 10303 18969 10304
rect 25736 10368 26052 10369
rect 25736 10304 25742 10368
rect 25806 10304 25822 10368
rect 25886 10304 25902 10368
rect 25966 10304 25982 10368
rect 26046 10304 26052 10368
rect 25736 10303 26052 10304
rect 19885 10162 19951 10165
rect 22645 10162 22711 10165
rect 19885 10160 22711 10162
rect 19885 10104 19890 10160
rect 19946 10104 22650 10160
rect 22706 10104 22711 10160
rect 19885 10102 22711 10104
rect 19885 10099 19951 10102
rect 22645 10099 22711 10102
rect 8028 9824 8344 9825
rect 8028 9760 8034 9824
rect 8098 9760 8114 9824
rect 8178 9760 8194 9824
rect 8258 9760 8274 9824
rect 8338 9760 8344 9824
rect 8028 9759 8344 9760
rect 15111 9824 15427 9825
rect 15111 9760 15117 9824
rect 15181 9760 15197 9824
rect 15261 9760 15277 9824
rect 15341 9760 15357 9824
rect 15421 9760 15427 9824
rect 15111 9759 15427 9760
rect 22194 9824 22510 9825
rect 22194 9760 22200 9824
rect 22264 9760 22280 9824
rect 22344 9760 22360 9824
rect 22424 9760 22440 9824
rect 22504 9760 22510 9824
rect 22194 9759 22510 9760
rect 29277 9824 29593 9825
rect 29277 9760 29283 9824
rect 29347 9760 29363 9824
rect 29427 9760 29443 9824
rect 29507 9760 29523 9824
rect 29587 9760 29593 9824
rect 29277 9759 29593 9760
rect 10317 9754 10383 9757
rect 10869 9754 10935 9757
rect 11145 9754 11211 9757
rect 10317 9752 11211 9754
rect 10317 9696 10322 9752
rect 10378 9696 10874 9752
rect 10930 9696 11150 9752
rect 11206 9696 11211 9752
rect 10317 9694 11211 9696
rect 10317 9691 10383 9694
rect 10869 9691 10935 9694
rect 11145 9691 11211 9694
rect 5441 9618 5507 9621
rect 12249 9618 12315 9621
rect 5441 9616 12315 9618
rect 5441 9560 5446 9616
rect 5502 9560 12254 9616
rect 12310 9560 12315 9616
rect 5441 9558 12315 9560
rect 5441 9555 5507 9558
rect 12249 9555 12315 9558
rect 13169 9618 13235 9621
rect 16021 9618 16087 9621
rect 17033 9618 17099 9621
rect 13169 9616 17099 9618
rect 13169 9560 13174 9616
rect 13230 9560 16026 9616
rect 16082 9560 17038 9616
rect 17094 9560 17099 9616
rect 13169 9558 17099 9560
rect 13169 9555 13235 9558
rect 16021 9555 16087 9558
rect 17033 9555 17099 9558
rect 4061 9482 4127 9485
rect 6913 9482 6979 9485
rect 4061 9480 6979 9482
rect 4061 9424 4066 9480
rect 4122 9424 6918 9480
rect 6974 9424 6979 9480
rect 4061 9422 6979 9424
rect 4061 9419 4127 9422
rect 6913 9419 6979 9422
rect 8845 9482 8911 9485
rect 10174 9482 10180 9484
rect 8845 9480 10180 9482
rect 8845 9424 8850 9480
rect 8906 9424 10180 9480
rect 8845 9422 10180 9424
rect 8845 9419 8911 9422
rect 10174 9420 10180 9422
rect 10244 9482 10250 9484
rect 17125 9482 17191 9485
rect 10244 9480 17191 9482
rect 10244 9424 17130 9480
rect 17186 9424 17191 9480
rect 10244 9422 17191 9424
rect 10244 9420 10250 9422
rect 17125 9419 17191 9422
rect 9765 9346 9831 9349
rect 10317 9346 10383 9349
rect 9765 9344 10383 9346
rect 9765 9288 9770 9344
rect 9826 9288 10322 9344
rect 10378 9288 10383 9344
rect 9765 9286 10383 9288
rect 9765 9283 9831 9286
rect 10317 9283 10383 9286
rect 4487 9280 4803 9281
rect 4487 9216 4493 9280
rect 4557 9216 4573 9280
rect 4637 9216 4653 9280
rect 4717 9216 4733 9280
rect 4797 9216 4803 9280
rect 4487 9215 4803 9216
rect 11570 9280 11886 9281
rect 11570 9216 11576 9280
rect 11640 9216 11656 9280
rect 11720 9216 11736 9280
rect 11800 9216 11816 9280
rect 11880 9216 11886 9280
rect 11570 9215 11886 9216
rect 18653 9280 18969 9281
rect 18653 9216 18659 9280
rect 18723 9216 18739 9280
rect 18803 9216 18819 9280
rect 18883 9216 18899 9280
rect 18963 9216 18969 9280
rect 18653 9215 18969 9216
rect 25736 9280 26052 9281
rect 25736 9216 25742 9280
rect 25806 9216 25822 9280
rect 25886 9216 25902 9280
rect 25966 9216 25982 9280
rect 26046 9216 26052 9280
rect 25736 9215 26052 9216
rect 8028 8736 8344 8737
rect 8028 8672 8034 8736
rect 8098 8672 8114 8736
rect 8178 8672 8194 8736
rect 8258 8672 8274 8736
rect 8338 8672 8344 8736
rect 8028 8671 8344 8672
rect 15111 8736 15427 8737
rect 15111 8672 15117 8736
rect 15181 8672 15197 8736
rect 15261 8672 15277 8736
rect 15341 8672 15357 8736
rect 15421 8672 15427 8736
rect 15111 8671 15427 8672
rect 22194 8736 22510 8737
rect 22194 8672 22200 8736
rect 22264 8672 22280 8736
rect 22344 8672 22360 8736
rect 22424 8672 22440 8736
rect 22504 8672 22510 8736
rect 22194 8671 22510 8672
rect 29277 8736 29593 8737
rect 29277 8672 29283 8736
rect 29347 8672 29363 8736
rect 29427 8672 29443 8736
rect 29507 8672 29523 8736
rect 29587 8672 29593 8736
rect 29277 8671 29593 8672
rect 5441 8530 5507 8533
rect 9029 8530 9095 8533
rect 5441 8528 9095 8530
rect 5441 8472 5446 8528
rect 5502 8472 9034 8528
rect 9090 8472 9095 8528
rect 5441 8470 9095 8472
rect 5441 8467 5507 8470
rect 9029 8467 9095 8470
rect 26141 8530 26207 8533
rect 27797 8530 27863 8533
rect 26141 8528 27863 8530
rect 26141 8472 26146 8528
rect 26202 8472 27802 8528
rect 27858 8472 27863 8528
rect 26141 8470 27863 8472
rect 26141 8467 26207 8470
rect 27797 8467 27863 8470
rect 10501 8260 10567 8261
rect 10501 8258 10548 8260
rect 10456 8256 10548 8258
rect 10456 8200 10506 8256
rect 10456 8198 10548 8200
rect 10501 8196 10548 8198
rect 10612 8196 10618 8260
rect 10501 8195 10567 8196
rect 4487 8192 4803 8193
rect 4487 8128 4493 8192
rect 4557 8128 4573 8192
rect 4637 8128 4653 8192
rect 4717 8128 4733 8192
rect 4797 8128 4803 8192
rect 4487 8127 4803 8128
rect 11570 8192 11886 8193
rect 11570 8128 11576 8192
rect 11640 8128 11656 8192
rect 11720 8128 11736 8192
rect 11800 8128 11816 8192
rect 11880 8128 11886 8192
rect 11570 8127 11886 8128
rect 18653 8192 18969 8193
rect 18653 8128 18659 8192
rect 18723 8128 18739 8192
rect 18803 8128 18819 8192
rect 18883 8128 18899 8192
rect 18963 8128 18969 8192
rect 18653 8127 18969 8128
rect 25736 8192 26052 8193
rect 25736 8128 25742 8192
rect 25806 8128 25822 8192
rect 25886 8128 25902 8192
rect 25966 8128 25982 8192
rect 26046 8128 26052 8192
rect 25736 8127 26052 8128
rect 17401 7986 17467 7989
rect 22829 7986 22895 7989
rect 17401 7984 22895 7986
rect 17401 7928 17406 7984
rect 17462 7928 22834 7984
rect 22890 7928 22895 7984
rect 17401 7926 22895 7928
rect 17401 7923 17467 7926
rect 22829 7923 22895 7926
rect 8028 7648 8344 7649
rect 0 7578 800 7608
rect 8028 7584 8034 7648
rect 8098 7584 8114 7648
rect 8178 7584 8194 7648
rect 8258 7584 8274 7648
rect 8338 7584 8344 7648
rect 8028 7583 8344 7584
rect 15111 7648 15427 7649
rect 15111 7584 15117 7648
rect 15181 7584 15197 7648
rect 15261 7584 15277 7648
rect 15341 7584 15357 7648
rect 15421 7584 15427 7648
rect 15111 7583 15427 7584
rect 22194 7648 22510 7649
rect 22194 7584 22200 7648
rect 22264 7584 22280 7648
rect 22344 7584 22360 7648
rect 22424 7584 22440 7648
rect 22504 7584 22510 7648
rect 22194 7583 22510 7584
rect 29277 7648 29593 7649
rect 29277 7584 29283 7648
rect 29347 7584 29363 7648
rect 29427 7584 29443 7648
rect 29507 7584 29523 7648
rect 29587 7584 29593 7648
rect 29277 7583 29593 7584
rect 4061 7578 4127 7581
rect 0 7576 4127 7578
rect 0 7520 4066 7576
rect 4122 7520 4127 7576
rect 0 7518 4127 7520
rect 0 7488 800 7518
rect 4061 7515 4127 7518
rect 17217 7442 17283 7445
rect 17861 7442 17927 7445
rect 17217 7440 17927 7442
rect 17217 7384 17222 7440
rect 17278 7384 17866 7440
rect 17922 7384 17927 7440
rect 17217 7382 17927 7384
rect 17217 7379 17283 7382
rect 17861 7379 17927 7382
rect 4487 7104 4803 7105
rect 4487 7040 4493 7104
rect 4557 7040 4573 7104
rect 4637 7040 4653 7104
rect 4717 7040 4733 7104
rect 4797 7040 4803 7104
rect 4487 7039 4803 7040
rect 11570 7104 11886 7105
rect 11570 7040 11576 7104
rect 11640 7040 11656 7104
rect 11720 7040 11736 7104
rect 11800 7040 11816 7104
rect 11880 7040 11886 7104
rect 11570 7039 11886 7040
rect 18653 7104 18969 7105
rect 18653 7040 18659 7104
rect 18723 7040 18739 7104
rect 18803 7040 18819 7104
rect 18883 7040 18899 7104
rect 18963 7040 18969 7104
rect 18653 7039 18969 7040
rect 25736 7104 26052 7105
rect 25736 7040 25742 7104
rect 25806 7040 25822 7104
rect 25886 7040 25902 7104
rect 25966 7040 25982 7104
rect 26046 7040 26052 7104
rect 25736 7039 26052 7040
rect 29085 6898 29151 6901
rect 29781 6898 30581 6928
rect 29085 6896 30581 6898
rect 29085 6840 29090 6896
rect 29146 6840 30581 6896
rect 29085 6838 30581 6840
rect 29085 6835 29151 6838
rect 29781 6808 30581 6838
rect 5993 6762 6059 6765
rect 7741 6762 7807 6765
rect 5993 6760 7807 6762
rect 5993 6704 5998 6760
rect 6054 6704 7746 6760
rect 7802 6704 7807 6760
rect 5993 6702 7807 6704
rect 5993 6699 6059 6702
rect 7741 6699 7807 6702
rect 10777 6762 10843 6765
rect 14089 6762 14155 6765
rect 10777 6760 14155 6762
rect 10777 6704 10782 6760
rect 10838 6704 14094 6760
rect 14150 6704 14155 6760
rect 10777 6702 14155 6704
rect 10777 6699 10843 6702
rect 14089 6699 14155 6702
rect 20069 6762 20135 6765
rect 28758 6762 28764 6764
rect 20069 6760 28764 6762
rect 20069 6704 20074 6760
rect 20130 6704 28764 6760
rect 20069 6702 28764 6704
rect 20069 6699 20135 6702
rect 28758 6700 28764 6702
rect 28828 6700 28834 6764
rect 10961 6626 11027 6629
rect 13905 6626 13971 6629
rect 10961 6624 13971 6626
rect 10961 6568 10966 6624
rect 11022 6568 13910 6624
rect 13966 6568 13971 6624
rect 10961 6566 13971 6568
rect 10961 6563 11027 6566
rect 13905 6563 13971 6566
rect 8028 6560 8344 6561
rect 8028 6496 8034 6560
rect 8098 6496 8114 6560
rect 8178 6496 8194 6560
rect 8258 6496 8274 6560
rect 8338 6496 8344 6560
rect 8028 6495 8344 6496
rect 15111 6560 15427 6561
rect 15111 6496 15117 6560
rect 15181 6496 15197 6560
rect 15261 6496 15277 6560
rect 15341 6496 15357 6560
rect 15421 6496 15427 6560
rect 15111 6495 15427 6496
rect 22194 6560 22510 6561
rect 22194 6496 22200 6560
rect 22264 6496 22280 6560
rect 22344 6496 22360 6560
rect 22424 6496 22440 6560
rect 22504 6496 22510 6560
rect 22194 6495 22510 6496
rect 29277 6560 29593 6561
rect 29277 6496 29283 6560
rect 29347 6496 29363 6560
rect 29427 6496 29443 6560
rect 29507 6496 29523 6560
rect 29587 6496 29593 6560
rect 29277 6495 29593 6496
rect 1485 6354 1551 6357
rect 20253 6354 20319 6357
rect 1485 6352 20319 6354
rect 1485 6296 1490 6352
rect 1546 6296 20258 6352
rect 20314 6296 20319 6352
rect 1485 6294 20319 6296
rect 1485 6291 1551 6294
rect 20253 6291 20319 6294
rect 4487 6016 4803 6017
rect 4487 5952 4493 6016
rect 4557 5952 4573 6016
rect 4637 5952 4653 6016
rect 4717 5952 4733 6016
rect 4797 5952 4803 6016
rect 4487 5951 4803 5952
rect 11570 6016 11886 6017
rect 11570 5952 11576 6016
rect 11640 5952 11656 6016
rect 11720 5952 11736 6016
rect 11800 5952 11816 6016
rect 11880 5952 11886 6016
rect 11570 5951 11886 5952
rect 18653 6016 18969 6017
rect 18653 5952 18659 6016
rect 18723 5952 18739 6016
rect 18803 5952 18819 6016
rect 18883 5952 18899 6016
rect 18963 5952 18969 6016
rect 18653 5951 18969 5952
rect 25736 6016 26052 6017
rect 25736 5952 25742 6016
rect 25806 5952 25822 6016
rect 25886 5952 25902 6016
rect 25966 5952 25982 6016
rect 26046 5952 26052 6016
rect 25736 5951 26052 5952
rect 24301 5540 24367 5541
rect 24301 5538 24348 5540
rect 24256 5536 24348 5538
rect 24256 5480 24306 5536
rect 24256 5478 24348 5480
rect 24301 5476 24348 5478
rect 24412 5476 24418 5540
rect 24301 5475 24367 5476
rect 8028 5472 8344 5473
rect 8028 5408 8034 5472
rect 8098 5408 8114 5472
rect 8178 5408 8194 5472
rect 8258 5408 8274 5472
rect 8338 5408 8344 5472
rect 8028 5407 8344 5408
rect 15111 5472 15427 5473
rect 15111 5408 15117 5472
rect 15181 5408 15197 5472
rect 15261 5408 15277 5472
rect 15341 5408 15357 5472
rect 15421 5408 15427 5472
rect 15111 5407 15427 5408
rect 22194 5472 22510 5473
rect 22194 5408 22200 5472
rect 22264 5408 22280 5472
rect 22344 5408 22360 5472
rect 22424 5408 22440 5472
rect 22504 5408 22510 5472
rect 22194 5407 22510 5408
rect 29277 5472 29593 5473
rect 29277 5408 29283 5472
rect 29347 5408 29363 5472
rect 29427 5408 29443 5472
rect 29507 5408 29523 5472
rect 29587 5408 29593 5472
rect 29277 5407 29593 5408
rect 17033 5130 17099 5133
rect 18229 5130 18295 5133
rect 17033 5128 18295 5130
rect 17033 5072 17038 5128
rect 17094 5072 18234 5128
rect 18290 5072 18295 5128
rect 17033 5070 18295 5072
rect 17033 5067 17099 5070
rect 18229 5067 18295 5070
rect 16205 4994 16271 4997
rect 18321 4994 18387 4997
rect 16205 4992 18387 4994
rect 16205 4936 16210 4992
rect 16266 4936 18326 4992
rect 18382 4936 18387 4992
rect 16205 4934 18387 4936
rect 16205 4931 16271 4934
rect 18321 4931 18387 4934
rect 4487 4928 4803 4929
rect 4487 4864 4493 4928
rect 4557 4864 4573 4928
rect 4637 4864 4653 4928
rect 4717 4864 4733 4928
rect 4797 4864 4803 4928
rect 4487 4863 4803 4864
rect 11570 4928 11886 4929
rect 11570 4864 11576 4928
rect 11640 4864 11656 4928
rect 11720 4864 11736 4928
rect 11800 4864 11816 4928
rect 11880 4864 11886 4928
rect 11570 4863 11886 4864
rect 18653 4928 18969 4929
rect 18653 4864 18659 4928
rect 18723 4864 18739 4928
rect 18803 4864 18819 4928
rect 18883 4864 18899 4928
rect 18963 4864 18969 4928
rect 18653 4863 18969 4864
rect 25736 4928 26052 4929
rect 25736 4864 25742 4928
rect 25806 4864 25822 4928
rect 25886 4864 25902 4928
rect 25966 4864 25982 4928
rect 26046 4864 26052 4928
rect 25736 4863 26052 4864
rect 8028 4384 8344 4385
rect 8028 4320 8034 4384
rect 8098 4320 8114 4384
rect 8178 4320 8194 4384
rect 8258 4320 8274 4384
rect 8338 4320 8344 4384
rect 8028 4319 8344 4320
rect 15111 4384 15427 4385
rect 15111 4320 15117 4384
rect 15181 4320 15197 4384
rect 15261 4320 15277 4384
rect 15341 4320 15357 4384
rect 15421 4320 15427 4384
rect 15111 4319 15427 4320
rect 22194 4384 22510 4385
rect 22194 4320 22200 4384
rect 22264 4320 22280 4384
rect 22344 4320 22360 4384
rect 22424 4320 22440 4384
rect 22504 4320 22510 4384
rect 22194 4319 22510 4320
rect 29277 4384 29593 4385
rect 29277 4320 29283 4384
rect 29347 4320 29363 4384
rect 29427 4320 29443 4384
rect 29507 4320 29523 4384
rect 29587 4320 29593 4384
rect 29277 4319 29593 4320
rect 2405 4042 2471 4045
rect 24209 4042 24275 4045
rect 2405 4040 24275 4042
rect 2405 3984 2410 4040
rect 2466 3984 24214 4040
rect 24270 3984 24275 4040
rect 2405 3982 24275 3984
rect 2405 3979 2471 3982
rect 24209 3979 24275 3982
rect 4487 3840 4803 3841
rect 4487 3776 4493 3840
rect 4557 3776 4573 3840
rect 4637 3776 4653 3840
rect 4717 3776 4733 3840
rect 4797 3776 4803 3840
rect 4487 3775 4803 3776
rect 11570 3840 11886 3841
rect 11570 3776 11576 3840
rect 11640 3776 11656 3840
rect 11720 3776 11736 3840
rect 11800 3776 11816 3840
rect 11880 3776 11886 3840
rect 11570 3775 11886 3776
rect 18653 3840 18969 3841
rect 18653 3776 18659 3840
rect 18723 3776 18739 3840
rect 18803 3776 18819 3840
rect 18883 3776 18899 3840
rect 18963 3776 18969 3840
rect 18653 3775 18969 3776
rect 25736 3840 26052 3841
rect 25736 3776 25742 3840
rect 25806 3776 25822 3840
rect 25886 3776 25902 3840
rect 25966 3776 25982 3840
rect 26046 3776 26052 3840
rect 25736 3775 26052 3776
rect 0 3498 800 3528
rect 933 3498 999 3501
rect 0 3496 999 3498
rect 0 3440 938 3496
rect 994 3440 999 3496
rect 0 3438 999 3440
rect 0 3408 800 3438
rect 933 3435 999 3438
rect 13169 3498 13235 3501
rect 15193 3498 15259 3501
rect 13169 3496 15259 3498
rect 13169 3440 13174 3496
rect 13230 3440 15198 3496
rect 15254 3440 15259 3496
rect 13169 3438 15259 3440
rect 13169 3435 13235 3438
rect 15193 3435 15259 3438
rect 8028 3296 8344 3297
rect 8028 3232 8034 3296
rect 8098 3232 8114 3296
rect 8178 3232 8194 3296
rect 8258 3232 8274 3296
rect 8338 3232 8344 3296
rect 8028 3231 8344 3232
rect 15111 3296 15427 3297
rect 15111 3232 15117 3296
rect 15181 3232 15197 3296
rect 15261 3232 15277 3296
rect 15341 3232 15357 3296
rect 15421 3232 15427 3296
rect 15111 3231 15427 3232
rect 22194 3296 22510 3297
rect 22194 3232 22200 3296
rect 22264 3232 22280 3296
rect 22344 3232 22360 3296
rect 22424 3232 22440 3296
rect 22504 3232 22510 3296
rect 22194 3231 22510 3232
rect 29277 3296 29593 3297
rect 29277 3232 29283 3296
rect 29347 3232 29363 3296
rect 29427 3232 29443 3296
rect 29507 3232 29523 3296
rect 29587 3232 29593 3296
rect 29277 3231 29593 3232
rect 28993 2818 29059 2821
rect 29781 2818 30581 2848
rect 28993 2816 30581 2818
rect 28993 2760 28998 2816
rect 29054 2760 30581 2816
rect 28993 2758 30581 2760
rect 28993 2755 29059 2758
rect 4487 2752 4803 2753
rect 4487 2688 4493 2752
rect 4557 2688 4573 2752
rect 4637 2688 4653 2752
rect 4717 2688 4733 2752
rect 4797 2688 4803 2752
rect 4487 2687 4803 2688
rect 11570 2752 11886 2753
rect 11570 2688 11576 2752
rect 11640 2688 11656 2752
rect 11720 2688 11736 2752
rect 11800 2688 11816 2752
rect 11880 2688 11886 2752
rect 11570 2687 11886 2688
rect 18653 2752 18969 2753
rect 18653 2688 18659 2752
rect 18723 2688 18739 2752
rect 18803 2688 18819 2752
rect 18883 2688 18899 2752
rect 18963 2688 18969 2752
rect 18653 2687 18969 2688
rect 25736 2752 26052 2753
rect 25736 2688 25742 2752
rect 25806 2688 25822 2752
rect 25886 2688 25902 2752
rect 25966 2688 25982 2752
rect 26046 2688 26052 2752
rect 29781 2728 30581 2758
rect 25736 2687 26052 2688
rect 8028 2208 8344 2209
rect 8028 2144 8034 2208
rect 8098 2144 8114 2208
rect 8178 2144 8194 2208
rect 8258 2144 8274 2208
rect 8338 2144 8344 2208
rect 8028 2143 8344 2144
rect 15111 2208 15427 2209
rect 15111 2144 15117 2208
rect 15181 2144 15197 2208
rect 15261 2144 15277 2208
rect 15341 2144 15357 2208
rect 15421 2144 15427 2208
rect 15111 2143 15427 2144
rect 22194 2208 22510 2209
rect 22194 2144 22200 2208
rect 22264 2144 22280 2208
rect 22344 2144 22360 2208
rect 22424 2144 22440 2208
rect 22504 2144 22510 2208
rect 22194 2143 22510 2144
rect 29277 2208 29593 2209
rect 29277 2144 29283 2208
rect 29347 2144 29363 2208
rect 29427 2144 29443 2208
rect 29507 2144 29523 2208
rect 29587 2144 29593 2208
rect 29277 2143 29593 2144
<< via3 >>
rect 8034 30492 8098 30496
rect 8034 30436 8038 30492
rect 8038 30436 8094 30492
rect 8094 30436 8098 30492
rect 8034 30432 8098 30436
rect 8114 30492 8178 30496
rect 8114 30436 8118 30492
rect 8118 30436 8174 30492
rect 8174 30436 8178 30492
rect 8114 30432 8178 30436
rect 8194 30492 8258 30496
rect 8194 30436 8198 30492
rect 8198 30436 8254 30492
rect 8254 30436 8258 30492
rect 8194 30432 8258 30436
rect 8274 30492 8338 30496
rect 8274 30436 8278 30492
rect 8278 30436 8334 30492
rect 8334 30436 8338 30492
rect 8274 30432 8338 30436
rect 15117 30492 15181 30496
rect 15117 30436 15121 30492
rect 15121 30436 15177 30492
rect 15177 30436 15181 30492
rect 15117 30432 15181 30436
rect 15197 30492 15261 30496
rect 15197 30436 15201 30492
rect 15201 30436 15257 30492
rect 15257 30436 15261 30492
rect 15197 30432 15261 30436
rect 15277 30492 15341 30496
rect 15277 30436 15281 30492
rect 15281 30436 15337 30492
rect 15337 30436 15341 30492
rect 15277 30432 15341 30436
rect 15357 30492 15421 30496
rect 15357 30436 15361 30492
rect 15361 30436 15417 30492
rect 15417 30436 15421 30492
rect 15357 30432 15421 30436
rect 22200 30492 22264 30496
rect 22200 30436 22204 30492
rect 22204 30436 22260 30492
rect 22260 30436 22264 30492
rect 22200 30432 22264 30436
rect 22280 30492 22344 30496
rect 22280 30436 22284 30492
rect 22284 30436 22340 30492
rect 22340 30436 22344 30492
rect 22280 30432 22344 30436
rect 22360 30492 22424 30496
rect 22360 30436 22364 30492
rect 22364 30436 22420 30492
rect 22420 30436 22424 30492
rect 22360 30432 22424 30436
rect 22440 30492 22504 30496
rect 22440 30436 22444 30492
rect 22444 30436 22500 30492
rect 22500 30436 22504 30492
rect 22440 30432 22504 30436
rect 29283 30492 29347 30496
rect 29283 30436 29287 30492
rect 29287 30436 29343 30492
rect 29343 30436 29347 30492
rect 29283 30432 29347 30436
rect 29363 30492 29427 30496
rect 29363 30436 29367 30492
rect 29367 30436 29423 30492
rect 29423 30436 29427 30492
rect 29363 30432 29427 30436
rect 29443 30492 29507 30496
rect 29443 30436 29447 30492
rect 29447 30436 29503 30492
rect 29503 30436 29507 30492
rect 29443 30432 29507 30436
rect 29523 30492 29587 30496
rect 29523 30436 29527 30492
rect 29527 30436 29583 30492
rect 29583 30436 29587 30492
rect 29523 30432 29587 30436
rect 4493 29948 4557 29952
rect 4493 29892 4497 29948
rect 4497 29892 4553 29948
rect 4553 29892 4557 29948
rect 4493 29888 4557 29892
rect 4573 29948 4637 29952
rect 4573 29892 4577 29948
rect 4577 29892 4633 29948
rect 4633 29892 4637 29948
rect 4573 29888 4637 29892
rect 4653 29948 4717 29952
rect 4653 29892 4657 29948
rect 4657 29892 4713 29948
rect 4713 29892 4717 29948
rect 4653 29888 4717 29892
rect 4733 29948 4797 29952
rect 4733 29892 4737 29948
rect 4737 29892 4793 29948
rect 4793 29892 4797 29948
rect 4733 29888 4797 29892
rect 11576 29948 11640 29952
rect 11576 29892 11580 29948
rect 11580 29892 11636 29948
rect 11636 29892 11640 29948
rect 11576 29888 11640 29892
rect 11656 29948 11720 29952
rect 11656 29892 11660 29948
rect 11660 29892 11716 29948
rect 11716 29892 11720 29948
rect 11656 29888 11720 29892
rect 11736 29948 11800 29952
rect 11736 29892 11740 29948
rect 11740 29892 11796 29948
rect 11796 29892 11800 29948
rect 11736 29888 11800 29892
rect 11816 29948 11880 29952
rect 11816 29892 11820 29948
rect 11820 29892 11876 29948
rect 11876 29892 11880 29948
rect 11816 29888 11880 29892
rect 18659 29948 18723 29952
rect 18659 29892 18663 29948
rect 18663 29892 18719 29948
rect 18719 29892 18723 29948
rect 18659 29888 18723 29892
rect 18739 29948 18803 29952
rect 18739 29892 18743 29948
rect 18743 29892 18799 29948
rect 18799 29892 18803 29948
rect 18739 29888 18803 29892
rect 18819 29948 18883 29952
rect 18819 29892 18823 29948
rect 18823 29892 18879 29948
rect 18879 29892 18883 29948
rect 18819 29888 18883 29892
rect 18899 29948 18963 29952
rect 18899 29892 18903 29948
rect 18903 29892 18959 29948
rect 18959 29892 18963 29948
rect 18899 29888 18963 29892
rect 25742 29948 25806 29952
rect 25742 29892 25746 29948
rect 25746 29892 25802 29948
rect 25802 29892 25806 29948
rect 25742 29888 25806 29892
rect 25822 29948 25886 29952
rect 25822 29892 25826 29948
rect 25826 29892 25882 29948
rect 25882 29892 25886 29948
rect 25822 29888 25886 29892
rect 25902 29948 25966 29952
rect 25902 29892 25906 29948
rect 25906 29892 25962 29948
rect 25962 29892 25966 29948
rect 25902 29888 25966 29892
rect 25982 29948 26046 29952
rect 25982 29892 25986 29948
rect 25986 29892 26042 29948
rect 26042 29892 26046 29948
rect 25982 29888 26046 29892
rect 8034 29404 8098 29408
rect 8034 29348 8038 29404
rect 8038 29348 8094 29404
rect 8094 29348 8098 29404
rect 8034 29344 8098 29348
rect 8114 29404 8178 29408
rect 8114 29348 8118 29404
rect 8118 29348 8174 29404
rect 8174 29348 8178 29404
rect 8114 29344 8178 29348
rect 8194 29404 8258 29408
rect 8194 29348 8198 29404
rect 8198 29348 8254 29404
rect 8254 29348 8258 29404
rect 8194 29344 8258 29348
rect 8274 29404 8338 29408
rect 8274 29348 8278 29404
rect 8278 29348 8334 29404
rect 8334 29348 8338 29404
rect 8274 29344 8338 29348
rect 15117 29404 15181 29408
rect 15117 29348 15121 29404
rect 15121 29348 15177 29404
rect 15177 29348 15181 29404
rect 15117 29344 15181 29348
rect 15197 29404 15261 29408
rect 15197 29348 15201 29404
rect 15201 29348 15257 29404
rect 15257 29348 15261 29404
rect 15197 29344 15261 29348
rect 15277 29404 15341 29408
rect 15277 29348 15281 29404
rect 15281 29348 15337 29404
rect 15337 29348 15341 29404
rect 15277 29344 15341 29348
rect 15357 29404 15421 29408
rect 15357 29348 15361 29404
rect 15361 29348 15417 29404
rect 15417 29348 15421 29404
rect 15357 29344 15421 29348
rect 22200 29404 22264 29408
rect 22200 29348 22204 29404
rect 22204 29348 22260 29404
rect 22260 29348 22264 29404
rect 22200 29344 22264 29348
rect 22280 29404 22344 29408
rect 22280 29348 22284 29404
rect 22284 29348 22340 29404
rect 22340 29348 22344 29404
rect 22280 29344 22344 29348
rect 22360 29404 22424 29408
rect 22360 29348 22364 29404
rect 22364 29348 22420 29404
rect 22420 29348 22424 29404
rect 22360 29344 22424 29348
rect 22440 29404 22504 29408
rect 22440 29348 22444 29404
rect 22444 29348 22500 29404
rect 22500 29348 22504 29404
rect 22440 29344 22504 29348
rect 29283 29404 29347 29408
rect 29283 29348 29287 29404
rect 29287 29348 29343 29404
rect 29343 29348 29347 29404
rect 29283 29344 29347 29348
rect 29363 29404 29427 29408
rect 29363 29348 29367 29404
rect 29367 29348 29423 29404
rect 29423 29348 29427 29404
rect 29363 29344 29427 29348
rect 29443 29404 29507 29408
rect 29443 29348 29447 29404
rect 29447 29348 29503 29404
rect 29503 29348 29507 29404
rect 29443 29344 29507 29348
rect 29523 29404 29587 29408
rect 29523 29348 29527 29404
rect 29527 29348 29583 29404
rect 29583 29348 29587 29404
rect 29523 29344 29587 29348
rect 28764 29064 28828 29068
rect 28764 29008 28778 29064
rect 28778 29008 28828 29064
rect 28764 29004 28828 29008
rect 4493 28860 4557 28864
rect 4493 28804 4497 28860
rect 4497 28804 4553 28860
rect 4553 28804 4557 28860
rect 4493 28800 4557 28804
rect 4573 28860 4637 28864
rect 4573 28804 4577 28860
rect 4577 28804 4633 28860
rect 4633 28804 4637 28860
rect 4573 28800 4637 28804
rect 4653 28860 4717 28864
rect 4653 28804 4657 28860
rect 4657 28804 4713 28860
rect 4713 28804 4717 28860
rect 4653 28800 4717 28804
rect 4733 28860 4797 28864
rect 4733 28804 4737 28860
rect 4737 28804 4793 28860
rect 4793 28804 4797 28860
rect 4733 28800 4797 28804
rect 11576 28860 11640 28864
rect 11576 28804 11580 28860
rect 11580 28804 11636 28860
rect 11636 28804 11640 28860
rect 11576 28800 11640 28804
rect 11656 28860 11720 28864
rect 11656 28804 11660 28860
rect 11660 28804 11716 28860
rect 11716 28804 11720 28860
rect 11656 28800 11720 28804
rect 11736 28860 11800 28864
rect 11736 28804 11740 28860
rect 11740 28804 11796 28860
rect 11796 28804 11800 28860
rect 11736 28800 11800 28804
rect 11816 28860 11880 28864
rect 11816 28804 11820 28860
rect 11820 28804 11876 28860
rect 11876 28804 11880 28860
rect 11816 28800 11880 28804
rect 18659 28860 18723 28864
rect 18659 28804 18663 28860
rect 18663 28804 18719 28860
rect 18719 28804 18723 28860
rect 18659 28800 18723 28804
rect 18739 28860 18803 28864
rect 18739 28804 18743 28860
rect 18743 28804 18799 28860
rect 18799 28804 18803 28860
rect 18739 28800 18803 28804
rect 18819 28860 18883 28864
rect 18819 28804 18823 28860
rect 18823 28804 18879 28860
rect 18879 28804 18883 28860
rect 18819 28800 18883 28804
rect 18899 28860 18963 28864
rect 18899 28804 18903 28860
rect 18903 28804 18959 28860
rect 18959 28804 18963 28860
rect 18899 28800 18963 28804
rect 25742 28860 25806 28864
rect 25742 28804 25746 28860
rect 25746 28804 25802 28860
rect 25802 28804 25806 28860
rect 25742 28800 25806 28804
rect 25822 28860 25886 28864
rect 25822 28804 25826 28860
rect 25826 28804 25882 28860
rect 25882 28804 25886 28860
rect 25822 28800 25886 28804
rect 25902 28860 25966 28864
rect 25902 28804 25906 28860
rect 25906 28804 25962 28860
rect 25962 28804 25966 28860
rect 25902 28800 25966 28804
rect 25982 28860 26046 28864
rect 25982 28804 25986 28860
rect 25986 28804 26042 28860
rect 26042 28804 26046 28860
rect 25982 28800 26046 28804
rect 8034 28316 8098 28320
rect 8034 28260 8038 28316
rect 8038 28260 8094 28316
rect 8094 28260 8098 28316
rect 8034 28256 8098 28260
rect 8114 28316 8178 28320
rect 8114 28260 8118 28316
rect 8118 28260 8174 28316
rect 8174 28260 8178 28316
rect 8114 28256 8178 28260
rect 8194 28316 8258 28320
rect 8194 28260 8198 28316
rect 8198 28260 8254 28316
rect 8254 28260 8258 28316
rect 8194 28256 8258 28260
rect 8274 28316 8338 28320
rect 8274 28260 8278 28316
rect 8278 28260 8334 28316
rect 8334 28260 8338 28316
rect 8274 28256 8338 28260
rect 15117 28316 15181 28320
rect 15117 28260 15121 28316
rect 15121 28260 15177 28316
rect 15177 28260 15181 28316
rect 15117 28256 15181 28260
rect 15197 28316 15261 28320
rect 15197 28260 15201 28316
rect 15201 28260 15257 28316
rect 15257 28260 15261 28316
rect 15197 28256 15261 28260
rect 15277 28316 15341 28320
rect 15277 28260 15281 28316
rect 15281 28260 15337 28316
rect 15337 28260 15341 28316
rect 15277 28256 15341 28260
rect 15357 28316 15421 28320
rect 15357 28260 15361 28316
rect 15361 28260 15417 28316
rect 15417 28260 15421 28316
rect 15357 28256 15421 28260
rect 22200 28316 22264 28320
rect 22200 28260 22204 28316
rect 22204 28260 22260 28316
rect 22260 28260 22264 28316
rect 22200 28256 22264 28260
rect 22280 28316 22344 28320
rect 22280 28260 22284 28316
rect 22284 28260 22340 28316
rect 22340 28260 22344 28316
rect 22280 28256 22344 28260
rect 22360 28316 22424 28320
rect 22360 28260 22364 28316
rect 22364 28260 22420 28316
rect 22420 28260 22424 28316
rect 22360 28256 22424 28260
rect 22440 28316 22504 28320
rect 22440 28260 22444 28316
rect 22444 28260 22500 28316
rect 22500 28260 22504 28316
rect 22440 28256 22504 28260
rect 29283 28316 29347 28320
rect 29283 28260 29287 28316
rect 29287 28260 29343 28316
rect 29343 28260 29347 28316
rect 29283 28256 29347 28260
rect 29363 28316 29427 28320
rect 29363 28260 29367 28316
rect 29367 28260 29423 28316
rect 29423 28260 29427 28316
rect 29363 28256 29427 28260
rect 29443 28316 29507 28320
rect 29443 28260 29447 28316
rect 29447 28260 29503 28316
rect 29503 28260 29507 28316
rect 29443 28256 29507 28260
rect 29523 28316 29587 28320
rect 29523 28260 29527 28316
rect 29527 28260 29583 28316
rect 29583 28260 29587 28316
rect 29523 28256 29587 28260
rect 4493 27772 4557 27776
rect 4493 27716 4497 27772
rect 4497 27716 4553 27772
rect 4553 27716 4557 27772
rect 4493 27712 4557 27716
rect 4573 27772 4637 27776
rect 4573 27716 4577 27772
rect 4577 27716 4633 27772
rect 4633 27716 4637 27772
rect 4573 27712 4637 27716
rect 4653 27772 4717 27776
rect 4653 27716 4657 27772
rect 4657 27716 4713 27772
rect 4713 27716 4717 27772
rect 4653 27712 4717 27716
rect 4733 27772 4797 27776
rect 4733 27716 4737 27772
rect 4737 27716 4793 27772
rect 4793 27716 4797 27772
rect 4733 27712 4797 27716
rect 11576 27772 11640 27776
rect 11576 27716 11580 27772
rect 11580 27716 11636 27772
rect 11636 27716 11640 27772
rect 11576 27712 11640 27716
rect 11656 27772 11720 27776
rect 11656 27716 11660 27772
rect 11660 27716 11716 27772
rect 11716 27716 11720 27772
rect 11656 27712 11720 27716
rect 11736 27772 11800 27776
rect 11736 27716 11740 27772
rect 11740 27716 11796 27772
rect 11796 27716 11800 27772
rect 11736 27712 11800 27716
rect 11816 27772 11880 27776
rect 11816 27716 11820 27772
rect 11820 27716 11876 27772
rect 11876 27716 11880 27772
rect 11816 27712 11880 27716
rect 18659 27772 18723 27776
rect 18659 27716 18663 27772
rect 18663 27716 18719 27772
rect 18719 27716 18723 27772
rect 18659 27712 18723 27716
rect 18739 27772 18803 27776
rect 18739 27716 18743 27772
rect 18743 27716 18799 27772
rect 18799 27716 18803 27772
rect 18739 27712 18803 27716
rect 18819 27772 18883 27776
rect 18819 27716 18823 27772
rect 18823 27716 18879 27772
rect 18879 27716 18883 27772
rect 18819 27712 18883 27716
rect 18899 27772 18963 27776
rect 18899 27716 18903 27772
rect 18903 27716 18959 27772
rect 18959 27716 18963 27772
rect 18899 27712 18963 27716
rect 25742 27772 25806 27776
rect 25742 27716 25746 27772
rect 25746 27716 25802 27772
rect 25802 27716 25806 27772
rect 25742 27712 25806 27716
rect 25822 27772 25886 27776
rect 25822 27716 25826 27772
rect 25826 27716 25882 27772
rect 25882 27716 25886 27772
rect 25822 27712 25886 27716
rect 25902 27772 25966 27776
rect 25902 27716 25906 27772
rect 25906 27716 25962 27772
rect 25962 27716 25966 27772
rect 25902 27712 25966 27716
rect 25982 27772 26046 27776
rect 25982 27716 25986 27772
rect 25986 27716 26042 27772
rect 26042 27716 26046 27772
rect 25982 27712 26046 27716
rect 8034 27228 8098 27232
rect 8034 27172 8038 27228
rect 8038 27172 8094 27228
rect 8094 27172 8098 27228
rect 8034 27168 8098 27172
rect 8114 27228 8178 27232
rect 8114 27172 8118 27228
rect 8118 27172 8174 27228
rect 8174 27172 8178 27228
rect 8114 27168 8178 27172
rect 8194 27228 8258 27232
rect 8194 27172 8198 27228
rect 8198 27172 8254 27228
rect 8254 27172 8258 27228
rect 8194 27168 8258 27172
rect 8274 27228 8338 27232
rect 8274 27172 8278 27228
rect 8278 27172 8334 27228
rect 8334 27172 8338 27228
rect 8274 27168 8338 27172
rect 15117 27228 15181 27232
rect 15117 27172 15121 27228
rect 15121 27172 15177 27228
rect 15177 27172 15181 27228
rect 15117 27168 15181 27172
rect 15197 27228 15261 27232
rect 15197 27172 15201 27228
rect 15201 27172 15257 27228
rect 15257 27172 15261 27228
rect 15197 27168 15261 27172
rect 15277 27228 15341 27232
rect 15277 27172 15281 27228
rect 15281 27172 15337 27228
rect 15337 27172 15341 27228
rect 15277 27168 15341 27172
rect 15357 27228 15421 27232
rect 15357 27172 15361 27228
rect 15361 27172 15417 27228
rect 15417 27172 15421 27228
rect 15357 27168 15421 27172
rect 22200 27228 22264 27232
rect 22200 27172 22204 27228
rect 22204 27172 22260 27228
rect 22260 27172 22264 27228
rect 22200 27168 22264 27172
rect 22280 27228 22344 27232
rect 22280 27172 22284 27228
rect 22284 27172 22340 27228
rect 22340 27172 22344 27228
rect 22280 27168 22344 27172
rect 22360 27228 22424 27232
rect 22360 27172 22364 27228
rect 22364 27172 22420 27228
rect 22420 27172 22424 27228
rect 22360 27168 22424 27172
rect 22440 27228 22504 27232
rect 22440 27172 22444 27228
rect 22444 27172 22500 27228
rect 22500 27172 22504 27228
rect 22440 27168 22504 27172
rect 29283 27228 29347 27232
rect 29283 27172 29287 27228
rect 29287 27172 29343 27228
rect 29343 27172 29347 27228
rect 29283 27168 29347 27172
rect 29363 27228 29427 27232
rect 29363 27172 29367 27228
rect 29367 27172 29423 27228
rect 29423 27172 29427 27228
rect 29363 27168 29427 27172
rect 29443 27228 29507 27232
rect 29443 27172 29447 27228
rect 29447 27172 29503 27228
rect 29503 27172 29507 27228
rect 29443 27168 29507 27172
rect 29523 27228 29587 27232
rect 29523 27172 29527 27228
rect 29527 27172 29583 27228
rect 29583 27172 29587 27228
rect 29523 27168 29587 27172
rect 4493 26684 4557 26688
rect 4493 26628 4497 26684
rect 4497 26628 4553 26684
rect 4553 26628 4557 26684
rect 4493 26624 4557 26628
rect 4573 26684 4637 26688
rect 4573 26628 4577 26684
rect 4577 26628 4633 26684
rect 4633 26628 4637 26684
rect 4573 26624 4637 26628
rect 4653 26684 4717 26688
rect 4653 26628 4657 26684
rect 4657 26628 4713 26684
rect 4713 26628 4717 26684
rect 4653 26624 4717 26628
rect 4733 26684 4797 26688
rect 4733 26628 4737 26684
rect 4737 26628 4793 26684
rect 4793 26628 4797 26684
rect 4733 26624 4797 26628
rect 11576 26684 11640 26688
rect 11576 26628 11580 26684
rect 11580 26628 11636 26684
rect 11636 26628 11640 26684
rect 11576 26624 11640 26628
rect 11656 26684 11720 26688
rect 11656 26628 11660 26684
rect 11660 26628 11716 26684
rect 11716 26628 11720 26684
rect 11656 26624 11720 26628
rect 11736 26684 11800 26688
rect 11736 26628 11740 26684
rect 11740 26628 11796 26684
rect 11796 26628 11800 26684
rect 11736 26624 11800 26628
rect 11816 26684 11880 26688
rect 11816 26628 11820 26684
rect 11820 26628 11876 26684
rect 11876 26628 11880 26684
rect 11816 26624 11880 26628
rect 18659 26684 18723 26688
rect 18659 26628 18663 26684
rect 18663 26628 18719 26684
rect 18719 26628 18723 26684
rect 18659 26624 18723 26628
rect 18739 26684 18803 26688
rect 18739 26628 18743 26684
rect 18743 26628 18799 26684
rect 18799 26628 18803 26684
rect 18739 26624 18803 26628
rect 18819 26684 18883 26688
rect 18819 26628 18823 26684
rect 18823 26628 18879 26684
rect 18879 26628 18883 26684
rect 18819 26624 18883 26628
rect 18899 26684 18963 26688
rect 18899 26628 18903 26684
rect 18903 26628 18959 26684
rect 18959 26628 18963 26684
rect 18899 26624 18963 26628
rect 25742 26684 25806 26688
rect 25742 26628 25746 26684
rect 25746 26628 25802 26684
rect 25802 26628 25806 26684
rect 25742 26624 25806 26628
rect 25822 26684 25886 26688
rect 25822 26628 25826 26684
rect 25826 26628 25882 26684
rect 25882 26628 25886 26684
rect 25822 26624 25886 26628
rect 25902 26684 25966 26688
rect 25902 26628 25906 26684
rect 25906 26628 25962 26684
rect 25962 26628 25966 26684
rect 25902 26624 25966 26628
rect 25982 26684 26046 26688
rect 25982 26628 25986 26684
rect 25986 26628 26042 26684
rect 26042 26628 26046 26684
rect 25982 26624 26046 26628
rect 8034 26140 8098 26144
rect 8034 26084 8038 26140
rect 8038 26084 8094 26140
rect 8094 26084 8098 26140
rect 8034 26080 8098 26084
rect 8114 26140 8178 26144
rect 8114 26084 8118 26140
rect 8118 26084 8174 26140
rect 8174 26084 8178 26140
rect 8114 26080 8178 26084
rect 8194 26140 8258 26144
rect 8194 26084 8198 26140
rect 8198 26084 8254 26140
rect 8254 26084 8258 26140
rect 8194 26080 8258 26084
rect 8274 26140 8338 26144
rect 8274 26084 8278 26140
rect 8278 26084 8334 26140
rect 8334 26084 8338 26140
rect 8274 26080 8338 26084
rect 15117 26140 15181 26144
rect 15117 26084 15121 26140
rect 15121 26084 15177 26140
rect 15177 26084 15181 26140
rect 15117 26080 15181 26084
rect 15197 26140 15261 26144
rect 15197 26084 15201 26140
rect 15201 26084 15257 26140
rect 15257 26084 15261 26140
rect 15197 26080 15261 26084
rect 15277 26140 15341 26144
rect 15277 26084 15281 26140
rect 15281 26084 15337 26140
rect 15337 26084 15341 26140
rect 15277 26080 15341 26084
rect 15357 26140 15421 26144
rect 15357 26084 15361 26140
rect 15361 26084 15417 26140
rect 15417 26084 15421 26140
rect 15357 26080 15421 26084
rect 22200 26140 22264 26144
rect 22200 26084 22204 26140
rect 22204 26084 22260 26140
rect 22260 26084 22264 26140
rect 22200 26080 22264 26084
rect 22280 26140 22344 26144
rect 22280 26084 22284 26140
rect 22284 26084 22340 26140
rect 22340 26084 22344 26140
rect 22280 26080 22344 26084
rect 22360 26140 22424 26144
rect 22360 26084 22364 26140
rect 22364 26084 22420 26140
rect 22420 26084 22424 26140
rect 22360 26080 22424 26084
rect 22440 26140 22504 26144
rect 22440 26084 22444 26140
rect 22444 26084 22500 26140
rect 22500 26084 22504 26140
rect 22440 26080 22504 26084
rect 29283 26140 29347 26144
rect 29283 26084 29287 26140
rect 29287 26084 29343 26140
rect 29343 26084 29347 26140
rect 29283 26080 29347 26084
rect 29363 26140 29427 26144
rect 29363 26084 29367 26140
rect 29367 26084 29423 26140
rect 29423 26084 29427 26140
rect 29363 26080 29427 26084
rect 29443 26140 29507 26144
rect 29443 26084 29447 26140
rect 29447 26084 29503 26140
rect 29503 26084 29507 26140
rect 29443 26080 29507 26084
rect 29523 26140 29587 26144
rect 29523 26084 29527 26140
rect 29527 26084 29583 26140
rect 29583 26084 29587 26140
rect 29523 26080 29587 26084
rect 4493 25596 4557 25600
rect 4493 25540 4497 25596
rect 4497 25540 4553 25596
rect 4553 25540 4557 25596
rect 4493 25536 4557 25540
rect 4573 25596 4637 25600
rect 4573 25540 4577 25596
rect 4577 25540 4633 25596
rect 4633 25540 4637 25596
rect 4573 25536 4637 25540
rect 4653 25596 4717 25600
rect 4653 25540 4657 25596
rect 4657 25540 4713 25596
rect 4713 25540 4717 25596
rect 4653 25536 4717 25540
rect 4733 25596 4797 25600
rect 4733 25540 4737 25596
rect 4737 25540 4793 25596
rect 4793 25540 4797 25596
rect 4733 25536 4797 25540
rect 11576 25596 11640 25600
rect 11576 25540 11580 25596
rect 11580 25540 11636 25596
rect 11636 25540 11640 25596
rect 11576 25536 11640 25540
rect 11656 25596 11720 25600
rect 11656 25540 11660 25596
rect 11660 25540 11716 25596
rect 11716 25540 11720 25596
rect 11656 25536 11720 25540
rect 11736 25596 11800 25600
rect 11736 25540 11740 25596
rect 11740 25540 11796 25596
rect 11796 25540 11800 25596
rect 11736 25536 11800 25540
rect 11816 25596 11880 25600
rect 11816 25540 11820 25596
rect 11820 25540 11876 25596
rect 11876 25540 11880 25596
rect 11816 25536 11880 25540
rect 18659 25596 18723 25600
rect 18659 25540 18663 25596
rect 18663 25540 18719 25596
rect 18719 25540 18723 25596
rect 18659 25536 18723 25540
rect 18739 25596 18803 25600
rect 18739 25540 18743 25596
rect 18743 25540 18799 25596
rect 18799 25540 18803 25596
rect 18739 25536 18803 25540
rect 18819 25596 18883 25600
rect 18819 25540 18823 25596
rect 18823 25540 18879 25596
rect 18879 25540 18883 25596
rect 18819 25536 18883 25540
rect 18899 25596 18963 25600
rect 18899 25540 18903 25596
rect 18903 25540 18959 25596
rect 18959 25540 18963 25596
rect 18899 25536 18963 25540
rect 25742 25596 25806 25600
rect 25742 25540 25746 25596
rect 25746 25540 25802 25596
rect 25802 25540 25806 25596
rect 25742 25536 25806 25540
rect 25822 25596 25886 25600
rect 25822 25540 25826 25596
rect 25826 25540 25882 25596
rect 25882 25540 25886 25596
rect 25822 25536 25886 25540
rect 25902 25596 25966 25600
rect 25902 25540 25906 25596
rect 25906 25540 25962 25596
rect 25962 25540 25966 25596
rect 25902 25536 25966 25540
rect 25982 25596 26046 25600
rect 25982 25540 25986 25596
rect 25986 25540 26042 25596
rect 26042 25540 26046 25596
rect 25982 25536 26046 25540
rect 8034 25052 8098 25056
rect 8034 24996 8038 25052
rect 8038 24996 8094 25052
rect 8094 24996 8098 25052
rect 8034 24992 8098 24996
rect 8114 25052 8178 25056
rect 8114 24996 8118 25052
rect 8118 24996 8174 25052
rect 8174 24996 8178 25052
rect 8114 24992 8178 24996
rect 8194 25052 8258 25056
rect 8194 24996 8198 25052
rect 8198 24996 8254 25052
rect 8254 24996 8258 25052
rect 8194 24992 8258 24996
rect 8274 25052 8338 25056
rect 8274 24996 8278 25052
rect 8278 24996 8334 25052
rect 8334 24996 8338 25052
rect 8274 24992 8338 24996
rect 15117 25052 15181 25056
rect 15117 24996 15121 25052
rect 15121 24996 15177 25052
rect 15177 24996 15181 25052
rect 15117 24992 15181 24996
rect 15197 25052 15261 25056
rect 15197 24996 15201 25052
rect 15201 24996 15257 25052
rect 15257 24996 15261 25052
rect 15197 24992 15261 24996
rect 15277 25052 15341 25056
rect 15277 24996 15281 25052
rect 15281 24996 15337 25052
rect 15337 24996 15341 25052
rect 15277 24992 15341 24996
rect 15357 25052 15421 25056
rect 15357 24996 15361 25052
rect 15361 24996 15417 25052
rect 15417 24996 15421 25052
rect 15357 24992 15421 24996
rect 22200 25052 22264 25056
rect 22200 24996 22204 25052
rect 22204 24996 22260 25052
rect 22260 24996 22264 25052
rect 22200 24992 22264 24996
rect 22280 25052 22344 25056
rect 22280 24996 22284 25052
rect 22284 24996 22340 25052
rect 22340 24996 22344 25052
rect 22280 24992 22344 24996
rect 22360 25052 22424 25056
rect 22360 24996 22364 25052
rect 22364 24996 22420 25052
rect 22420 24996 22424 25052
rect 22360 24992 22424 24996
rect 22440 25052 22504 25056
rect 22440 24996 22444 25052
rect 22444 24996 22500 25052
rect 22500 24996 22504 25052
rect 22440 24992 22504 24996
rect 29283 25052 29347 25056
rect 29283 24996 29287 25052
rect 29287 24996 29343 25052
rect 29343 24996 29347 25052
rect 29283 24992 29347 24996
rect 29363 25052 29427 25056
rect 29363 24996 29367 25052
rect 29367 24996 29423 25052
rect 29423 24996 29427 25052
rect 29363 24992 29427 24996
rect 29443 25052 29507 25056
rect 29443 24996 29447 25052
rect 29447 24996 29503 25052
rect 29503 24996 29507 25052
rect 29443 24992 29507 24996
rect 29523 25052 29587 25056
rect 29523 24996 29527 25052
rect 29527 24996 29583 25052
rect 29583 24996 29587 25052
rect 29523 24992 29587 24996
rect 4493 24508 4557 24512
rect 4493 24452 4497 24508
rect 4497 24452 4553 24508
rect 4553 24452 4557 24508
rect 4493 24448 4557 24452
rect 4573 24508 4637 24512
rect 4573 24452 4577 24508
rect 4577 24452 4633 24508
rect 4633 24452 4637 24508
rect 4573 24448 4637 24452
rect 4653 24508 4717 24512
rect 4653 24452 4657 24508
rect 4657 24452 4713 24508
rect 4713 24452 4717 24508
rect 4653 24448 4717 24452
rect 4733 24508 4797 24512
rect 4733 24452 4737 24508
rect 4737 24452 4793 24508
rect 4793 24452 4797 24508
rect 4733 24448 4797 24452
rect 11576 24508 11640 24512
rect 11576 24452 11580 24508
rect 11580 24452 11636 24508
rect 11636 24452 11640 24508
rect 11576 24448 11640 24452
rect 11656 24508 11720 24512
rect 11656 24452 11660 24508
rect 11660 24452 11716 24508
rect 11716 24452 11720 24508
rect 11656 24448 11720 24452
rect 11736 24508 11800 24512
rect 11736 24452 11740 24508
rect 11740 24452 11796 24508
rect 11796 24452 11800 24508
rect 11736 24448 11800 24452
rect 11816 24508 11880 24512
rect 11816 24452 11820 24508
rect 11820 24452 11876 24508
rect 11876 24452 11880 24508
rect 11816 24448 11880 24452
rect 18659 24508 18723 24512
rect 18659 24452 18663 24508
rect 18663 24452 18719 24508
rect 18719 24452 18723 24508
rect 18659 24448 18723 24452
rect 18739 24508 18803 24512
rect 18739 24452 18743 24508
rect 18743 24452 18799 24508
rect 18799 24452 18803 24508
rect 18739 24448 18803 24452
rect 18819 24508 18883 24512
rect 18819 24452 18823 24508
rect 18823 24452 18879 24508
rect 18879 24452 18883 24508
rect 18819 24448 18883 24452
rect 18899 24508 18963 24512
rect 18899 24452 18903 24508
rect 18903 24452 18959 24508
rect 18959 24452 18963 24508
rect 18899 24448 18963 24452
rect 25742 24508 25806 24512
rect 25742 24452 25746 24508
rect 25746 24452 25802 24508
rect 25802 24452 25806 24508
rect 25742 24448 25806 24452
rect 25822 24508 25886 24512
rect 25822 24452 25826 24508
rect 25826 24452 25882 24508
rect 25882 24452 25886 24508
rect 25822 24448 25886 24452
rect 25902 24508 25966 24512
rect 25902 24452 25906 24508
rect 25906 24452 25962 24508
rect 25962 24452 25966 24508
rect 25902 24448 25966 24452
rect 25982 24508 26046 24512
rect 25982 24452 25986 24508
rect 25986 24452 26042 24508
rect 26042 24452 26046 24508
rect 25982 24448 26046 24452
rect 8034 23964 8098 23968
rect 8034 23908 8038 23964
rect 8038 23908 8094 23964
rect 8094 23908 8098 23964
rect 8034 23904 8098 23908
rect 8114 23964 8178 23968
rect 8114 23908 8118 23964
rect 8118 23908 8174 23964
rect 8174 23908 8178 23964
rect 8114 23904 8178 23908
rect 8194 23964 8258 23968
rect 8194 23908 8198 23964
rect 8198 23908 8254 23964
rect 8254 23908 8258 23964
rect 8194 23904 8258 23908
rect 8274 23964 8338 23968
rect 8274 23908 8278 23964
rect 8278 23908 8334 23964
rect 8334 23908 8338 23964
rect 8274 23904 8338 23908
rect 15117 23964 15181 23968
rect 15117 23908 15121 23964
rect 15121 23908 15177 23964
rect 15177 23908 15181 23964
rect 15117 23904 15181 23908
rect 15197 23964 15261 23968
rect 15197 23908 15201 23964
rect 15201 23908 15257 23964
rect 15257 23908 15261 23964
rect 15197 23904 15261 23908
rect 15277 23964 15341 23968
rect 15277 23908 15281 23964
rect 15281 23908 15337 23964
rect 15337 23908 15341 23964
rect 15277 23904 15341 23908
rect 15357 23964 15421 23968
rect 15357 23908 15361 23964
rect 15361 23908 15417 23964
rect 15417 23908 15421 23964
rect 15357 23904 15421 23908
rect 22200 23964 22264 23968
rect 22200 23908 22204 23964
rect 22204 23908 22260 23964
rect 22260 23908 22264 23964
rect 22200 23904 22264 23908
rect 22280 23964 22344 23968
rect 22280 23908 22284 23964
rect 22284 23908 22340 23964
rect 22340 23908 22344 23964
rect 22280 23904 22344 23908
rect 22360 23964 22424 23968
rect 22360 23908 22364 23964
rect 22364 23908 22420 23964
rect 22420 23908 22424 23964
rect 22360 23904 22424 23908
rect 22440 23964 22504 23968
rect 22440 23908 22444 23964
rect 22444 23908 22500 23964
rect 22500 23908 22504 23964
rect 22440 23904 22504 23908
rect 29283 23964 29347 23968
rect 29283 23908 29287 23964
rect 29287 23908 29343 23964
rect 29343 23908 29347 23964
rect 29283 23904 29347 23908
rect 29363 23964 29427 23968
rect 29363 23908 29367 23964
rect 29367 23908 29423 23964
rect 29423 23908 29427 23964
rect 29363 23904 29427 23908
rect 29443 23964 29507 23968
rect 29443 23908 29447 23964
rect 29447 23908 29503 23964
rect 29503 23908 29507 23964
rect 29443 23904 29507 23908
rect 29523 23964 29587 23968
rect 29523 23908 29527 23964
rect 29527 23908 29583 23964
rect 29583 23908 29587 23964
rect 29523 23904 29587 23908
rect 4493 23420 4557 23424
rect 4493 23364 4497 23420
rect 4497 23364 4553 23420
rect 4553 23364 4557 23420
rect 4493 23360 4557 23364
rect 4573 23420 4637 23424
rect 4573 23364 4577 23420
rect 4577 23364 4633 23420
rect 4633 23364 4637 23420
rect 4573 23360 4637 23364
rect 4653 23420 4717 23424
rect 4653 23364 4657 23420
rect 4657 23364 4713 23420
rect 4713 23364 4717 23420
rect 4653 23360 4717 23364
rect 4733 23420 4797 23424
rect 4733 23364 4737 23420
rect 4737 23364 4793 23420
rect 4793 23364 4797 23420
rect 4733 23360 4797 23364
rect 11576 23420 11640 23424
rect 11576 23364 11580 23420
rect 11580 23364 11636 23420
rect 11636 23364 11640 23420
rect 11576 23360 11640 23364
rect 11656 23420 11720 23424
rect 11656 23364 11660 23420
rect 11660 23364 11716 23420
rect 11716 23364 11720 23420
rect 11656 23360 11720 23364
rect 11736 23420 11800 23424
rect 11736 23364 11740 23420
rect 11740 23364 11796 23420
rect 11796 23364 11800 23420
rect 11736 23360 11800 23364
rect 11816 23420 11880 23424
rect 11816 23364 11820 23420
rect 11820 23364 11876 23420
rect 11876 23364 11880 23420
rect 11816 23360 11880 23364
rect 18659 23420 18723 23424
rect 18659 23364 18663 23420
rect 18663 23364 18719 23420
rect 18719 23364 18723 23420
rect 18659 23360 18723 23364
rect 18739 23420 18803 23424
rect 18739 23364 18743 23420
rect 18743 23364 18799 23420
rect 18799 23364 18803 23420
rect 18739 23360 18803 23364
rect 18819 23420 18883 23424
rect 18819 23364 18823 23420
rect 18823 23364 18879 23420
rect 18879 23364 18883 23420
rect 18819 23360 18883 23364
rect 18899 23420 18963 23424
rect 18899 23364 18903 23420
rect 18903 23364 18959 23420
rect 18959 23364 18963 23420
rect 18899 23360 18963 23364
rect 25742 23420 25806 23424
rect 25742 23364 25746 23420
rect 25746 23364 25802 23420
rect 25802 23364 25806 23420
rect 25742 23360 25806 23364
rect 25822 23420 25886 23424
rect 25822 23364 25826 23420
rect 25826 23364 25882 23420
rect 25882 23364 25886 23420
rect 25822 23360 25886 23364
rect 25902 23420 25966 23424
rect 25902 23364 25906 23420
rect 25906 23364 25962 23420
rect 25962 23364 25966 23420
rect 25902 23360 25966 23364
rect 25982 23420 26046 23424
rect 25982 23364 25986 23420
rect 25986 23364 26042 23420
rect 26042 23364 26046 23420
rect 25982 23360 26046 23364
rect 8034 22876 8098 22880
rect 8034 22820 8038 22876
rect 8038 22820 8094 22876
rect 8094 22820 8098 22876
rect 8034 22816 8098 22820
rect 8114 22876 8178 22880
rect 8114 22820 8118 22876
rect 8118 22820 8174 22876
rect 8174 22820 8178 22876
rect 8114 22816 8178 22820
rect 8194 22876 8258 22880
rect 8194 22820 8198 22876
rect 8198 22820 8254 22876
rect 8254 22820 8258 22876
rect 8194 22816 8258 22820
rect 8274 22876 8338 22880
rect 8274 22820 8278 22876
rect 8278 22820 8334 22876
rect 8334 22820 8338 22876
rect 8274 22816 8338 22820
rect 15117 22876 15181 22880
rect 15117 22820 15121 22876
rect 15121 22820 15177 22876
rect 15177 22820 15181 22876
rect 15117 22816 15181 22820
rect 15197 22876 15261 22880
rect 15197 22820 15201 22876
rect 15201 22820 15257 22876
rect 15257 22820 15261 22876
rect 15197 22816 15261 22820
rect 15277 22876 15341 22880
rect 15277 22820 15281 22876
rect 15281 22820 15337 22876
rect 15337 22820 15341 22876
rect 15277 22816 15341 22820
rect 15357 22876 15421 22880
rect 15357 22820 15361 22876
rect 15361 22820 15417 22876
rect 15417 22820 15421 22876
rect 15357 22816 15421 22820
rect 22200 22876 22264 22880
rect 22200 22820 22204 22876
rect 22204 22820 22260 22876
rect 22260 22820 22264 22876
rect 22200 22816 22264 22820
rect 22280 22876 22344 22880
rect 22280 22820 22284 22876
rect 22284 22820 22340 22876
rect 22340 22820 22344 22876
rect 22280 22816 22344 22820
rect 22360 22876 22424 22880
rect 22360 22820 22364 22876
rect 22364 22820 22420 22876
rect 22420 22820 22424 22876
rect 22360 22816 22424 22820
rect 22440 22876 22504 22880
rect 22440 22820 22444 22876
rect 22444 22820 22500 22876
rect 22500 22820 22504 22876
rect 22440 22816 22504 22820
rect 29283 22876 29347 22880
rect 29283 22820 29287 22876
rect 29287 22820 29343 22876
rect 29343 22820 29347 22876
rect 29283 22816 29347 22820
rect 29363 22876 29427 22880
rect 29363 22820 29367 22876
rect 29367 22820 29423 22876
rect 29423 22820 29427 22876
rect 29363 22816 29427 22820
rect 29443 22876 29507 22880
rect 29443 22820 29447 22876
rect 29447 22820 29503 22876
rect 29503 22820 29507 22876
rect 29443 22816 29507 22820
rect 29523 22876 29587 22880
rect 29523 22820 29527 22876
rect 29527 22820 29583 22876
rect 29583 22820 29587 22876
rect 29523 22816 29587 22820
rect 24348 22536 24412 22540
rect 24348 22480 24398 22536
rect 24398 22480 24412 22536
rect 24348 22476 24412 22480
rect 4493 22332 4557 22336
rect 4493 22276 4497 22332
rect 4497 22276 4553 22332
rect 4553 22276 4557 22332
rect 4493 22272 4557 22276
rect 4573 22332 4637 22336
rect 4573 22276 4577 22332
rect 4577 22276 4633 22332
rect 4633 22276 4637 22332
rect 4573 22272 4637 22276
rect 4653 22332 4717 22336
rect 4653 22276 4657 22332
rect 4657 22276 4713 22332
rect 4713 22276 4717 22332
rect 4653 22272 4717 22276
rect 4733 22332 4797 22336
rect 4733 22276 4737 22332
rect 4737 22276 4793 22332
rect 4793 22276 4797 22332
rect 4733 22272 4797 22276
rect 11576 22332 11640 22336
rect 11576 22276 11580 22332
rect 11580 22276 11636 22332
rect 11636 22276 11640 22332
rect 11576 22272 11640 22276
rect 11656 22332 11720 22336
rect 11656 22276 11660 22332
rect 11660 22276 11716 22332
rect 11716 22276 11720 22332
rect 11656 22272 11720 22276
rect 11736 22332 11800 22336
rect 11736 22276 11740 22332
rect 11740 22276 11796 22332
rect 11796 22276 11800 22332
rect 11736 22272 11800 22276
rect 11816 22332 11880 22336
rect 11816 22276 11820 22332
rect 11820 22276 11876 22332
rect 11876 22276 11880 22332
rect 11816 22272 11880 22276
rect 18659 22332 18723 22336
rect 18659 22276 18663 22332
rect 18663 22276 18719 22332
rect 18719 22276 18723 22332
rect 18659 22272 18723 22276
rect 18739 22332 18803 22336
rect 18739 22276 18743 22332
rect 18743 22276 18799 22332
rect 18799 22276 18803 22332
rect 18739 22272 18803 22276
rect 18819 22332 18883 22336
rect 18819 22276 18823 22332
rect 18823 22276 18879 22332
rect 18879 22276 18883 22332
rect 18819 22272 18883 22276
rect 18899 22332 18963 22336
rect 18899 22276 18903 22332
rect 18903 22276 18959 22332
rect 18959 22276 18963 22332
rect 18899 22272 18963 22276
rect 25742 22332 25806 22336
rect 25742 22276 25746 22332
rect 25746 22276 25802 22332
rect 25802 22276 25806 22332
rect 25742 22272 25806 22276
rect 25822 22332 25886 22336
rect 25822 22276 25826 22332
rect 25826 22276 25882 22332
rect 25882 22276 25886 22332
rect 25822 22272 25886 22276
rect 25902 22332 25966 22336
rect 25902 22276 25906 22332
rect 25906 22276 25962 22332
rect 25962 22276 25966 22332
rect 25902 22272 25966 22276
rect 25982 22332 26046 22336
rect 25982 22276 25986 22332
rect 25986 22276 26042 22332
rect 26042 22276 26046 22332
rect 25982 22272 26046 22276
rect 8034 21788 8098 21792
rect 8034 21732 8038 21788
rect 8038 21732 8094 21788
rect 8094 21732 8098 21788
rect 8034 21728 8098 21732
rect 8114 21788 8178 21792
rect 8114 21732 8118 21788
rect 8118 21732 8174 21788
rect 8174 21732 8178 21788
rect 8114 21728 8178 21732
rect 8194 21788 8258 21792
rect 8194 21732 8198 21788
rect 8198 21732 8254 21788
rect 8254 21732 8258 21788
rect 8194 21728 8258 21732
rect 8274 21788 8338 21792
rect 8274 21732 8278 21788
rect 8278 21732 8334 21788
rect 8334 21732 8338 21788
rect 8274 21728 8338 21732
rect 15117 21788 15181 21792
rect 15117 21732 15121 21788
rect 15121 21732 15177 21788
rect 15177 21732 15181 21788
rect 15117 21728 15181 21732
rect 15197 21788 15261 21792
rect 15197 21732 15201 21788
rect 15201 21732 15257 21788
rect 15257 21732 15261 21788
rect 15197 21728 15261 21732
rect 15277 21788 15341 21792
rect 15277 21732 15281 21788
rect 15281 21732 15337 21788
rect 15337 21732 15341 21788
rect 15277 21728 15341 21732
rect 15357 21788 15421 21792
rect 15357 21732 15361 21788
rect 15361 21732 15417 21788
rect 15417 21732 15421 21788
rect 15357 21728 15421 21732
rect 22200 21788 22264 21792
rect 22200 21732 22204 21788
rect 22204 21732 22260 21788
rect 22260 21732 22264 21788
rect 22200 21728 22264 21732
rect 22280 21788 22344 21792
rect 22280 21732 22284 21788
rect 22284 21732 22340 21788
rect 22340 21732 22344 21788
rect 22280 21728 22344 21732
rect 22360 21788 22424 21792
rect 22360 21732 22364 21788
rect 22364 21732 22420 21788
rect 22420 21732 22424 21788
rect 22360 21728 22424 21732
rect 22440 21788 22504 21792
rect 22440 21732 22444 21788
rect 22444 21732 22500 21788
rect 22500 21732 22504 21788
rect 22440 21728 22504 21732
rect 29283 21788 29347 21792
rect 29283 21732 29287 21788
rect 29287 21732 29343 21788
rect 29343 21732 29347 21788
rect 29283 21728 29347 21732
rect 29363 21788 29427 21792
rect 29363 21732 29367 21788
rect 29367 21732 29423 21788
rect 29423 21732 29427 21788
rect 29363 21728 29427 21732
rect 29443 21788 29507 21792
rect 29443 21732 29447 21788
rect 29447 21732 29503 21788
rect 29503 21732 29507 21788
rect 29443 21728 29507 21732
rect 29523 21788 29587 21792
rect 29523 21732 29527 21788
rect 29527 21732 29583 21788
rect 29583 21732 29587 21788
rect 29523 21728 29587 21732
rect 4493 21244 4557 21248
rect 4493 21188 4497 21244
rect 4497 21188 4553 21244
rect 4553 21188 4557 21244
rect 4493 21184 4557 21188
rect 4573 21244 4637 21248
rect 4573 21188 4577 21244
rect 4577 21188 4633 21244
rect 4633 21188 4637 21244
rect 4573 21184 4637 21188
rect 4653 21244 4717 21248
rect 4653 21188 4657 21244
rect 4657 21188 4713 21244
rect 4713 21188 4717 21244
rect 4653 21184 4717 21188
rect 4733 21244 4797 21248
rect 4733 21188 4737 21244
rect 4737 21188 4793 21244
rect 4793 21188 4797 21244
rect 4733 21184 4797 21188
rect 11576 21244 11640 21248
rect 11576 21188 11580 21244
rect 11580 21188 11636 21244
rect 11636 21188 11640 21244
rect 11576 21184 11640 21188
rect 11656 21244 11720 21248
rect 11656 21188 11660 21244
rect 11660 21188 11716 21244
rect 11716 21188 11720 21244
rect 11656 21184 11720 21188
rect 11736 21244 11800 21248
rect 11736 21188 11740 21244
rect 11740 21188 11796 21244
rect 11796 21188 11800 21244
rect 11736 21184 11800 21188
rect 11816 21244 11880 21248
rect 11816 21188 11820 21244
rect 11820 21188 11876 21244
rect 11876 21188 11880 21244
rect 11816 21184 11880 21188
rect 18659 21244 18723 21248
rect 18659 21188 18663 21244
rect 18663 21188 18719 21244
rect 18719 21188 18723 21244
rect 18659 21184 18723 21188
rect 18739 21244 18803 21248
rect 18739 21188 18743 21244
rect 18743 21188 18799 21244
rect 18799 21188 18803 21244
rect 18739 21184 18803 21188
rect 18819 21244 18883 21248
rect 18819 21188 18823 21244
rect 18823 21188 18879 21244
rect 18879 21188 18883 21244
rect 18819 21184 18883 21188
rect 18899 21244 18963 21248
rect 18899 21188 18903 21244
rect 18903 21188 18959 21244
rect 18959 21188 18963 21244
rect 18899 21184 18963 21188
rect 25742 21244 25806 21248
rect 25742 21188 25746 21244
rect 25746 21188 25802 21244
rect 25802 21188 25806 21244
rect 25742 21184 25806 21188
rect 25822 21244 25886 21248
rect 25822 21188 25826 21244
rect 25826 21188 25882 21244
rect 25882 21188 25886 21244
rect 25822 21184 25886 21188
rect 25902 21244 25966 21248
rect 25902 21188 25906 21244
rect 25906 21188 25962 21244
rect 25962 21188 25966 21244
rect 25902 21184 25966 21188
rect 25982 21244 26046 21248
rect 25982 21188 25986 21244
rect 25986 21188 26042 21244
rect 26042 21188 26046 21244
rect 25982 21184 26046 21188
rect 16252 20768 16316 20772
rect 16252 20712 16302 20768
rect 16302 20712 16316 20768
rect 16252 20708 16316 20712
rect 8034 20700 8098 20704
rect 8034 20644 8038 20700
rect 8038 20644 8094 20700
rect 8094 20644 8098 20700
rect 8034 20640 8098 20644
rect 8114 20700 8178 20704
rect 8114 20644 8118 20700
rect 8118 20644 8174 20700
rect 8174 20644 8178 20700
rect 8114 20640 8178 20644
rect 8194 20700 8258 20704
rect 8194 20644 8198 20700
rect 8198 20644 8254 20700
rect 8254 20644 8258 20700
rect 8194 20640 8258 20644
rect 8274 20700 8338 20704
rect 8274 20644 8278 20700
rect 8278 20644 8334 20700
rect 8334 20644 8338 20700
rect 8274 20640 8338 20644
rect 15117 20700 15181 20704
rect 15117 20644 15121 20700
rect 15121 20644 15177 20700
rect 15177 20644 15181 20700
rect 15117 20640 15181 20644
rect 15197 20700 15261 20704
rect 15197 20644 15201 20700
rect 15201 20644 15257 20700
rect 15257 20644 15261 20700
rect 15197 20640 15261 20644
rect 15277 20700 15341 20704
rect 15277 20644 15281 20700
rect 15281 20644 15337 20700
rect 15337 20644 15341 20700
rect 15277 20640 15341 20644
rect 15357 20700 15421 20704
rect 15357 20644 15361 20700
rect 15361 20644 15417 20700
rect 15417 20644 15421 20700
rect 15357 20640 15421 20644
rect 22200 20700 22264 20704
rect 22200 20644 22204 20700
rect 22204 20644 22260 20700
rect 22260 20644 22264 20700
rect 22200 20640 22264 20644
rect 22280 20700 22344 20704
rect 22280 20644 22284 20700
rect 22284 20644 22340 20700
rect 22340 20644 22344 20700
rect 22280 20640 22344 20644
rect 22360 20700 22424 20704
rect 22360 20644 22364 20700
rect 22364 20644 22420 20700
rect 22420 20644 22424 20700
rect 22360 20640 22424 20644
rect 22440 20700 22504 20704
rect 22440 20644 22444 20700
rect 22444 20644 22500 20700
rect 22500 20644 22504 20700
rect 22440 20640 22504 20644
rect 29283 20700 29347 20704
rect 29283 20644 29287 20700
rect 29287 20644 29343 20700
rect 29343 20644 29347 20700
rect 29283 20640 29347 20644
rect 29363 20700 29427 20704
rect 29363 20644 29367 20700
rect 29367 20644 29423 20700
rect 29423 20644 29427 20700
rect 29363 20640 29427 20644
rect 29443 20700 29507 20704
rect 29443 20644 29447 20700
rect 29447 20644 29503 20700
rect 29503 20644 29507 20700
rect 29443 20640 29507 20644
rect 29523 20700 29587 20704
rect 29523 20644 29527 20700
rect 29527 20644 29583 20700
rect 29583 20644 29587 20700
rect 29523 20640 29587 20644
rect 4493 20156 4557 20160
rect 4493 20100 4497 20156
rect 4497 20100 4553 20156
rect 4553 20100 4557 20156
rect 4493 20096 4557 20100
rect 4573 20156 4637 20160
rect 4573 20100 4577 20156
rect 4577 20100 4633 20156
rect 4633 20100 4637 20156
rect 4573 20096 4637 20100
rect 4653 20156 4717 20160
rect 4653 20100 4657 20156
rect 4657 20100 4713 20156
rect 4713 20100 4717 20156
rect 4653 20096 4717 20100
rect 4733 20156 4797 20160
rect 4733 20100 4737 20156
rect 4737 20100 4793 20156
rect 4793 20100 4797 20156
rect 4733 20096 4797 20100
rect 11576 20156 11640 20160
rect 11576 20100 11580 20156
rect 11580 20100 11636 20156
rect 11636 20100 11640 20156
rect 11576 20096 11640 20100
rect 11656 20156 11720 20160
rect 11656 20100 11660 20156
rect 11660 20100 11716 20156
rect 11716 20100 11720 20156
rect 11656 20096 11720 20100
rect 11736 20156 11800 20160
rect 11736 20100 11740 20156
rect 11740 20100 11796 20156
rect 11796 20100 11800 20156
rect 11736 20096 11800 20100
rect 11816 20156 11880 20160
rect 11816 20100 11820 20156
rect 11820 20100 11876 20156
rect 11876 20100 11880 20156
rect 11816 20096 11880 20100
rect 18659 20156 18723 20160
rect 18659 20100 18663 20156
rect 18663 20100 18719 20156
rect 18719 20100 18723 20156
rect 18659 20096 18723 20100
rect 18739 20156 18803 20160
rect 18739 20100 18743 20156
rect 18743 20100 18799 20156
rect 18799 20100 18803 20156
rect 18739 20096 18803 20100
rect 18819 20156 18883 20160
rect 18819 20100 18823 20156
rect 18823 20100 18879 20156
rect 18879 20100 18883 20156
rect 18819 20096 18883 20100
rect 18899 20156 18963 20160
rect 18899 20100 18903 20156
rect 18903 20100 18959 20156
rect 18959 20100 18963 20156
rect 18899 20096 18963 20100
rect 25742 20156 25806 20160
rect 25742 20100 25746 20156
rect 25746 20100 25802 20156
rect 25802 20100 25806 20156
rect 25742 20096 25806 20100
rect 25822 20156 25886 20160
rect 25822 20100 25826 20156
rect 25826 20100 25882 20156
rect 25882 20100 25886 20156
rect 25822 20096 25886 20100
rect 25902 20156 25966 20160
rect 25902 20100 25906 20156
rect 25906 20100 25962 20156
rect 25962 20100 25966 20156
rect 25902 20096 25966 20100
rect 25982 20156 26046 20160
rect 25982 20100 25986 20156
rect 25986 20100 26042 20156
rect 26042 20100 26046 20156
rect 25982 20096 26046 20100
rect 8034 19612 8098 19616
rect 8034 19556 8038 19612
rect 8038 19556 8094 19612
rect 8094 19556 8098 19612
rect 8034 19552 8098 19556
rect 8114 19612 8178 19616
rect 8114 19556 8118 19612
rect 8118 19556 8174 19612
rect 8174 19556 8178 19612
rect 8114 19552 8178 19556
rect 8194 19612 8258 19616
rect 8194 19556 8198 19612
rect 8198 19556 8254 19612
rect 8254 19556 8258 19612
rect 8194 19552 8258 19556
rect 8274 19612 8338 19616
rect 8274 19556 8278 19612
rect 8278 19556 8334 19612
rect 8334 19556 8338 19612
rect 8274 19552 8338 19556
rect 15117 19612 15181 19616
rect 15117 19556 15121 19612
rect 15121 19556 15177 19612
rect 15177 19556 15181 19612
rect 15117 19552 15181 19556
rect 15197 19612 15261 19616
rect 15197 19556 15201 19612
rect 15201 19556 15257 19612
rect 15257 19556 15261 19612
rect 15197 19552 15261 19556
rect 15277 19612 15341 19616
rect 15277 19556 15281 19612
rect 15281 19556 15337 19612
rect 15337 19556 15341 19612
rect 15277 19552 15341 19556
rect 15357 19612 15421 19616
rect 15357 19556 15361 19612
rect 15361 19556 15417 19612
rect 15417 19556 15421 19612
rect 15357 19552 15421 19556
rect 22200 19612 22264 19616
rect 22200 19556 22204 19612
rect 22204 19556 22260 19612
rect 22260 19556 22264 19612
rect 22200 19552 22264 19556
rect 22280 19612 22344 19616
rect 22280 19556 22284 19612
rect 22284 19556 22340 19612
rect 22340 19556 22344 19612
rect 22280 19552 22344 19556
rect 22360 19612 22424 19616
rect 22360 19556 22364 19612
rect 22364 19556 22420 19612
rect 22420 19556 22424 19612
rect 22360 19552 22424 19556
rect 22440 19612 22504 19616
rect 22440 19556 22444 19612
rect 22444 19556 22500 19612
rect 22500 19556 22504 19612
rect 22440 19552 22504 19556
rect 29283 19612 29347 19616
rect 29283 19556 29287 19612
rect 29287 19556 29343 19612
rect 29343 19556 29347 19612
rect 29283 19552 29347 19556
rect 29363 19612 29427 19616
rect 29363 19556 29367 19612
rect 29367 19556 29423 19612
rect 29423 19556 29427 19612
rect 29363 19552 29427 19556
rect 29443 19612 29507 19616
rect 29443 19556 29447 19612
rect 29447 19556 29503 19612
rect 29503 19556 29507 19612
rect 29443 19552 29507 19556
rect 29523 19612 29587 19616
rect 29523 19556 29527 19612
rect 29527 19556 29583 19612
rect 29583 19556 29587 19612
rect 29523 19552 29587 19556
rect 10180 19408 10244 19412
rect 10180 19352 10194 19408
rect 10194 19352 10244 19408
rect 10180 19348 10244 19352
rect 4493 19068 4557 19072
rect 4493 19012 4497 19068
rect 4497 19012 4553 19068
rect 4553 19012 4557 19068
rect 4493 19008 4557 19012
rect 4573 19068 4637 19072
rect 4573 19012 4577 19068
rect 4577 19012 4633 19068
rect 4633 19012 4637 19068
rect 4573 19008 4637 19012
rect 4653 19068 4717 19072
rect 4653 19012 4657 19068
rect 4657 19012 4713 19068
rect 4713 19012 4717 19068
rect 4653 19008 4717 19012
rect 4733 19068 4797 19072
rect 4733 19012 4737 19068
rect 4737 19012 4793 19068
rect 4793 19012 4797 19068
rect 4733 19008 4797 19012
rect 11576 19068 11640 19072
rect 11576 19012 11580 19068
rect 11580 19012 11636 19068
rect 11636 19012 11640 19068
rect 11576 19008 11640 19012
rect 11656 19068 11720 19072
rect 11656 19012 11660 19068
rect 11660 19012 11716 19068
rect 11716 19012 11720 19068
rect 11656 19008 11720 19012
rect 11736 19068 11800 19072
rect 11736 19012 11740 19068
rect 11740 19012 11796 19068
rect 11796 19012 11800 19068
rect 11736 19008 11800 19012
rect 11816 19068 11880 19072
rect 11816 19012 11820 19068
rect 11820 19012 11876 19068
rect 11876 19012 11880 19068
rect 11816 19008 11880 19012
rect 18659 19068 18723 19072
rect 18659 19012 18663 19068
rect 18663 19012 18719 19068
rect 18719 19012 18723 19068
rect 18659 19008 18723 19012
rect 18739 19068 18803 19072
rect 18739 19012 18743 19068
rect 18743 19012 18799 19068
rect 18799 19012 18803 19068
rect 18739 19008 18803 19012
rect 18819 19068 18883 19072
rect 18819 19012 18823 19068
rect 18823 19012 18879 19068
rect 18879 19012 18883 19068
rect 18819 19008 18883 19012
rect 18899 19068 18963 19072
rect 18899 19012 18903 19068
rect 18903 19012 18959 19068
rect 18959 19012 18963 19068
rect 18899 19008 18963 19012
rect 25742 19068 25806 19072
rect 25742 19012 25746 19068
rect 25746 19012 25802 19068
rect 25802 19012 25806 19068
rect 25742 19008 25806 19012
rect 25822 19068 25886 19072
rect 25822 19012 25826 19068
rect 25826 19012 25882 19068
rect 25882 19012 25886 19068
rect 25822 19008 25886 19012
rect 25902 19068 25966 19072
rect 25902 19012 25906 19068
rect 25906 19012 25962 19068
rect 25962 19012 25966 19068
rect 25902 19008 25966 19012
rect 25982 19068 26046 19072
rect 25982 19012 25986 19068
rect 25986 19012 26042 19068
rect 26042 19012 26046 19068
rect 25982 19008 26046 19012
rect 8034 18524 8098 18528
rect 8034 18468 8038 18524
rect 8038 18468 8094 18524
rect 8094 18468 8098 18524
rect 8034 18464 8098 18468
rect 8114 18524 8178 18528
rect 8114 18468 8118 18524
rect 8118 18468 8174 18524
rect 8174 18468 8178 18524
rect 8114 18464 8178 18468
rect 8194 18524 8258 18528
rect 8194 18468 8198 18524
rect 8198 18468 8254 18524
rect 8254 18468 8258 18524
rect 8194 18464 8258 18468
rect 8274 18524 8338 18528
rect 8274 18468 8278 18524
rect 8278 18468 8334 18524
rect 8334 18468 8338 18524
rect 8274 18464 8338 18468
rect 15117 18524 15181 18528
rect 15117 18468 15121 18524
rect 15121 18468 15177 18524
rect 15177 18468 15181 18524
rect 15117 18464 15181 18468
rect 15197 18524 15261 18528
rect 15197 18468 15201 18524
rect 15201 18468 15257 18524
rect 15257 18468 15261 18524
rect 15197 18464 15261 18468
rect 15277 18524 15341 18528
rect 15277 18468 15281 18524
rect 15281 18468 15337 18524
rect 15337 18468 15341 18524
rect 15277 18464 15341 18468
rect 15357 18524 15421 18528
rect 15357 18468 15361 18524
rect 15361 18468 15417 18524
rect 15417 18468 15421 18524
rect 15357 18464 15421 18468
rect 22200 18524 22264 18528
rect 22200 18468 22204 18524
rect 22204 18468 22260 18524
rect 22260 18468 22264 18524
rect 22200 18464 22264 18468
rect 22280 18524 22344 18528
rect 22280 18468 22284 18524
rect 22284 18468 22340 18524
rect 22340 18468 22344 18524
rect 22280 18464 22344 18468
rect 22360 18524 22424 18528
rect 22360 18468 22364 18524
rect 22364 18468 22420 18524
rect 22420 18468 22424 18524
rect 22360 18464 22424 18468
rect 22440 18524 22504 18528
rect 22440 18468 22444 18524
rect 22444 18468 22500 18524
rect 22500 18468 22504 18524
rect 22440 18464 22504 18468
rect 29283 18524 29347 18528
rect 29283 18468 29287 18524
rect 29287 18468 29343 18524
rect 29343 18468 29347 18524
rect 29283 18464 29347 18468
rect 29363 18524 29427 18528
rect 29363 18468 29367 18524
rect 29367 18468 29423 18524
rect 29423 18468 29427 18524
rect 29363 18464 29427 18468
rect 29443 18524 29507 18528
rect 29443 18468 29447 18524
rect 29447 18468 29503 18524
rect 29503 18468 29507 18524
rect 29443 18464 29507 18468
rect 29523 18524 29587 18528
rect 29523 18468 29527 18524
rect 29527 18468 29583 18524
rect 29583 18468 29587 18524
rect 29523 18464 29587 18468
rect 4493 17980 4557 17984
rect 4493 17924 4497 17980
rect 4497 17924 4553 17980
rect 4553 17924 4557 17980
rect 4493 17920 4557 17924
rect 4573 17980 4637 17984
rect 4573 17924 4577 17980
rect 4577 17924 4633 17980
rect 4633 17924 4637 17980
rect 4573 17920 4637 17924
rect 4653 17980 4717 17984
rect 4653 17924 4657 17980
rect 4657 17924 4713 17980
rect 4713 17924 4717 17980
rect 4653 17920 4717 17924
rect 4733 17980 4797 17984
rect 4733 17924 4737 17980
rect 4737 17924 4793 17980
rect 4793 17924 4797 17980
rect 4733 17920 4797 17924
rect 11576 17980 11640 17984
rect 11576 17924 11580 17980
rect 11580 17924 11636 17980
rect 11636 17924 11640 17980
rect 11576 17920 11640 17924
rect 11656 17980 11720 17984
rect 11656 17924 11660 17980
rect 11660 17924 11716 17980
rect 11716 17924 11720 17980
rect 11656 17920 11720 17924
rect 11736 17980 11800 17984
rect 11736 17924 11740 17980
rect 11740 17924 11796 17980
rect 11796 17924 11800 17980
rect 11736 17920 11800 17924
rect 11816 17980 11880 17984
rect 11816 17924 11820 17980
rect 11820 17924 11876 17980
rect 11876 17924 11880 17980
rect 11816 17920 11880 17924
rect 18659 17980 18723 17984
rect 18659 17924 18663 17980
rect 18663 17924 18719 17980
rect 18719 17924 18723 17980
rect 18659 17920 18723 17924
rect 18739 17980 18803 17984
rect 18739 17924 18743 17980
rect 18743 17924 18799 17980
rect 18799 17924 18803 17980
rect 18739 17920 18803 17924
rect 18819 17980 18883 17984
rect 18819 17924 18823 17980
rect 18823 17924 18879 17980
rect 18879 17924 18883 17980
rect 18819 17920 18883 17924
rect 18899 17980 18963 17984
rect 18899 17924 18903 17980
rect 18903 17924 18959 17980
rect 18959 17924 18963 17980
rect 18899 17920 18963 17924
rect 25742 17980 25806 17984
rect 25742 17924 25746 17980
rect 25746 17924 25802 17980
rect 25802 17924 25806 17980
rect 25742 17920 25806 17924
rect 25822 17980 25886 17984
rect 25822 17924 25826 17980
rect 25826 17924 25882 17980
rect 25882 17924 25886 17980
rect 25822 17920 25886 17924
rect 25902 17980 25966 17984
rect 25902 17924 25906 17980
rect 25906 17924 25962 17980
rect 25962 17924 25966 17980
rect 25902 17920 25966 17924
rect 25982 17980 26046 17984
rect 25982 17924 25986 17980
rect 25986 17924 26042 17980
rect 26042 17924 26046 17980
rect 25982 17920 26046 17924
rect 8034 17436 8098 17440
rect 8034 17380 8038 17436
rect 8038 17380 8094 17436
rect 8094 17380 8098 17436
rect 8034 17376 8098 17380
rect 8114 17436 8178 17440
rect 8114 17380 8118 17436
rect 8118 17380 8174 17436
rect 8174 17380 8178 17436
rect 8114 17376 8178 17380
rect 8194 17436 8258 17440
rect 8194 17380 8198 17436
rect 8198 17380 8254 17436
rect 8254 17380 8258 17436
rect 8194 17376 8258 17380
rect 8274 17436 8338 17440
rect 8274 17380 8278 17436
rect 8278 17380 8334 17436
rect 8334 17380 8338 17436
rect 8274 17376 8338 17380
rect 15117 17436 15181 17440
rect 15117 17380 15121 17436
rect 15121 17380 15177 17436
rect 15177 17380 15181 17436
rect 15117 17376 15181 17380
rect 15197 17436 15261 17440
rect 15197 17380 15201 17436
rect 15201 17380 15257 17436
rect 15257 17380 15261 17436
rect 15197 17376 15261 17380
rect 15277 17436 15341 17440
rect 15277 17380 15281 17436
rect 15281 17380 15337 17436
rect 15337 17380 15341 17436
rect 15277 17376 15341 17380
rect 15357 17436 15421 17440
rect 15357 17380 15361 17436
rect 15361 17380 15417 17436
rect 15417 17380 15421 17436
rect 15357 17376 15421 17380
rect 22200 17436 22264 17440
rect 22200 17380 22204 17436
rect 22204 17380 22260 17436
rect 22260 17380 22264 17436
rect 22200 17376 22264 17380
rect 22280 17436 22344 17440
rect 22280 17380 22284 17436
rect 22284 17380 22340 17436
rect 22340 17380 22344 17436
rect 22280 17376 22344 17380
rect 22360 17436 22424 17440
rect 22360 17380 22364 17436
rect 22364 17380 22420 17436
rect 22420 17380 22424 17436
rect 22360 17376 22424 17380
rect 22440 17436 22504 17440
rect 22440 17380 22444 17436
rect 22444 17380 22500 17436
rect 22500 17380 22504 17436
rect 22440 17376 22504 17380
rect 29283 17436 29347 17440
rect 29283 17380 29287 17436
rect 29287 17380 29343 17436
rect 29343 17380 29347 17436
rect 29283 17376 29347 17380
rect 29363 17436 29427 17440
rect 29363 17380 29367 17436
rect 29367 17380 29423 17436
rect 29423 17380 29427 17436
rect 29363 17376 29427 17380
rect 29443 17436 29507 17440
rect 29443 17380 29447 17436
rect 29447 17380 29503 17436
rect 29503 17380 29507 17436
rect 29443 17376 29507 17380
rect 29523 17436 29587 17440
rect 29523 17380 29527 17436
rect 29527 17380 29583 17436
rect 29583 17380 29587 17436
rect 29523 17376 29587 17380
rect 27660 17232 27724 17236
rect 27660 17176 27710 17232
rect 27710 17176 27724 17232
rect 27660 17172 27724 17176
rect 4493 16892 4557 16896
rect 4493 16836 4497 16892
rect 4497 16836 4553 16892
rect 4553 16836 4557 16892
rect 4493 16832 4557 16836
rect 4573 16892 4637 16896
rect 4573 16836 4577 16892
rect 4577 16836 4633 16892
rect 4633 16836 4637 16892
rect 4573 16832 4637 16836
rect 4653 16892 4717 16896
rect 4653 16836 4657 16892
rect 4657 16836 4713 16892
rect 4713 16836 4717 16892
rect 4653 16832 4717 16836
rect 4733 16892 4797 16896
rect 4733 16836 4737 16892
rect 4737 16836 4793 16892
rect 4793 16836 4797 16892
rect 4733 16832 4797 16836
rect 11576 16892 11640 16896
rect 11576 16836 11580 16892
rect 11580 16836 11636 16892
rect 11636 16836 11640 16892
rect 11576 16832 11640 16836
rect 11656 16892 11720 16896
rect 11656 16836 11660 16892
rect 11660 16836 11716 16892
rect 11716 16836 11720 16892
rect 11656 16832 11720 16836
rect 11736 16892 11800 16896
rect 11736 16836 11740 16892
rect 11740 16836 11796 16892
rect 11796 16836 11800 16892
rect 11736 16832 11800 16836
rect 11816 16892 11880 16896
rect 11816 16836 11820 16892
rect 11820 16836 11876 16892
rect 11876 16836 11880 16892
rect 11816 16832 11880 16836
rect 18659 16892 18723 16896
rect 18659 16836 18663 16892
rect 18663 16836 18719 16892
rect 18719 16836 18723 16892
rect 18659 16832 18723 16836
rect 18739 16892 18803 16896
rect 18739 16836 18743 16892
rect 18743 16836 18799 16892
rect 18799 16836 18803 16892
rect 18739 16832 18803 16836
rect 18819 16892 18883 16896
rect 18819 16836 18823 16892
rect 18823 16836 18879 16892
rect 18879 16836 18883 16892
rect 18819 16832 18883 16836
rect 18899 16892 18963 16896
rect 18899 16836 18903 16892
rect 18903 16836 18959 16892
rect 18959 16836 18963 16892
rect 18899 16832 18963 16836
rect 25742 16892 25806 16896
rect 25742 16836 25746 16892
rect 25746 16836 25802 16892
rect 25802 16836 25806 16892
rect 25742 16832 25806 16836
rect 25822 16892 25886 16896
rect 25822 16836 25826 16892
rect 25826 16836 25882 16892
rect 25882 16836 25886 16892
rect 25822 16832 25886 16836
rect 25902 16892 25966 16896
rect 25902 16836 25906 16892
rect 25906 16836 25962 16892
rect 25962 16836 25966 16892
rect 25902 16832 25966 16836
rect 25982 16892 26046 16896
rect 25982 16836 25986 16892
rect 25986 16836 26042 16892
rect 26042 16836 26046 16892
rect 25982 16832 26046 16836
rect 8034 16348 8098 16352
rect 8034 16292 8038 16348
rect 8038 16292 8094 16348
rect 8094 16292 8098 16348
rect 8034 16288 8098 16292
rect 8114 16348 8178 16352
rect 8114 16292 8118 16348
rect 8118 16292 8174 16348
rect 8174 16292 8178 16348
rect 8114 16288 8178 16292
rect 8194 16348 8258 16352
rect 8194 16292 8198 16348
rect 8198 16292 8254 16348
rect 8254 16292 8258 16348
rect 8194 16288 8258 16292
rect 8274 16348 8338 16352
rect 8274 16292 8278 16348
rect 8278 16292 8334 16348
rect 8334 16292 8338 16348
rect 8274 16288 8338 16292
rect 15117 16348 15181 16352
rect 15117 16292 15121 16348
rect 15121 16292 15177 16348
rect 15177 16292 15181 16348
rect 15117 16288 15181 16292
rect 15197 16348 15261 16352
rect 15197 16292 15201 16348
rect 15201 16292 15257 16348
rect 15257 16292 15261 16348
rect 15197 16288 15261 16292
rect 15277 16348 15341 16352
rect 15277 16292 15281 16348
rect 15281 16292 15337 16348
rect 15337 16292 15341 16348
rect 15277 16288 15341 16292
rect 15357 16348 15421 16352
rect 15357 16292 15361 16348
rect 15361 16292 15417 16348
rect 15417 16292 15421 16348
rect 15357 16288 15421 16292
rect 22200 16348 22264 16352
rect 22200 16292 22204 16348
rect 22204 16292 22260 16348
rect 22260 16292 22264 16348
rect 22200 16288 22264 16292
rect 22280 16348 22344 16352
rect 22280 16292 22284 16348
rect 22284 16292 22340 16348
rect 22340 16292 22344 16348
rect 22280 16288 22344 16292
rect 22360 16348 22424 16352
rect 22360 16292 22364 16348
rect 22364 16292 22420 16348
rect 22420 16292 22424 16348
rect 22360 16288 22424 16292
rect 22440 16348 22504 16352
rect 22440 16292 22444 16348
rect 22444 16292 22500 16348
rect 22500 16292 22504 16348
rect 22440 16288 22504 16292
rect 29283 16348 29347 16352
rect 29283 16292 29287 16348
rect 29287 16292 29343 16348
rect 29343 16292 29347 16348
rect 29283 16288 29347 16292
rect 29363 16348 29427 16352
rect 29363 16292 29367 16348
rect 29367 16292 29423 16348
rect 29423 16292 29427 16348
rect 29363 16288 29427 16292
rect 29443 16348 29507 16352
rect 29443 16292 29447 16348
rect 29447 16292 29503 16348
rect 29503 16292 29507 16348
rect 29443 16288 29507 16292
rect 29523 16348 29587 16352
rect 29523 16292 29527 16348
rect 29527 16292 29583 16348
rect 29583 16292 29587 16348
rect 29523 16288 29587 16292
rect 4493 15804 4557 15808
rect 4493 15748 4497 15804
rect 4497 15748 4553 15804
rect 4553 15748 4557 15804
rect 4493 15744 4557 15748
rect 4573 15804 4637 15808
rect 4573 15748 4577 15804
rect 4577 15748 4633 15804
rect 4633 15748 4637 15804
rect 4573 15744 4637 15748
rect 4653 15804 4717 15808
rect 4653 15748 4657 15804
rect 4657 15748 4713 15804
rect 4713 15748 4717 15804
rect 4653 15744 4717 15748
rect 4733 15804 4797 15808
rect 4733 15748 4737 15804
rect 4737 15748 4793 15804
rect 4793 15748 4797 15804
rect 4733 15744 4797 15748
rect 11576 15804 11640 15808
rect 11576 15748 11580 15804
rect 11580 15748 11636 15804
rect 11636 15748 11640 15804
rect 11576 15744 11640 15748
rect 11656 15804 11720 15808
rect 11656 15748 11660 15804
rect 11660 15748 11716 15804
rect 11716 15748 11720 15804
rect 11656 15744 11720 15748
rect 11736 15804 11800 15808
rect 11736 15748 11740 15804
rect 11740 15748 11796 15804
rect 11796 15748 11800 15804
rect 11736 15744 11800 15748
rect 11816 15804 11880 15808
rect 11816 15748 11820 15804
rect 11820 15748 11876 15804
rect 11876 15748 11880 15804
rect 11816 15744 11880 15748
rect 18659 15804 18723 15808
rect 18659 15748 18663 15804
rect 18663 15748 18719 15804
rect 18719 15748 18723 15804
rect 18659 15744 18723 15748
rect 18739 15804 18803 15808
rect 18739 15748 18743 15804
rect 18743 15748 18799 15804
rect 18799 15748 18803 15804
rect 18739 15744 18803 15748
rect 18819 15804 18883 15808
rect 18819 15748 18823 15804
rect 18823 15748 18879 15804
rect 18879 15748 18883 15804
rect 18819 15744 18883 15748
rect 18899 15804 18963 15808
rect 18899 15748 18903 15804
rect 18903 15748 18959 15804
rect 18959 15748 18963 15804
rect 18899 15744 18963 15748
rect 25742 15804 25806 15808
rect 25742 15748 25746 15804
rect 25746 15748 25802 15804
rect 25802 15748 25806 15804
rect 25742 15744 25806 15748
rect 25822 15804 25886 15808
rect 25822 15748 25826 15804
rect 25826 15748 25882 15804
rect 25882 15748 25886 15804
rect 25822 15744 25886 15748
rect 25902 15804 25966 15808
rect 25902 15748 25906 15804
rect 25906 15748 25962 15804
rect 25962 15748 25966 15804
rect 25902 15744 25966 15748
rect 25982 15804 26046 15808
rect 25982 15748 25986 15804
rect 25986 15748 26042 15804
rect 26042 15748 26046 15804
rect 25982 15744 26046 15748
rect 8034 15260 8098 15264
rect 8034 15204 8038 15260
rect 8038 15204 8094 15260
rect 8094 15204 8098 15260
rect 8034 15200 8098 15204
rect 8114 15260 8178 15264
rect 8114 15204 8118 15260
rect 8118 15204 8174 15260
rect 8174 15204 8178 15260
rect 8114 15200 8178 15204
rect 8194 15260 8258 15264
rect 8194 15204 8198 15260
rect 8198 15204 8254 15260
rect 8254 15204 8258 15260
rect 8194 15200 8258 15204
rect 8274 15260 8338 15264
rect 8274 15204 8278 15260
rect 8278 15204 8334 15260
rect 8334 15204 8338 15260
rect 8274 15200 8338 15204
rect 15117 15260 15181 15264
rect 15117 15204 15121 15260
rect 15121 15204 15177 15260
rect 15177 15204 15181 15260
rect 15117 15200 15181 15204
rect 15197 15260 15261 15264
rect 15197 15204 15201 15260
rect 15201 15204 15257 15260
rect 15257 15204 15261 15260
rect 15197 15200 15261 15204
rect 15277 15260 15341 15264
rect 15277 15204 15281 15260
rect 15281 15204 15337 15260
rect 15337 15204 15341 15260
rect 15277 15200 15341 15204
rect 15357 15260 15421 15264
rect 15357 15204 15361 15260
rect 15361 15204 15417 15260
rect 15417 15204 15421 15260
rect 15357 15200 15421 15204
rect 22200 15260 22264 15264
rect 22200 15204 22204 15260
rect 22204 15204 22260 15260
rect 22260 15204 22264 15260
rect 22200 15200 22264 15204
rect 22280 15260 22344 15264
rect 22280 15204 22284 15260
rect 22284 15204 22340 15260
rect 22340 15204 22344 15260
rect 22280 15200 22344 15204
rect 22360 15260 22424 15264
rect 22360 15204 22364 15260
rect 22364 15204 22420 15260
rect 22420 15204 22424 15260
rect 22360 15200 22424 15204
rect 22440 15260 22504 15264
rect 22440 15204 22444 15260
rect 22444 15204 22500 15260
rect 22500 15204 22504 15260
rect 22440 15200 22504 15204
rect 29283 15260 29347 15264
rect 29283 15204 29287 15260
rect 29287 15204 29343 15260
rect 29343 15204 29347 15260
rect 29283 15200 29347 15204
rect 29363 15260 29427 15264
rect 29363 15204 29367 15260
rect 29367 15204 29423 15260
rect 29423 15204 29427 15260
rect 29363 15200 29427 15204
rect 29443 15260 29507 15264
rect 29443 15204 29447 15260
rect 29447 15204 29503 15260
rect 29503 15204 29507 15260
rect 29443 15200 29507 15204
rect 29523 15260 29587 15264
rect 29523 15204 29527 15260
rect 29527 15204 29583 15260
rect 29583 15204 29587 15260
rect 29523 15200 29587 15204
rect 16252 15192 16316 15196
rect 16252 15136 16302 15192
rect 16302 15136 16316 15192
rect 16252 15132 16316 15136
rect 4493 14716 4557 14720
rect 4493 14660 4497 14716
rect 4497 14660 4553 14716
rect 4553 14660 4557 14716
rect 4493 14656 4557 14660
rect 4573 14716 4637 14720
rect 4573 14660 4577 14716
rect 4577 14660 4633 14716
rect 4633 14660 4637 14716
rect 4573 14656 4637 14660
rect 4653 14716 4717 14720
rect 4653 14660 4657 14716
rect 4657 14660 4713 14716
rect 4713 14660 4717 14716
rect 4653 14656 4717 14660
rect 4733 14716 4797 14720
rect 4733 14660 4737 14716
rect 4737 14660 4793 14716
rect 4793 14660 4797 14716
rect 4733 14656 4797 14660
rect 11576 14716 11640 14720
rect 11576 14660 11580 14716
rect 11580 14660 11636 14716
rect 11636 14660 11640 14716
rect 11576 14656 11640 14660
rect 11656 14716 11720 14720
rect 11656 14660 11660 14716
rect 11660 14660 11716 14716
rect 11716 14660 11720 14716
rect 11656 14656 11720 14660
rect 11736 14716 11800 14720
rect 11736 14660 11740 14716
rect 11740 14660 11796 14716
rect 11796 14660 11800 14716
rect 11736 14656 11800 14660
rect 11816 14716 11880 14720
rect 11816 14660 11820 14716
rect 11820 14660 11876 14716
rect 11876 14660 11880 14716
rect 11816 14656 11880 14660
rect 18659 14716 18723 14720
rect 18659 14660 18663 14716
rect 18663 14660 18719 14716
rect 18719 14660 18723 14716
rect 18659 14656 18723 14660
rect 18739 14716 18803 14720
rect 18739 14660 18743 14716
rect 18743 14660 18799 14716
rect 18799 14660 18803 14716
rect 18739 14656 18803 14660
rect 18819 14716 18883 14720
rect 18819 14660 18823 14716
rect 18823 14660 18879 14716
rect 18879 14660 18883 14716
rect 18819 14656 18883 14660
rect 18899 14716 18963 14720
rect 18899 14660 18903 14716
rect 18903 14660 18959 14716
rect 18959 14660 18963 14716
rect 18899 14656 18963 14660
rect 25742 14716 25806 14720
rect 25742 14660 25746 14716
rect 25746 14660 25802 14716
rect 25802 14660 25806 14716
rect 25742 14656 25806 14660
rect 25822 14716 25886 14720
rect 25822 14660 25826 14716
rect 25826 14660 25882 14716
rect 25882 14660 25886 14716
rect 25822 14656 25886 14660
rect 25902 14716 25966 14720
rect 25902 14660 25906 14716
rect 25906 14660 25962 14716
rect 25962 14660 25966 14716
rect 25902 14656 25966 14660
rect 25982 14716 26046 14720
rect 25982 14660 25986 14716
rect 25986 14660 26042 14716
rect 26042 14660 26046 14716
rect 25982 14656 26046 14660
rect 8034 14172 8098 14176
rect 8034 14116 8038 14172
rect 8038 14116 8094 14172
rect 8094 14116 8098 14172
rect 8034 14112 8098 14116
rect 8114 14172 8178 14176
rect 8114 14116 8118 14172
rect 8118 14116 8174 14172
rect 8174 14116 8178 14172
rect 8114 14112 8178 14116
rect 8194 14172 8258 14176
rect 8194 14116 8198 14172
rect 8198 14116 8254 14172
rect 8254 14116 8258 14172
rect 8194 14112 8258 14116
rect 8274 14172 8338 14176
rect 8274 14116 8278 14172
rect 8278 14116 8334 14172
rect 8334 14116 8338 14172
rect 8274 14112 8338 14116
rect 15117 14172 15181 14176
rect 15117 14116 15121 14172
rect 15121 14116 15177 14172
rect 15177 14116 15181 14172
rect 15117 14112 15181 14116
rect 15197 14172 15261 14176
rect 15197 14116 15201 14172
rect 15201 14116 15257 14172
rect 15257 14116 15261 14172
rect 15197 14112 15261 14116
rect 15277 14172 15341 14176
rect 15277 14116 15281 14172
rect 15281 14116 15337 14172
rect 15337 14116 15341 14172
rect 15277 14112 15341 14116
rect 15357 14172 15421 14176
rect 15357 14116 15361 14172
rect 15361 14116 15417 14172
rect 15417 14116 15421 14172
rect 15357 14112 15421 14116
rect 22200 14172 22264 14176
rect 22200 14116 22204 14172
rect 22204 14116 22260 14172
rect 22260 14116 22264 14172
rect 22200 14112 22264 14116
rect 22280 14172 22344 14176
rect 22280 14116 22284 14172
rect 22284 14116 22340 14172
rect 22340 14116 22344 14172
rect 22280 14112 22344 14116
rect 22360 14172 22424 14176
rect 22360 14116 22364 14172
rect 22364 14116 22420 14172
rect 22420 14116 22424 14172
rect 22360 14112 22424 14116
rect 22440 14172 22504 14176
rect 22440 14116 22444 14172
rect 22444 14116 22500 14172
rect 22500 14116 22504 14172
rect 22440 14112 22504 14116
rect 29283 14172 29347 14176
rect 29283 14116 29287 14172
rect 29287 14116 29343 14172
rect 29343 14116 29347 14172
rect 29283 14112 29347 14116
rect 29363 14172 29427 14176
rect 29363 14116 29367 14172
rect 29367 14116 29423 14172
rect 29423 14116 29427 14172
rect 29363 14112 29427 14116
rect 29443 14172 29507 14176
rect 29443 14116 29447 14172
rect 29447 14116 29503 14172
rect 29503 14116 29507 14172
rect 29443 14112 29507 14116
rect 29523 14172 29587 14176
rect 29523 14116 29527 14172
rect 29527 14116 29583 14172
rect 29583 14116 29587 14172
rect 29523 14112 29587 14116
rect 4493 13628 4557 13632
rect 4493 13572 4497 13628
rect 4497 13572 4553 13628
rect 4553 13572 4557 13628
rect 4493 13568 4557 13572
rect 4573 13628 4637 13632
rect 4573 13572 4577 13628
rect 4577 13572 4633 13628
rect 4633 13572 4637 13628
rect 4573 13568 4637 13572
rect 4653 13628 4717 13632
rect 4653 13572 4657 13628
rect 4657 13572 4713 13628
rect 4713 13572 4717 13628
rect 4653 13568 4717 13572
rect 4733 13628 4797 13632
rect 4733 13572 4737 13628
rect 4737 13572 4793 13628
rect 4793 13572 4797 13628
rect 4733 13568 4797 13572
rect 11576 13628 11640 13632
rect 11576 13572 11580 13628
rect 11580 13572 11636 13628
rect 11636 13572 11640 13628
rect 11576 13568 11640 13572
rect 11656 13628 11720 13632
rect 11656 13572 11660 13628
rect 11660 13572 11716 13628
rect 11716 13572 11720 13628
rect 11656 13568 11720 13572
rect 11736 13628 11800 13632
rect 11736 13572 11740 13628
rect 11740 13572 11796 13628
rect 11796 13572 11800 13628
rect 11736 13568 11800 13572
rect 11816 13628 11880 13632
rect 11816 13572 11820 13628
rect 11820 13572 11876 13628
rect 11876 13572 11880 13628
rect 11816 13568 11880 13572
rect 18659 13628 18723 13632
rect 18659 13572 18663 13628
rect 18663 13572 18719 13628
rect 18719 13572 18723 13628
rect 18659 13568 18723 13572
rect 18739 13628 18803 13632
rect 18739 13572 18743 13628
rect 18743 13572 18799 13628
rect 18799 13572 18803 13628
rect 18739 13568 18803 13572
rect 18819 13628 18883 13632
rect 18819 13572 18823 13628
rect 18823 13572 18879 13628
rect 18879 13572 18883 13628
rect 18819 13568 18883 13572
rect 18899 13628 18963 13632
rect 18899 13572 18903 13628
rect 18903 13572 18959 13628
rect 18959 13572 18963 13628
rect 18899 13568 18963 13572
rect 25742 13628 25806 13632
rect 25742 13572 25746 13628
rect 25746 13572 25802 13628
rect 25802 13572 25806 13628
rect 25742 13568 25806 13572
rect 25822 13628 25886 13632
rect 25822 13572 25826 13628
rect 25826 13572 25882 13628
rect 25882 13572 25886 13628
rect 25822 13568 25886 13572
rect 25902 13628 25966 13632
rect 25902 13572 25906 13628
rect 25906 13572 25962 13628
rect 25962 13572 25966 13628
rect 25902 13568 25966 13572
rect 25982 13628 26046 13632
rect 25982 13572 25986 13628
rect 25986 13572 26042 13628
rect 26042 13572 26046 13628
rect 25982 13568 26046 13572
rect 10548 13228 10612 13292
rect 8034 13084 8098 13088
rect 8034 13028 8038 13084
rect 8038 13028 8094 13084
rect 8094 13028 8098 13084
rect 8034 13024 8098 13028
rect 8114 13084 8178 13088
rect 8114 13028 8118 13084
rect 8118 13028 8174 13084
rect 8174 13028 8178 13084
rect 8114 13024 8178 13028
rect 8194 13084 8258 13088
rect 8194 13028 8198 13084
rect 8198 13028 8254 13084
rect 8254 13028 8258 13084
rect 8194 13024 8258 13028
rect 8274 13084 8338 13088
rect 8274 13028 8278 13084
rect 8278 13028 8334 13084
rect 8334 13028 8338 13084
rect 8274 13024 8338 13028
rect 15117 13084 15181 13088
rect 15117 13028 15121 13084
rect 15121 13028 15177 13084
rect 15177 13028 15181 13084
rect 15117 13024 15181 13028
rect 15197 13084 15261 13088
rect 15197 13028 15201 13084
rect 15201 13028 15257 13084
rect 15257 13028 15261 13084
rect 15197 13024 15261 13028
rect 15277 13084 15341 13088
rect 15277 13028 15281 13084
rect 15281 13028 15337 13084
rect 15337 13028 15341 13084
rect 15277 13024 15341 13028
rect 15357 13084 15421 13088
rect 15357 13028 15361 13084
rect 15361 13028 15417 13084
rect 15417 13028 15421 13084
rect 15357 13024 15421 13028
rect 22200 13084 22264 13088
rect 22200 13028 22204 13084
rect 22204 13028 22260 13084
rect 22260 13028 22264 13084
rect 22200 13024 22264 13028
rect 22280 13084 22344 13088
rect 22280 13028 22284 13084
rect 22284 13028 22340 13084
rect 22340 13028 22344 13084
rect 22280 13024 22344 13028
rect 22360 13084 22424 13088
rect 22360 13028 22364 13084
rect 22364 13028 22420 13084
rect 22420 13028 22424 13084
rect 22360 13024 22424 13028
rect 22440 13084 22504 13088
rect 22440 13028 22444 13084
rect 22444 13028 22500 13084
rect 22500 13028 22504 13084
rect 22440 13024 22504 13028
rect 29283 13084 29347 13088
rect 29283 13028 29287 13084
rect 29287 13028 29343 13084
rect 29343 13028 29347 13084
rect 29283 13024 29347 13028
rect 29363 13084 29427 13088
rect 29363 13028 29367 13084
rect 29367 13028 29423 13084
rect 29423 13028 29427 13084
rect 29363 13024 29427 13028
rect 29443 13084 29507 13088
rect 29443 13028 29447 13084
rect 29447 13028 29503 13084
rect 29503 13028 29507 13084
rect 29443 13024 29507 13028
rect 29523 13084 29587 13088
rect 29523 13028 29527 13084
rect 29527 13028 29583 13084
rect 29583 13028 29587 13084
rect 29523 13024 29587 13028
rect 4493 12540 4557 12544
rect 4493 12484 4497 12540
rect 4497 12484 4553 12540
rect 4553 12484 4557 12540
rect 4493 12480 4557 12484
rect 4573 12540 4637 12544
rect 4573 12484 4577 12540
rect 4577 12484 4633 12540
rect 4633 12484 4637 12540
rect 4573 12480 4637 12484
rect 4653 12540 4717 12544
rect 4653 12484 4657 12540
rect 4657 12484 4713 12540
rect 4713 12484 4717 12540
rect 4653 12480 4717 12484
rect 4733 12540 4797 12544
rect 4733 12484 4737 12540
rect 4737 12484 4793 12540
rect 4793 12484 4797 12540
rect 4733 12480 4797 12484
rect 11576 12540 11640 12544
rect 11576 12484 11580 12540
rect 11580 12484 11636 12540
rect 11636 12484 11640 12540
rect 11576 12480 11640 12484
rect 11656 12540 11720 12544
rect 11656 12484 11660 12540
rect 11660 12484 11716 12540
rect 11716 12484 11720 12540
rect 11656 12480 11720 12484
rect 11736 12540 11800 12544
rect 11736 12484 11740 12540
rect 11740 12484 11796 12540
rect 11796 12484 11800 12540
rect 11736 12480 11800 12484
rect 11816 12540 11880 12544
rect 11816 12484 11820 12540
rect 11820 12484 11876 12540
rect 11876 12484 11880 12540
rect 11816 12480 11880 12484
rect 18659 12540 18723 12544
rect 18659 12484 18663 12540
rect 18663 12484 18719 12540
rect 18719 12484 18723 12540
rect 18659 12480 18723 12484
rect 18739 12540 18803 12544
rect 18739 12484 18743 12540
rect 18743 12484 18799 12540
rect 18799 12484 18803 12540
rect 18739 12480 18803 12484
rect 18819 12540 18883 12544
rect 18819 12484 18823 12540
rect 18823 12484 18879 12540
rect 18879 12484 18883 12540
rect 18819 12480 18883 12484
rect 18899 12540 18963 12544
rect 18899 12484 18903 12540
rect 18903 12484 18959 12540
rect 18959 12484 18963 12540
rect 18899 12480 18963 12484
rect 25742 12540 25806 12544
rect 25742 12484 25746 12540
rect 25746 12484 25802 12540
rect 25802 12484 25806 12540
rect 25742 12480 25806 12484
rect 25822 12540 25886 12544
rect 25822 12484 25826 12540
rect 25826 12484 25882 12540
rect 25882 12484 25886 12540
rect 25822 12480 25886 12484
rect 25902 12540 25966 12544
rect 25902 12484 25906 12540
rect 25906 12484 25962 12540
rect 25962 12484 25966 12540
rect 25902 12480 25966 12484
rect 25982 12540 26046 12544
rect 25982 12484 25986 12540
rect 25986 12484 26042 12540
rect 26042 12484 26046 12540
rect 25982 12480 26046 12484
rect 8034 11996 8098 12000
rect 8034 11940 8038 11996
rect 8038 11940 8094 11996
rect 8094 11940 8098 11996
rect 8034 11936 8098 11940
rect 8114 11996 8178 12000
rect 8114 11940 8118 11996
rect 8118 11940 8174 11996
rect 8174 11940 8178 11996
rect 8114 11936 8178 11940
rect 8194 11996 8258 12000
rect 8194 11940 8198 11996
rect 8198 11940 8254 11996
rect 8254 11940 8258 11996
rect 8194 11936 8258 11940
rect 8274 11996 8338 12000
rect 8274 11940 8278 11996
rect 8278 11940 8334 11996
rect 8334 11940 8338 11996
rect 8274 11936 8338 11940
rect 15117 11996 15181 12000
rect 15117 11940 15121 11996
rect 15121 11940 15177 11996
rect 15177 11940 15181 11996
rect 15117 11936 15181 11940
rect 15197 11996 15261 12000
rect 15197 11940 15201 11996
rect 15201 11940 15257 11996
rect 15257 11940 15261 11996
rect 15197 11936 15261 11940
rect 15277 11996 15341 12000
rect 15277 11940 15281 11996
rect 15281 11940 15337 11996
rect 15337 11940 15341 11996
rect 15277 11936 15341 11940
rect 15357 11996 15421 12000
rect 15357 11940 15361 11996
rect 15361 11940 15417 11996
rect 15417 11940 15421 11996
rect 15357 11936 15421 11940
rect 22200 11996 22264 12000
rect 22200 11940 22204 11996
rect 22204 11940 22260 11996
rect 22260 11940 22264 11996
rect 22200 11936 22264 11940
rect 22280 11996 22344 12000
rect 22280 11940 22284 11996
rect 22284 11940 22340 11996
rect 22340 11940 22344 11996
rect 22280 11936 22344 11940
rect 22360 11996 22424 12000
rect 22360 11940 22364 11996
rect 22364 11940 22420 11996
rect 22420 11940 22424 11996
rect 22360 11936 22424 11940
rect 22440 11996 22504 12000
rect 22440 11940 22444 11996
rect 22444 11940 22500 11996
rect 22500 11940 22504 11996
rect 22440 11936 22504 11940
rect 29283 11996 29347 12000
rect 29283 11940 29287 11996
rect 29287 11940 29343 11996
rect 29343 11940 29347 11996
rect 29283 11936 29347 11940
rect 29363 11996 29427 12000
rect 29363 11940 29367 11996
rect 29367 11940 29423 11996
rect 29423 11940 29427 11996
rect 29363 11936 29427 11940
rect 29443 11996 29507 12000
rect 29443 11940 29447 11996
rect 29447 11940 29503 11996
rect 29503 11940 29507 11996
rect 29443 11936 29507 11940
rect 29523 11996 29587 12000
rect 29523 11940 29527 11996
rect 29527 11940 29583 11996
rect 29583 11940 29587 11996
rect 29523 11936 29587 11940
rect 27660 11732 27724 11796
rect 4493 11452 4557 11456
rect 4493 11396 4497 11452
rect 4497 11396 4553 11452
rect 4553 11396 4557 11452
rect 4493 11392 4557 11396
rect 4573 11452 4637 11456
rect 4573 11396 4577 11452
rect 4577 11396 4633 11452
rect 4633 11396 4637 11452
rect 4573 11392 4637 11396
rect 4653 11452 4717 11456
rect 4653 11396 4657 11452
rect 4657 11396 4713 11452
rect 4713 11396 4717 11452
rect 4653 11392 4717 11396
rect 4733 11452 4797 11456
rect 4733 11396 4737 11452
rect 4737 11396 4793 11452
rect 4793 11396 4797 11452
rect 4733 11392 4797 11396
rect 11576 11452 11640 11456
rect 11576 11396 11580 11452
rect 11580 11396 11636 11452
rect 11636 11396 11640 11452
rect 11576 11392 11640 11396
rect 11656 11452 11720 11456
rect 11656 11396 11660 11452
rect 11660 11396 11716 11452
rect 11716 11396 11720 11452
rect 11656 11392 11720 11396
rect 11736 11452 11800 11456
rect 11736 11396 11740 11452
rect 11740 11396 11796 11452
rect 11796 11396 11800 11452
rect 11736 11392 11800 11396
rect 11816 11452 11880 11456
rect 11816 11396 11820 11452
rect 11820 11396 11876 11452
rect 11876 11396 11880 11452
rect 11816 11392 11880 11396
rect 18659 11452 18723 11456
rect 18659 11396 18663 11452
rect 18663 11396 18719 11452
rect 18719 11396 18723 11452
rect 18659 11392 18723 11396
rect 18739 11452 18803 11456
rect 18739 11396 18743 11452
rect 18743 11396 18799 11452
rect 18799 11396 18803 11452
rect 18739 11392 18803 11396
rect 18819 11452 18883 11456
rect 18819 11396 18823 11452
rect 18823 11396 18879 11452
rect 18879 11396 18883 11452
rect 18819 11392 18883 11396
rect 18899 11452 18963 11456
rect 18899 11396 18903 11452
rect 18903 11396 18959 11452
rect 18959 11396 18963 11452
rect 18899 11392 18963 11396
rect 25742 11452 25806 11456
rect 25742 11396 25746 11452
rect 25746 11396 25802 11452
rect 25802 11396 25806 11452
rect 25742 11392 25806 11396
rect 25822 11452 25886 11456
rect 25822 11396 25826 11452
rect 25826 11396 25882 11452
rect 25882 11396 25886 11452
rect 25822 11392 25886 11396
rect 25902 11452 25966 11456
rect 25902 11396 25906 11452
rect 25906 11396 25962 11452
rect 25962 11396 25966 11452
rect 25902 11392 25966 11396
rect 25982 11452 26046 11456
rect 25982 11396 25986 11452
rect 25986 11396 26042 11452
rect 26042 11396 26046 11452
rect 25982 11392 26046 11396
rect 8034 10908 8098 10912
rect 8034 10852 8038 10908
rect 8038 10852 8094 10908
rect 8094 10852 8098 10908
rect 8034 10848 8098 10852
rect 8114 10908 8178 10912
rect 8114 10852 8118 10908
rect 8118 10852 8174 10908
rect 8174 10852 8178 10908
rect 8114 10848 8178 10852
rect 8194 10908 8258 10912
rect 8194 10852 8198 10908
rect 8198 10852 8254 10908
rect 8254 10852 8258 10908
rect 8194 10848 8258 10852
rect 8274 10908 8338 10912
rect 8274 10852 8278 10908
rect 8278 10852 8334 10908
rect 8334 10852 8338 10908
rect 8274 10848 8338 10852
rect 15117 10908 15181 10912
rect 15117 10852 15121 10908
rect 15121 10852 15177 10908
rect 15177 10852 15181 10908
rect 15117 10848 15181 10852
rect 15197 10908 15261 10912
rect 15197 10852 15201 10908
rect 15201 10852 15257 10908
rect 15257 10852 15261 10908
rect 15197 10848 15261 10852
rect 15277 10908 15341 10912
rect 15277 10852 15281 10908
rect 15281 10852 15337 10908
rect 15337 10852 15341 10908
rect 15277 10848 15341 10852
rect 15357 10908 15421 10912
rect 15357 10852 15361 10908
rect 15361 10852 15417 10908
rect 15417 10852 15421 10908
rect 15357 10848 15421 10852
rect 22200 10908 22264 10912
rect 22200 10852 22204 10908
rect 22204 10852 22260 10908
rect 22260 10852 22264 10908
rect 22200 10848 22264 10852
rect 22280 10908 22344 10912
rect 22280 10852 22284 10908
rect 22284 10852 22340 10908
rect 22340 10852 22344 10908
rect 22280 10848 22344 10852
rect 22360 10908 22424 10912
rect 22360 10852 22364 10908
rect 22364 10852 22420 10908
rect 22420 10852 22424 10908
rect 22360 10848 22424 10852
rect 22440 10908 22504 10912
rect 22440 10852 22444 10908
rect 22444 10852 22500 10908
rect 22500 10852 22504 10908
rect 22440 10848 22504 10852
rect 29283 10908 29347 10912
rect 29283 10852 29287 10908
rect 29287 10852 29343 10908
rect 29343 10852 29347 10908
rect 29283 10848 29347 10852
rect 29363 10908 29427 10912
rect 29363 10852 29367 10908
rect 29367 10852 29423 10908
rect 29423 10852 29427 10908
rect 29363 10848 29427 10852
rect 29443 10908 29507 10912
rect 29443 10852 29447 10908
rect 29447 10852 29503 10908
rect 29503 10852 29507 10908
rect 29443 10848 29507 10852
rect 29523 10908 29587 10912
rect 29523 10852 29527 10908
rect 29527 10852 29583 10908
rect 29583 10852 29587 10908
rect 29523 10848 29587 10852
rect 4493 10364 4557 10368
rect 4493 10308 4497 10364
rect 4497 10308 4553 10364
rect 4553 10308 4557 10364
rect 4493 10304 4557 10308
rect 4573 10364 4637 10368
rect 4573 10308 4577 10364
rect 4577 10308 4633 10364
rect 4633 10308 4637 10364
rect 4573 10304 4637 10308
rect 4653 10364 4717 10368
rect 4653 10308 4657 10364
rect 4657 10308 4713 10364
rect 4713 10308 4717 10364
rect 4653 10304 4717 10308
rect 4733 10364 4797 10368
rect 4733 10308 4737 10364
rect 4737 10308 4793 10364
rect 4793 10308 4797 10364
rect 4733 10304 4797 10308
rect 11576 10364 11640 10368
rect 11576 10308 11580 10364
rect 11580 10308 11636 10364
rect 11636 10308 11640 10364
rect 11576 10304 11640 10308
rect 11656 10364 11720 10368
rect 11656 10308 11660 10364
rect 11660 10308 11716 10364
rect 11716 10308 11720 10364
rect 11656 10304 11720 10308
rect 11736 10364 11800 10368
rect 11736 10308 11740 10364
rect 11740 10308 11796 10364
rect 11796 10308 11800 10364
rect 11736 10304 11800 10308
rect 11816 10364 11880 10368
rect 11816 10308 11820 10364
rect 11820 10308 11876 10364
rect 11876 10308 11880 10364
rect 11816 10304 11880 10308
rect 18659 10364 18723 10368
rect 18659 10308 18663 10364
rect 18663 10308 18719 10364
rect 18719 10308 18723 10364
rect 18659 10304 18723 10308
rect 18739 10364 18803 10368
rect 18739 10308 18743 10364
rect 18743 10308 18799 10364
rect 18799 10308 18803 10364
rect 18739 10304 18803 10308
rect 18819 10364 18883 10368
rect 18819 10308 18823 10364
rect 18823 10308 18879 10364
rect 18879 10308 18883 10364
rect 18819 10304 18883 10308
rect 18899 10364 18963 10368
rect 18899 10308 18903 10364
rect 18903 10308 18959 10364
rect 18959 10308 18963 10364
rect 18899 10304 18963 10308
rect 25742 10364 25806 10368
rect 25742 10308 25746 10364
rect 25746 10308 25802 10364
rect 25802 10308 25806 10364
rect 25742 10304 25806 10308
rect 25822 10364 25886 10368
rect 25822 10308 25826 10364
rect 25826 10308 25882 10364
rect 25882 10308 25886 10364
rect 25822 10304 25886 10308
rect 25902 10364 25966 10368
rect 25902 10308 25906 10364
rect 25906 10308 25962 10364
rect 25962 10308 25966 10364
rect 25902 10304 25966 10308
rect 25982 10364 26046 10368
rect 25982 10308 25986 10364
rect 25986 10308 26042 10364
rect 26042 10308 26046 10364
rect 25982 10304 26046 10308
rect 8034 9820 8098 9824
rect 8034 9764 8038 9820
rect 8038 9764 8094 9820
rect 8094 9764 8098 9820
rect 8034 9760 8098 9764
rect 8114 9820 8178 9824
rect 8114 9764 8118 9820
rect 8118 9764 8174 9820
rect 8174 9764 8178 9820
rect 8114 9760 8178 9764
rect 8194 9820 8258 9824
rect 8194 9764 8198 9820
rect 8198 9764 8254 9820
rect 8254 9764 8258 9820
rect 8194 9760 8258 9764
rect 8274 9820 8338 9824
rect 8274 9764 8278 9820
rect 8278 9764 8334 9820
rect 8334 9764 8338 9820
rect 8274 9760 8338 9764
rect 15117 9820 15181 9824
rect 15117 9764 15121 9820
rect 15121 9764 15177 9820
rect 15177 9764 15181 9820
rect 15117 9760 15181 9764
rect 15197 9820 15261 9824
rect 15197 9764 15201 9820
rect 15201 9764 15257 9820
rect 15257 9764 15261 9820
rect 15197 9760 15261 9764
rect 15277 9820 15341 9824
rect 15277 9764 15281 9820
rect 15281 9764 15337 9820
rect 15337 9764 15341 9820
rect 15277 9760 15341 9764
rect 15357 9820 15421 9824
rect 15357 9764 15361 9820
rect 15361 9764 15417 9820
rect 15417 9764 15421 9820
rect 15357 9760 15421 9764
rect 22200 9820 22264 9824
rect 22200 9764 22204 9820
rect 22204 9764 22260 9820
rect 22260 9764 22264 9820
rect 22200 9760 22264 9764
rect 22280 9820 22344 9824
rect 22280 9764 22284 9820
rect 22284 9764 22340 9820
rect 22340 9764 22344 9820
rect 22280 9760 22344 9764
rect 22360 9820 22424 9824
rect 22360 9764 22364 9820
rect 22364 9764 22420 9820
rect 22420 9764 22424 9820
rect 22360 9760 22424 9764
rect 22440 9820 22504 9824
rect 22440 9764 22444 9820
rect 22444 9764 22500 9820
rect 22500 9764 22504 9820
rect 22440 9760 22504 9764
rect 29283 9820 29347 9824
rect 29283 9764 29287 9820
rect 29287 9764 29343 9820
rect 29343 9764 29347 9820
rect 29283 9760 29347 9764
rect 29363 9820 29427 9824
rect 29363 9764 29367 9820
rect 29367 9764 29423 9820
rect 29423 9764 29427 9820
rect 29363 9760 29427 9764
rect 29443 9820 29507 9824
rect 29443 9764 29447 9820
rect 29447 9764 29503 9820
rect 29503 9764 29507 9820
rect 29443 9760 29507 9764
rect 29523 9820 29587 9824
rect 29523 9764 29527 9820
rect 29527 9764 29583 9820
rect 29583 9764 29587 9820
rect 29523 9760 29587 9764
rect 10180 9420 10244 9484
rect 4493 9276 4557 9280
rect 4493 9220 4497 9276
rect 4497 9220 4553 9276
rect 4553 9220 4557 9276
rect 4493 9216 4557 9220
rect 4573 9276 4637 9280
rect 4573 9220 4577 9276
rect 4577 9220 4633 9276
rect 4633 9220 4637 9276
rect 4573 9216 4637 9220
rect 4653 9276 4717 9280
rect 4653 9220 4657 9276
rect 4657 9220 4713 9276
rect 4713 9220 4717 9276
rect 4653 9216 4717 9220
rect 4733 9276 4797 9280
rect 4733 9220 4737 9276
rect 4737 9220 4793 9276
rect 4793 9220 4797 9276
rect 4733 9216 4797 9220
rect 11576 9276 11640 9280
rect 11576 9220 11580 9276
rect 11580 9220 11636 9276
rect 11636 9220 11640 9276
rect 11576 9216 11640 9220
rect 11656 9276 11720 9280
rect 11656 9220 11660 9276
rect 11660 9220 11716 9276
rect 11716 9220 11720 9276
rect 11656 9216 11720 9220
rect 11736 9276 11800 9280
rect 11736 9220 11740 9276
rect 11740 9220 11796 9276
rect 11796 9220 11800 9276
rect 11736 9216 11800 9220
rect 11816 9276 11880 9280
rect 11816 9220 11820 9276
rect 11820 9220 11876 9276
rect 11876 9220 11880 9276
rect 11816 9216 11880 9220
rect 18659 9276 18723 9280
rect 18659 9220 18663 9276
rect 18663 9220 18719 9276
rect 18719 9220 18723 9276
rect 18659 9216 18723 9220
rect 18739 9276 18803 9280
rect 18739 9220 18743 9276
rect 18743 9220 18799 9276
rect 18799 9220 18803 9276
rect 18739 9216 18803 9220
rect 18819 9276 18883 9280
rect 18819 9220 18823 9276
rect 18823 9220 18879 9276
rect 18879 9220 18883 9276
rect 18819 9216 18883 9220
rect 18899 9276 18963 9280
rect 18899 9220 18903 9276
rect 18903 9220 18959 9276
rect 18959 9220 18963 9276
rect 18899 9216 18963 9220
rect 25742 9276 25806 9280
rect 25742 9220 25746 9276
rect 25746 9220 25802 9276
rect 25802 9220 25806 9276
rect 25742 9216 25806 9220
rect 25822 9276 25886 9280
rect 25822 9220 25826 9276
rect 25826 9220 25882 9276
rect 25882 9220 25886 9276
rect 25822 9216 25886 9220
rect 25902 9276 25966 9280
rect 25902 9220 25906 9276
rect 25906 9220 25962 9276
rect 25962 9220 25966 9276
rect 25902 9216 25966 9220
rect 25982 9276 26046 9280
rect 25982 9220 25986 9276
rect 25986 9220 26042 9276
rect 26042 9220 26046 9276
rect 25982 9216 26046 9220
rect 8034 8732 8098 8736
rect 8034 8676 8038 8732
rect 8038 8676 8094 8732
rect 8094 8676 8098 8732
rect 8034 8672 8098 8676
rect 8114 8732 8178 8736
rect 8114 8676 8118 8732
rect 8118 8676 8174 8732
rect 8174 8676 8178 8732
rect 8114 8672 8178 8676
rect 8194 8732 8258 8736
rect 8194 8676 8198 8732
rect 8198 8676 8254 8732
rect 8254 8676 8258 8732
rect 8194 8672 8258 8676
rect 8274 8732 8338 8736
rect 8274 8676 8278 8732
rect 8278 8676 8334 8732
rect 8334 8676 8338 8732
rect 8274 8672 8338 8676
rect 15117 8732 15181 8736
rect 15117 8676 15121 8732
rect 15121 8676 15177 8732
rect 15177 8676 15181 8732
rect 15117 8672 15181 8676
rect 15197 8732 15261 8736
rect 15197 8676 15201 8732
rect 15201 8676 15257 8732
rect 15257 8676 15261 8732
rect 15197 8672 15261 8676
rect 15277 8732 15341 8736
rect 15277 8676 15281 8732
rect 15281 8676 15337 8732
rect 15337 8676 15341 8732
rect 15277 8672 15341 8676
rect 15357 8732 15421 8736
rect 15357 8676 15361 8732
rect 15361 8676 15417 8732
rect 15417 8676 15421 8732
rect 15357 8672 15421 8676
rect 22200 8732 22264 8736
rect 22200 8676 22204 8732
rect 22204 8676 22260 8732
rect 22260 8676 22264 8732
rect 22200 8672 22264 8676
rect 22280 8732 22344 8736
rect 22280 8676 22284 8732
rect 22284 8676 22340 8732
rect 22340 8676 22344 8732
rect 22280 8672 22344 8676
rect 22360 8732 22424 8736
rect 22360 8676 22364 8732
rect 22364 8676 22420 8732
rect 22420 8676 22424 8732
rect 22360 8672 22424 8676
rect 22440 8732 22504 8736
rect 22440 8676 22444 8732
rect 22444 8676 22500 8732
rect 22500 8676 22504 8732
rect 22440 8672 22504 8676
rect 29283 8732 29347 8736
rect 29283 8676 29287 8732
rect 29287 8676 29343 8732
rect 29343 8676 29347 8732
rect 29283 8672 29347 8676
rect 29363 8732 29427 8736
rect 29363 8676 29367 8732
rect 29367 8676 29423 8732
rect 29423 8676 29427 8732
rect 29363 8672 29427 8676
rect 29443 8732 29507 8736
rect 29443 8676 29447 8732
rect 29447 8676 29503 8732
rect 29503 8676 29507 8732
rect 29443 8672 29507 8676
rect 29523 8732 29587 8736
rect 29523 8676 29527 8732
rect 29527 8676 29583 8732
rect 29583 8676 29587 8732
rect 29523 8672 29587 8676
rect 10548 8256 10612 8260
rect 10548 8200 10562 8256
rect 10562 8200 10612 8256
rect 10548 8196 10612 8200
rect 4493 8188 4557 8192
rect 4493 8132 4497 8188
rect 4497 8132 4553 8188
rect 4553 8132 4557 8188
rect 4493 8128 4557 8132
rect 4573 8188 4637 8192
rect 4573 8132 4577 8188
rect 4577 8132 4633 8188
rect 4633 8132 4637 8188
rect 4573 8128 4637 8132
rect 4653 8188 4717 8192
rect 4653 8132 4657 8188
rect 4657 8132 4713 8188
rect 4713 8132 4717 8188
rect 4653 8128 4717 8132
rect 4733 8188 4797 8192
rect 4733 8132 4737 8188
rect 4737 8132 4793 8188
rect 4793 8132 4797 8188
rect 4733 8128 4797 8132
rect 11576 8188 11640 8192
rect 11576 8132 11580 8188
rect 11580 8132 11636 8188
rect 11636 8132 11640 8188
rect 11576 8128 11640 8132
rect 11656 8188 11720 8192
rect 11656 8132 11660 8188
rect 11660 8132 11716 8188
rect 11716 8132 11720 8188
rect 11656 8128 11720 8132
rect 11736 8188 11800 8192
rect 11736 8132 11740 8188
rect 11740 8132 11796 8188
rect 11796 8132 11800 8188
rect 11736 8128 11800 8132
rect 11816 8188 11880 8192
rect 11816 8132 11820 8188
rect 11820 8132 11876 8188
rect 11876 8132 11880 8188
rect 11816 8128 11880 8132
rect 18659 8188 18723 8192
rect 18659 8132 18663 8188
rect 18663 8132 18719 8188
rect 18719 8132 18723 8188
rect 18659 8128 18723 8132
rect 18739 8188 18803 8192
rect 18739 8132 18743 8188
rect 18743 8132 18799 8188
rect 18799 8132 18803 8188
rect 18739 8128 18803 8132
rect 18819 8188 18883 8192
rect 18819 8132 18823 8188
rect 18823 8132 18879 8188
rect 18879 8132 18883 8188
rect 18819 8128 18883 8132
rect 18899 8188 18963 8192
rect 18899 8132 18903 8188
rect 18903 8132 18959 8188
rect 18959 8132 18963 8188
rect 18899 8128 18963 8132
rect 25742 8188 25806 8192
rect 25742 8132 25746 8188
rect 25746 8132 25802 8188
rect 25802 8132 25806 8188
rect 25742 8128 25806 8132
rect 25822 8188 25886 8192
rect 25822 8132 25826 8188
rect 25826 8132 25882 8188
rect 25882 8132 25886 8188
rect 25822 8128 25886 8132
rect 25902 8188 25966 8192
rect 25902 8132 25906 8188
rect 25906 8132 25962 8188
rect 25962 8132 25966 8188
rect 25902 8128 25966 8132
rect 25982 8188 26046 8192
rect 25982 8132 25986 8188
rect 25986 8132 26042 8188
rect 26042 8132 26046 8188
rect 25982 8128 26046 8132
rect 8034 7644 8098 7648
rect 8034 7588 8038 7644
rect 8038 7588 8094 7644
rect 8094 7588 8098 7644
rect 8034 7584 8098 7588
rect 8114 7644 8178 7648
rect 8114 7588 8118 7644
rect 8118 7588 8174 7644
rect 8174 7588 8178 7644
rect 8114 7584 8178 7588
rect 8194 7644 8258 7648
rect 8194 7588 8198 7644
rect 8198 7588 8254 7644
rect 8254 7588 8258 7644
rect 8194 7584 8258 7588
rect 8274 7644 8338 7648
rect 8274 7588 8278 7644
rect 8278 7588 8334 7644
rect 8334 7588 8338 7644
rect 8274 7584 8338 7588
rect 15117 7644 15181 7648
rect 15117 7588 15121 7644
rect 15121 7588 15177 7644
rect 15177 7588 15181 7644
rect 15117 7584 15181 7588
rect 15197 7644 15261 7648
rect 15197 7588 15201 7644
rect 15201 7588 15257 7644
rect 15257 7588 15261 7644
rect 15197 7584 15261 7588
rect 15277 7644 15341 7648
rect 15277 7588 15281 7644
rect 15281 7588 15337 7644
rect 15337 7588 15341 7644
rect 15277 7584 15341 7588
rect 15357 7644 15421 7648
rect 15357 7588 15361 7644
rect 15361 7588 15417 7644
rect 15417 7588 15421 7644
rect 15357 7584 15421 7588
rect 22200 7644 22264 7648
rect 22200 7588 22204 7644
rect 22204 7588 22260 7644
rect 22260 7588 22264 7644
rect 22200 7584 22264 7588
rect 22280 7644 22344 7648
rect 22280 7588 22284 7644
rect 22284 7588 22340 7644
rect 22340 7588 22344 7644
rect 22280 7584 22344 7588
rect 22360 7644 22424 7648
rect 22360 7588 22364 7644
rect 22364 7588 22420 7644
rect 22420 7588 22424 7644
rect 22360 7584 22424 7588
rect 22440 7644 22504 7648
rect 22440 7588 22444 7644
rect 22444 7588 22500 7644
rect 22500 7588 22504 7644
rect 22440 7584 22504 7588
rect 29283 7644 29347 7648
rect 29283 7588 29287 7644
rect 29287 7588 29343 7644
rect 29343 7588 29347 7644
rect 29283 7584 29347 7588
rect 29363 7644 29427 7648
rect 29363 7588 29367 7644
rect 29367 7588 29423 7644
rect 29423 7588 29427 7644
rect 29363 7584 29427 7588
rect 29443 7644 29507 7648
rect 29443 7588 29447 7644
rect 29447 7588 29503 7644
rect 29503 7588 29507 7644
rect 29443 7584 29507 7588
rect 29523 7644 29587 7648
rect 29523 7588 29527 7644
rect 29527 7588 29583 7644
rect 29583 7588 29587 7644
rect 29523 7584 29587 7588
rect 4493 7100 4557 7104
rect 4493 7044 4497 7100
rect 4497 7044 4553 7100
rect 4553 7044 4557 7100
rect 4493 7040 4557 7044
rect 4573 7100 4637 7104
rect 4573 7044 4577 7100
rect 4577 7044 4633 7100
rect 4633 7044 4637 7100
rect 4573 7040 4637 7044
rect 4653 7100 4717 7104
rect 4653 7044 4657 7100
rect 4657 7044 4713 7100
rect 4713 7044 4717 7100
rect 4653 7040 4717 7044
rect 4733 7100 4797 7104
rect 4733 7044 4737 7100
rect 4737 7044 4793 7100
rect 4793 7044 4797 7100
rect 4733 7040 4797 7044
rect 11576 7100 11640 7104
rect 11576 7044 11580 7100
rect 11580 7044 11636 7100
rect 11636 7044 11640 7100
rect 11576 7040 11640 7044
rect 11656 7100 11720 7104
rect 11656 7044 11660 7100
rect 11660 7044 11716 7100
rect 11716 7044 11720 7100
rect 11656 7040 11720 7044
rect 11736 7100 11800 7104
rect 11736 7044 11740 7100
rect 11740 7044 11796 7100
rect 11796 7044 11800 7100
rect 11736 7040 11800 7044
rect 11816 7100 11880 7104
rect 11816 7044 11820 7100
rect 11820 7044 11876 7100
rect 11876 7044 11880 7100
rect 11816 7040 11880 7044
rect 18659 7100 18723 7104
rect 18659 7044 18663 7100
rect 18663 7044 18719 7100
rect 18719 7044 18723 7100
rect 18659 7040 18723 7044
rect 18739 7100 18803 7104
rect 18739 7044 18743 7100
rect 18743 7044 18799 7100
rect 18799 7044 18803 7100
rect 18739 7040 18803 7044
rect 18819 7100 18883 7104
rect 18819 7044 18823 7100
rect 18823 7044 18879 7100
rect 18879 7044 18883 7100
rect 18819 7040 18883 7044
rect 18899 7100 18963 7104
rect 18899 7044 18903 7100
rect 18903 7044 18959 7100
rect 18959 7044 18963 7100
rect 18899 7040 18963 7044
rect 25742 7100 25806 7104
rect 25742 7044 25746 7100
rect 25746 7044 25802 7100
rect 25802 7044 25806 7100
rect 25742 7040 25806 7044
rect 25822 7100 25886 7104
rect 25822 7044 25826 7100
rect 25826 7044 25882 7100
rect 25882 7044 25886 7100
rect 25822 7040 25886 7044
rect 25902 7100 25966 7104
rect 25902 7044 25906 7100
rect 25906 7044 25962 7100
rect 25962 7044 25966 7100
rect 25902 7040 25966 7044
rect 25982 7100 26046 7104
rect 25982 7044 25986 7100
rect 25986 7044 26042 7100
rect 26042 7044 26046 7100
rect 25982 7040 26046 7044
rect 28764 6700 28828 6764
rect 8034 6556 8098 6560
rect 8034 6500 8038 6556
rect 8038 6500 8094 6556
rect 8094 6500 8098 6556
rect 8034 6496 8098 6500
rect 8114 6556 8178 6560
rect 8114 6500 8118 6556
rect 8118 6500 8174 6556
rect 8174 6500 8178 6556
rect 8114 6496 8178 6500
rect 8194 6556 8258 6560
rect 8194 6500 8198 6556
rect 8198 6500 8254 6556
rect 8254 6500 8258 6556
rect 8194 6496 8258 6500
rect 8274 6556 8338 6560
rect 8274 6500 8278 6556
rect 8278 6500 8334 6556
rect 8334 6500 8338 6556
rect 8274 6496 8338 6500
rect 15117 6556 15181 6560
rect 15117 6500 15121 6556
rect 15121 6500 15177 6556
rect 15177 6500 15181 6556
rect 15117 6496 15181 6500
rect 15197 6556 15261 6560
rect 15197 6500 15201 6556
rect 15201 6500 15257 6556
rect 15257 6500 15261 6556
rect 15197 6496 15261 6500
rect 15277 6556 15341 6560
rect 15277 6500 15281 6556
rect 15281 6500 15337 6556
rect 15337 6500 15341 6556
rect 15277 6496 15341 6500
rect 15357 6556 15421 6560
rect 15357 6500 15361 6556
rect 15361 6500 15417 6556
rect 15417 6500 15421 6556
rect 15357 6496 15421 6500
rect 22200 6556 22264 6560
rect 22200 6500 22204 6556
rect 22204 6500 22260 6556
rect 22260 6500 22264 6556
rect 22200 6496 22264 6500
rect 22280 6556 22344 6560
rect 22280 6500 22284 6556
rect 22284 6500 22340 6556
rect 22340 6500 22344 6556
rect 22280 6496 22344 6500
rect 22360 6556 22424 6560
rect 22360 6500 22364 6556
rect 22364 6500 22420 6556
rect 22420 6500 22424 6556
rect 22360 6496 22424 6500
rect 22440 6556 22504 6560
rect 22440 6500 22444 6556
rect 22444 6500 22500 6556
rect 22500 6500 22504 6556
rect 22440 6496 22504 6500
rect 29283 6556 29347 6560
rect 29283 6500 29287 6556
rect 29287 6500 29343 6556
rect 29343 6500 29347 6556
rect 29283 6496 29347 6500
rect 29363 6556 29427 6560
rect 29363 6500 29367 6556
rect 29367 6500 29423 6556
rect 29423 6500 29427 6556
rect 29363 6496 29427 6500
rect 29443 6556 29507 6560
rect 29443 6500 29447 6556
rect 29447 6500 29503 6556
rect 29503 6500 29507 6556
rect 29443 6496 29507 6500
rect 29523 6556 29587 6560
rect 29523 6500 29527 6556
rect 29527 6500 29583 6556
rect 29583 6500 29587 6556
rect 29523 6496 29587 6500
rect 4493 6012 4557 6016
rect 4493 5956 4497 6012
rect 4497 5956 4553 6012
rect 4553 5956 4557 6012
rect 4493 5952 4557 5956
rect 4573 6012 4637 6016
rect 4573 5956 4577 6012
rect 4577 5956 4633 6012
rect 4633 5956 4637 6012
rect 4573 5952 4637 5956
rect 4653 6012 4717 6016
rect 4653 5956 4657 6012
rect 4657 5956 4713 6012
rect 4713 5956 4717 6012
rect 4653 5952 4717 5956
rect 4733 6012 4797 6016
rect 4733 5956 4737 6012
rect 4737 5956 4793 6012
rect 4793 5956 4797 6012
rect 4733 5952 4797 5956
rect 11576 6012 11640 6016
rect 11576 5956 11580 6012
rect 11580 5956 11636 6012
rect 11636 5956 11640 6012
rect 11576 5952 11640 5956
rect 11656 6012 11720 6016
rect 11656 5956 11660 6012
rect 11660 5956 11716 6012
rect 11716 5956 11720 6012
rect 11656 5952 11720 5956
rect 11736 6012 11800 6016
rect 11736 5956 11740 6012
rect 11740 5956 11796 6012
rect 11796 5956 11800 6012
rect 11736 5952 11800 5956
rect 11816 6012 11880 6016
rect 11816 5956 11820 6012
rect 11820 5956 11876 6012
rect 11876 5956 11880 6012
rect 11816 5952 11880 5956
rect 18659 6012 18723 6016
rect 18659 5956 18663 6012
rect 18663 5956 18719 6012
rect 18719 5956 18723 6012
rect 18659 5952 18723 5956
rect 18739 6012 18803 6016
rect 18739 5956 18743 6012
rect 18743 5956 18799 6012
rect 18799 5956 18803 6012
rect 18739 5952 18803 5956
rect 18819 6012 18883 6016
rect 18819 5956 18823 6012
rect 18823 5956 18879 6012
rect 18879 5956 18883 6012
rect 18819 5952 18883 5956
rect 18899 6012 18963 6016
rect 18899 5956 18903 6012
rect 18903 5956 18959 6012
rect 18959 5956 18963 6012
rect 18899 5952 18963 5956
rect 25742 6012 25806 6016
rect 25742 5956 25746 6012
rect 25746 5956 25802 6012
rect 25802 5956 25806 6012
rect 25742 5952 25806 5956
rect 25822 6012 25886 6016
rect 25822 5956 25826 6012
rect 25826 5956 25882 6012
rect 25882 5956 25886 6012
rect 25822 5952 25886 5956
rect 25902 6012 25966 6016
rect 25902 5956 25906 6012
rect 25906 5956 25962 6012
rect 25962 5956 25966 6012
rect 25902 5952 25966 5956
rect 25982 6012 26046 6016
rect 25982 5956 25986 6012
rect 25986 5956 26042 6012
rect 26042 5956 26046 6012
rect 25982 5952 26046 5956
rect 24348 5536 24412 5540
rect 24348 5480 24362 5536
rect 24362 5480 24412 5536
rect 24348 5476 24412 5480
rect 8034 5468 8098 5472
rect 8034 5412 8038 5468
rect 8038 5412 8094 5468
rect 8094 5412 8098 5468
rect 8034 5408 8098 5412
rect 8114 5468 8178 5472
rect 8114 5412 8118 5468
rect 8118 5412 8174 5468
rect 8174 5412 8178 5468
rect 8114 5408 8178 5412
rect 8194 5468 8258 5472
rect 8194 5412 8198 5468
rect 8198 5412 8254 5468
rect 8254 5412 8258 5468
rect 8194 5408 8258 5412
rect 8274 5468 8338 5472
rect 8274 5412 8278 5468
rect 8278 5412 8334 5468
rect 8334 5412 8338 5468
rect 8274 5408 8338 5412
rect 15117 5468 15181 5472
rect 15117 5412 15121 5468
rect 15121 5412 15177 5468
rect 15177 5412 15181 5468
rect 15117 5408 15181 5412
rect 15197 5468 15261 5472
rect 15197 5412 15201 5468
rect 15201 5412 15257 5468
rect 15257 5412 15261 5468
rect 15197 5408 15261 5412
rect 15277 5468 15341 5472
rect 15277 5412 15281 5468
rect 15281 5412 15337 5468
rect 15337 5412 15341 5468
rect 15277 5408 15341 5412
rect 15357 5468 15421 5472
rect 15357 5412 15361 5468
rect 15361 5412 15417 5468
rect 15417 5412 15421 5468
rect 15357 5408 15421 5412
rect 22200 5468 22264 5472
rect 22200 5412 22204 5468
rect 22204 5412 22260 5468
rect 22260 5412 22264 5468
rect 22200 5408 22264 5412
rect 22280 5468 22344 5472
rect 22280 5412 22284 5468
rect 22284 5412 22340 5468
rect 22340 5412 22344 5468
rect 22280 5408 22344 5412
rect 22360 5468 22424 5472
rect 22360 5412 22364 5468
rect 22364 5412 22420 5468
rect 22420 5412 22424 5468
rect 22360 5408 22424 5412
rect 22440 5468 22504 5472
rect 22440 5412 22444 5468
rect 22444 5412 22500 5468
rect 22500 5412 22504 5468
rect 22440 5408 22504 5412
rect 29283 5468 29347 5472
rect 29283 5412 29287 5468
rect 29287 5412 29343 5468
rect 29343 5412 29347 5468
rect 29283 5408 29347 5412
rect 29363 5468 29427 5472
rect 29363 5412 29367 5468
rect 29367 5412 29423 5468
rect 29423 5412 29427 5468
rect 29363 5408 29427 5412
rect 29443 5468 29507 5472
rect 29443 5412 29447 5468
rect 29447 5412 29503 5468
rect 29503 5412 29507 5468
rect 29443 5408 29507 5412
rect 29523 5468 29587 5472
rect 29523 5412 29527 5468
rect 29527 5412 29583 5468
rect 29583 5412 29587 5468
rect 29523 5408 29587 5412
rect 4493 4924 4557 4928
rect 4493 4868 4497 4924
rect 4497 4868 4553 4924
rect 4553 4868 4557 4924
rect 4493 4864 4557 4868
rect 4573 4924 4637 4928
rect 4573 4868 4577 4924
rect 4577 4868 4633 4924
rect 4633 4868 4637 4924
rect 4573 4864 4637 4868
rect 4653 4924 4717 4928
rect 4653 4868 4657 4924
rect 4657 4868 4713 4924
rect 4713 4868 4717 4924
rect 4653 4864 4717 4868
rect 4733 4924 4797 4928
rect 4733 4868 4737 4924
rect 4737 4868 4793 4924
rect 4793 4868 4797 4924
rect 4733 4864 4797 4868
rect 11576 4924 11640 4928
rect 11576 4868 11580 4924
rect 11580 4868 11636 4924
rect 11636 4868 11640 4924
rect 11576 4864 11640 4868
rect 11656 4924 11720 4928
rect 11656 4868 11660 4924
rect 11660 4868 11716 4924
rect 11716 4868 11720 4924
rect 11656 4864 11720 4868
rect 11736 4924 11800 4928
rect 11736 4868 11740 4924
rect 11740 4868 11796 4924
rect 11796 4868 11800 4924
rect 11736 4864 11800 4868
rect 11816 4924 11880 4928
rect 11816 4868 11820 4924
rect 11820 4868 11876 4924
rect 11876 4868 11880 4924
rect 11816 4864 11880 4868
rect 18659 4924 18723 4928
rect 18659 4868 18663 4924
rect 18663 4868 18719 4924
rect 18719 4868 18723 4924
rect 18659 4864 18723 4868
rect 18739 4924 18803 4928
rect 18739 4868 18743 4924
rect 18743 4868 18799 4924
rect 18799 4868 18803 4924
rect 18739 4864 18803 4868
rect 18819 4924 18883 4928
rect 18819 4868 18823 4924
rect 18823 4868 18879 4924
rect 18879 4868 18883 4924
rect 18819 4864 18883 4868
rect 18899 4924 18963 4928
rect 18899 4868 18903 4924
rect 18903 4868 18959 4924
rect 18959 4868 18963 4924
rect 18899 4864 18963 4868
rect 25742 4924 25806 4928
rect 25742 4868 25746 4924
rect 25746 4868 25802 4924
rect 25802 4868 25806 4924
rect 25742 4864 25806 4868
rect 25822 4924 25886 4928
rect 25822 4868 25826 4924
rect 25826 4868 25882 4924
rect 25882 4868 25886 4924
rect 25822 4864 25886 4868
rect 25902 4924 25966 4928
rect 25902 4868 25906 4924
rect 25906 4868 25962 4924
rect 25962 4868 25966 4924
rect 25902 4864 25966 4868
rect 25982 4924 26046 4928
rect 25982 4868 25986 4924
rect 25986 4868 26042 4924
rect 26042 4868 26046 4924
rect 25982 4864 26046 4868
rect 8034 4380 8098 4384
rect 8034 4324 8038 4380
rect 8038 4324 8094 4380
rect 8094 4324 8098 4380
rect 8034 4320 8098 4324
rect 8114 4380 8178 4384
rect 8114 4324 8118 4380
rect 8118 4324 8174 4380
rect 8174 4324 8178 4380
rect 8114 4320 8178 4324
rect 8194 4380 8258 4384
rect 8194 4324 8198 4380
rect 8198 4324 8254 4380
rect 8254 4324 8258 4380
rect 8194 4320 8258 4324
rect 8274 4380 8338 4384
rect 8274 4324 8278 4380
rect 8278 4324 8334 4380
rect 8334 4324 8338 4380
rect 8274 4320 8338 4324
rect 15117 4380 15181 4384
rect 15117 4324 15121 4380
rect 15121 4324 15177 4380
rect 15177 4324 15181 4380
rect 15117 4320 15181 4324
rect 15197 4380 15261 4384
rect 15197 4324 15201 4380
rect 15201 4324 15257 4380
rect 15257 4324 15261 4380
rect 15197 4320 15261 4324
rect 15277 4380 15341 4384
rect 15277 4324 15281 4380
rect 15281 4324 15337 4380
rect 15337 4324 15341 4380
rect 15277 4320 15341 4324
rect 15357 4380 15421 4384
rect 15357 4324 15361 4380
rect 15361 4324 15417 4380
rect 15417 4324 15421 4380
rect 15357 4320 15421 4324
rect 22200 4380 22264 4384
rect 22200 4324 22204 4380
rect 22204 4324 22260 4380
rect 22260 4324 22264 4380
rect 22200 4320 22264 4324
rect 22280 4380 22344 4384
rect 22280 4324 22284 4380
rect 22284 4324 22340 4380
rect 22340 4324 22344 4380
rect 22280 4320 22344 4324
rect 22360 4380 22424 4384
rect 22360 4324 22364 4380
rect 22364 4324 22420 4380
rect 22420 4324 22424 4380
rect 22360 4320 22424 4324
rect 22440 4380 22504 4384
rect 22440 4324 22444 4380
rect 22444 4324 22500 4380
rect 22500 4324 22504 4380
rect 22440 4320 22504 4324
rect 29283 4380 29347 4384
rect 29283 4324 29287 4380
rect 29287 4324 29343 4380
rect 29343 4324 29347 4380
rect 29283 4320 29347 4324
rect 29363 4380 29427 4384
rect 29363 4324 29367 4380
rect 29367 4324 29423 4380
rect 29423 4324 29427 4380
rect 29363 4320 29427 4324
rect 29443 4380 29507 4384
rect 29443 4324 29447 4380
rect 29447 4324 29503 4380
rect 29503 4324 29507 4380
rect 29443 4320 29507 4324
rect 29523 4380 29587 4384
rect 29523 4324 29527 4380
rect 29527 4324 29583 4380
rect 29583 4324 29587 4380
rect 29523 4320 29587 4324
rect 4493 3836 4557 3840
rect 4493 3780 4497 3836
rect 4497 3780 4553 3836
rect 4553 3780 4557 3836
rect 4493 3776 4557 3780
rect 4573 3836 4637 3840
rect 4573 3780 4577 3836
rect 4577 3780 4633 3836
rect 4633 3780 4637 3836
rect 4573 3776 4637 3780
rect 4653 3836 4717 3840
rect 4653 3780 4657 3836
rect 4657 3780 4713 3836
rect 4713 3780 4717 3836
rect 4653 3776 4717 3780
rect 4733 3836 4797 3840
rect 4733 3780 4737 3836
rect 4737 3780 4793 3836
rect 4793 3780 4797 3836
rect 4733 3776 4797 3780
rect 11576 3836 11640 3840
rect 11576 3780 11580 3836
rect 11580 3780 11636 3836
rect 11636 3780 11640 3836
rect 11576 3776 11640 3780
rect 11656 3836 11720 3840
rect 11656 3780 11660 3836
rect 11660 3780 11716 3836
rect 11716 3780 11720 3836
rect 11656 3776 11720 3780
rect 11736 3836 11800 3840
rect 11736 3780 11740 3836
rect 11740 3780 11796 3836
rect 11796 3780 11800 3836
rect 11736 3776 11800 3780
rect 11816 3836 11880 3840
rect 11816 3780 11820 3836
rect 11820 3780 11876 3836
rect 11876 3780 11880 3836
rect 11816 3776 11880 3780
rect 18659 3836 18723 3840
rect 18659 3780 18663 3836
rect 18663 3780 18719 3836
rect 18719 3780 18723 3836
rect 18659 3776 18723 3780
rect 18739 3836 18803 3840
rect 18739 3780 18743 3836
rect 18743 3780 18799 3836
rect 18799 3780 18803 3836
rect 18739 3776 18803 3780
rect 18819 3836 18883 3840
rect 18819 3780 18823 3836
rect 18823 3780 18879 3836
rect 18879 3780 18883 3836
rect 18819 3776 18883 3780
rect 18899 3836 18963 3840
rect 18899 3780 18903 3836
rect 18903 3780 18959 3836
rect 18959 3780 18963 3836
rect 18899 3776 18963 3780
rect 25742 3836 25806 3840
rect 25742 3780 25746 3836
rect 25746 3780 25802 3836
rect 25802 3780 25806 3836
rect 25742 3776 25806 3780
rect 25822 3836 25886 3840
rect 25822 3780 25826 3836
rect 25826 3780 25882 3836
rect 25882 3780 25886 3836
rect 25822 3776 25886 3780
rect 25902 3836 25966 3840
rect 25902 3780 25906 3836
rect 25906 3780 25962 3836
rect 25962 3780 25966 3836
rect 25902 3776 25966 3780
rect 25982 3836 26046 3840
rect 25982 3780 25986 3836
rect 25986 3780 26042 3836
rect 26042 3780 26046 3836
rect 25982 3776 26046 3780
rect 8034 3292 8098 3296
rect 8034 3236 8038 3292
rect 8038 3236 8094 3292
rect 8094 3236 8098 3292
rect 8034 3232 8098 3236
rect 8114 3292 8178 3296
rect 8114 3236 8118 3292
rect 8118 3236 8174 3292
rect 8174 3236 8178 3292
rect 8114 3232 8178 3236
rect 8194 3292 8258 3296
rect 8194 3236 8198 3292
rect 8198 3236 8254 3292
rect 8254 3236 8258 3292
rect 8194 3232 8258 3236
rect 8274 3292 8338 3296
rect 8274 3236 8278 3292
rect 8278 3236 8334 3292
rect 8334 3236 8338 3292
rect 8274 3232 8338 3236
rect 15117 3292 15181 3296
rect 15117 3236 15121 3292
rect 15121 3236 15177 3292
rect 15177 3236 15181 3292
rect 15117 3232 15181 3236
rect 15197 3292 15261 3296
rect 15197 3236 15201 3292
rect 15201 3236 15257 3292
rect 15257 3236 15261 3292
rect 15197 3232 15261 3236
rect 15277 3292 15341 3296
rect 15277 3236 15281 3292
rect 15281 3236 15337 3292
rect 15337 3236 15341 3292
rect 15277 3232 15341 3236
rect 15357 3292 15421 3296
rect 15357 3236 15361 3292
rect 15361 3236 15417 3292
rect 15417 3236 15421 3292
rect 15357 3232 15421 3236
rect 22200 3292 22264 3296
rect 22200 3236 22204 3292
rect 22204 3236 22260 3292
rect 22260 3236 22264 3292
rect 22200 3232 22264 3236
rect 22280 3292 22344 3296
rect 22280 3236 22284 3292
rect 22284 3236 22340 3292
rect 22340 3236 22344 3292
rect 22280 3232 22344 3236
rect 22360 3292 22424 3296
rect 22360 3236 22364 3292
rect 22364 3236 22420 3292
rect 22420 3236 22424 3292
rect 22360 3232 22424 3236
rect 22440 3292 22504 3296
rect 22440 3236 22444 3292
rect 22444 3236 22500 3292
rect 22500 3236 22504 3292
rect 22440 3232 22504 3236
rect 29283 3292 29347 3296
rect 29283 3236 29287 3292
rect 29287 3236 29343 3292
rect 29343 3236 29347 3292
rect 29283 3232 29347 3236
rect 29363 3292 29427 3296
rect 29363 3236 29367 3292
rect 29367 3236 29423 3292
rect 29423 3236 29427 3292
rect 29363 3232 29427 3236
rect 29443 3292 29507 3296
rect 29443 3236 29447 3292
rect 29447 3236 29503 3292
rect 29503 3236 29507 3292
rect 29443 3232 29507 3236
rect 29523 3292 29587 3296
rect 29523 3236 29527 3292
rect 29527 3236 29583 3292
rect 29583 3236 29587 3292
rect 29523 3232 29587 3236
rect 4493 2748 4557 2752
rect 4493 2692 4497 2748
rect 4497 2692 4553 2748
rect 4553 2692 4557 2748
rect 4493 2688 4557 2692
rect 4573 2748 4637 2752
rect 4573 2692 4577 2748
rect 4577 2692 4633 2748
rect 4633 2692 4637 2748
rect 4573 2688 4637 2692
rect 4653 2748 4717 2752
rect 4653 2692 4657 2748
rect 4657 2692 4713 2748
rect 4713 2692 4717 2748
rect 4653 2688 4717 2692
rect 4733 2748 4797 2752
rect 4733 2692 4737 2748
rect 4737 2692 4793 2748
rect 4793 2692 4797 2748
rect 4733 2688 4797 2692
rect 11576 2748 11640 2752
rect 11576 2692 11580 2748
rect 11580 2692 11636 2748
rect 11636 2692 11640 2748
rect 11576 2688 11640 2692
rect 11656 2748 11720 2752
rect 11656 2692 11660 2748
rect 11660 2692 11716 2748
rect 11716 2692 11720 2748
rect 11656 2688 11720 2692
rect 11736 2748 11800 2752
rect 11736 2692 11740 2748
rect 11740 2692 11796 2748
rect 11796 2692 11800 2748
rect 11736 2688 11800 2692
rect 11816 2748 11880 2752
rect 11816 2692 11820 2748
rect 11820 2692 11876 2748
rect 11876 2692 11880 2748
rect 11816 2688 11880 2692
rect 18659 2748 18723 2752
rect 18659 2692 18663 2748
rect 18663 2692 18719 2748
rect 18719 2692 18723 2748
rect 18659 2688 18723 2692
rect 18739 2748 18803 2752
rect 18739 2692 18743 2748
rect 18743 2692 18799 2748
rect 18799 2692 18803 2748
rect 18739 2688 18803 2692
rect 18819 2748 18883 2752
rect 18819 2692 18823 2748
rect 18823 2692 18879 2748
rect 18879 2692 18883 2748
rect 18819 2688 18883 2692
rect 18899 2748 18963 2752
rect 18899 2692 18903 2748
rect 18903 2692 18959 2748
rect 18959 2692 18963 2748
rect 18899 2688 18963 2692
rect 25742 2748 25806 2752
rect 25742 2692 25746 2748
rect 25746 2692 25802 2748
rect 25802 2692 25806 2748
rect 25742 2688 25806 2692
rect 25822 2748 25886 2752
rect 25822 2692 25826 2748
rect 25826 2692 25882 2748
rect 25882 2692 25886 2748
rect 25822 2688 25886 2692
rect 25902 2748 25966 2752
rect 25902 2692 25906 2748
rect 25906 2692 25962 2748
rect 25962 2692 25966 2748
rect 25902 2688 25966 2692
rect 25982 2748 26046 2752
rect 25982 2692 25986 2748
rect 25986 2692 26042 2748
rect 26042 2692 26046 2748
rect 25982 2688 26046 2692
rect 8034 2204 8098 2208
rect 8034 2148 8038 2204
rect 8038 2148 8094 2204
rect 8094 2148 8098 2204
rect 8034 2144 8098 2148
rect 8114 2204 8178 2208
rect 8114 2148 8118 2204
rect 8118 2148 8174 2204
rect 8174 2148 8178 2204
rect 8114 2144 8178 2148
rect 8194 2204 8258 2208
rect 8194 2148 8198 2204
rect 8198 2148 8254 2204
rect 8254 2148 8258 2204
rect 8194 2144 8258 2148
rect 8274 2204 8338 2208
rect 8274 2148 8278 2204
rect 8278 2148 8334 2204
rect 8334 2148 8338 2204
rect 8274 2144 8338 2148
rect 15117 2204 15181 2208
rect 15117 2148 15121 2204
rect 15121 2148 15177 2204
rect 15177 2148 15181 2204
rect 15117 2144 15181 2148
rect 15197 2204 15261 2208
rect 15197 2148 15201 2204
rect 15201 2148 15257 2204
rect 15257 2148 15261 2204
rect 15197 2144 15261 2148
rect 15277 2204 15341 2208
rect 15277 2148 15281 2204
rect 15281 2148 15337 2204
rect 15337 2148 15341 2204
rect 15277 2144 15341 2148
rect 15357 2204 15421 2208
rect 15357 2148 15361 2204
rect 15361 2148 15417 2204
rect 15417 2148 15421 2204
rect 15357 2144 15421 2148
rect 22200 2204 22264 2208
rect 22200 2148 22204 2204
rect 22204 2148 22260 2204
rect 22260 2148 22264 2204
rect 22200 2144 22264 2148
rect 22280 2204 22344 2208
rect 22280 2148 22284 2204
rect 22284 2148 22340 2204
rect 22340 2148 22344 2204
rect 22280 2144 22344 2148
rect 22360 2204 22424 2208
rect 22360 2148 22364 2204
rect 22364 2148 22420 2204
rect 22420 2148 22424 2204
rect 22360 2144 22424 2148
rect 22440 2204 22504 2208
rect 22440 2148 22444 2204
rect 22444 2148 22500 2204
rect 22500 2148 22504 2204
rect 22440 2144 22504 2148
rect 29283 2204 29347 2208
rect 29283 2148 29287 2204
rect 29287 2148 29343 2204
rect 29343 2148 29347 2204
rect 29283 2144 29347 2148
rect 29363 2204 29427 2208
rect 29363 2148 29367 2204
rect 29367 2148 29423 2204
rect 29423 2148 29427 2204
rect 29363 2144 29427 2148
rect 29443 2204 29507 2208
rect 29443 2148 29447 2204
rect 29447 2148 29503 2204
rect 29503 2148 29507 2204
rect 29443 2144 29507 2148
rect 29523 2204 29587 2208
rect 29523 2148 29527 2204
rect 29527 2148 29583 2204
rect 29583 2148 29587 2204
rect 29523 2144 29587 2148
<< metal4 >>
rect 4485 29952 4805 30512
rect 4485 29888 4493 29952
rect 4557 29888 4573 29952
rect 4637 29888 4653 29952
rect 4717 29888 4733 29952
rect 4797 29888 4805 29952
rect 4485 28864 4805 29888
rect 4485 28800 4493 28864
rect 4557 28800 4573 28864
rect 4637 28800 4653 28864
rect 4717 28800 4733 28864
rect 4797 28800 4805 28864
rect 4485 27776 4805 28800
rect 4485 27712 4493 27776
rect 4557 27712 4573 27776
rect 4637 27712 4653 27776
rect 4717 27712 4733 27776
rect 4797 27712 4805 27776
rect 4485 26688 4805 27712
rect 4485 26624 4493 26688
rect 4557 26624 4573 26688
rect 4637 26624 4653 26688
rect 4717 26624 4733 26688
rect 4797 26624 4805 26688
rect 4485 25600 4805 26624
rect 4485 25536 4493 25600
rect 4557 25536 4573 25600
rect 4637 25536 4653 25600
rect 4717 25536 4733 25600
rect 4797 25536 4805 25600
rect 4485 24512 4805 25536
rect 4485 24448 4493 24512
rect 4557 24448 4573 24512
rect 4637 24448 4653 24512
rect 4717 24448 4733 24512
rect 4797 24448 4805 24512
rect 4485 23424 4805 24448
rect 4485 23360 4493 23424
rect 4557 23360 4573 23424
rect 4637 23360 4653 23424
rect 4717 23360 4733 23424
rect 4797 23360 4805 23424
rect 4485 22336 4805 23360
rect 4485 22272 4493 22336
rect 4557 22272 4573 22336
rect 4637 22272 4653 22336
rect 4717 22272 4733 22336
rect 4797 22272 4805 22336
rect 4485 21248 4805 22272
rect 4485 21184 4493 21248
rect 4557 21184 4573 21248
rect 4637 21184 4653 21248
rect 4717 21184 4733 21248
rect 4797 21184 4805 21248
rect 4485 20160 4805 21184
rect 4485 20096 4493 20160
rect 4557 20096 4573 20160
rect 4637 20096 4653 20160
rect 4717 20096 4733 20160
rect 4797 20096 4805 20160
rect 4485 19072 4805 20096
rect 4485 19008 4493 19072
rect 4557 19008 4573 19072
rect 4637 19008 4653 19072
rect 4717 19008 4733 19072
rect 4797 19008 4805 19072
rect 4485 17984 4805 19008
rect 4485 17920 4493 17984
rect 4557 17920 4573 17984
rect 4637 17920 4653 17984
rect 4717 17920 4733 17984
rect 4797 17920 4805 17984
rect 4485 16896 4805 17920
rect 4485 16832 4493 16896
rect 4557 16832 4573 16896
rect 4637 16832 4653 16896
rect 4717 16832 4733 16896
rect 4797 16832 4805 16896
rect 4485 15808 4805 16832
rect 4485 15744 4493 15808
rect 4557 15744 4573 15808
rect 4637 15744 4653 15808
rect 4717 15744 4733 15808
rect 4797 15744 4805 15808
rect 4485 14720 4805 15744
rect 4485 14656 4493 14720
rect 4557 14656 4573 14720
rect 4637 14656 4653 14720
rect 4717 14656 4733 14720
rect 4797 14656 4805 14720
rect 4485 13632 4805 14656
rect 4485 13568 4493 13632
rect 4557 13568 4573 13632
rect 4637 13568 4653 13632
rect 4717 13568 4733 13632
rect 4797 13568 4805 13632
rect 4485 12544 4805 13568
rect 4485 12480 4493 12544
rect 4557 12480 4573 12544
rect 4637 12480 4653 12544
rect 4717 12480 4733 12544
rect 4797 12480 4805 12544
rect 4485 11456 4805 12480
rect 4485 11392 4493 11456
rect 4557 11392 4573 11456
rect 4637 11392 4653 11456
rect 4717 11392 4733 11456
rect 4797 11392 4805 11456
rect 4485 10368 4805 11392
rect 4485 10304 4493 10368
rect 4557 10304 4573 10368
rect 4637 10304 4653 10368
rect 4717 10304 4733 10368
rect 4797 10304 4805 10368
rect 4485 9280 4805 10304
rect 4485 9216 4493 9280
rect 4557 9216 4573 9280
rect 4637 9216 4653 9280
rect 4717 9216 4733 9280
rect 4797 9216 4805 9280
rect 4485 8192 4805 9216
rect 4485 8128 4493 8192
rect 4557 8128 4573 8192
rect 4637 8128 4653 8192
rect 4717 8128 4733 8192
rect 4797 8128 4805 8192
rect 4485 7104 4805 8128
rect 4485 7040 4493 7104
rect 4557 7040 4573 7104
rect 4637 7040 4653 7104
rect 4717 7040 4733 7104
rect 4797 7040 4805 7104
rect 4485 6016 4805 7040
rect 4485 5952 4493 6016
rect 4557 5952 4573 6016
rect 4637 5952 4653 6016
rect 4717 5952 4733 6016
rect 4797 5952 4805 6016
rect 4485 4928 4805 5952
rect 4485 4864 4493 4928
rect 4557 4864 4573 4928
rect 4637 4864 4653 4928
rect 4717 4864 4733 4928
rect 4797 4864 4805 4928
rect 4485 3840 4805 4864
rect 4485 3776 4493 3840
rect 4557 3776 4573 3840
rect 4637 3776 4653 3840
rect 4717 3776 4733 3840
rect 4797 3776 4805 3840
rect 4485 2752 4805 3776
rect 4485 2688 4493 2752
rect 4557 2688 4573 2752
rect 4637 2688 4653 2752
rect 4717 2688 4733 2752
rect 4797 2688 4805 2752
rect 4485 2128 4805 2688
rect 8026 30496 8346 30512
rect 8026 30432 8034 30496
rect 8098 30432 8114 30496
rect 8178 30432 8194 30496
rect 8258 30432 8274 30496
rect 8338 30432 8346 30496
rect 8026 29408 8346 30432
rect 8026 29344 8034 29408
rect 8098 29344 8114 29408
rect 8178 29344 8194 29408
rect 8258 29344 8274 29408
rect 8338 29344 8346 29408
rect 8026 28320 8346 29344
rect 8026 28256 8034 28320
rect 8098 28256 8114 28320
rect 8178 28256 8194 28320
rect 8258 28256 8274 28320
rect 8338 28256 8346 28320
rect 8026 27232 8346 28256
rect 8026 27168 8034 27232
rect 8098 27168 8114 27232
rect 8178 27168 8194 27232
rect 8258 27168 8274 27232
rect 8338 27168 8346 27232
rect 8026 26144 8346 27168
rect 8026 26080 8034 26144
rect 8098 26080 8114 26144
rect 8178 26080 8194 26144
rect 8258 26080 8274 26144
rect 8338 26080 8346 26144
rect 8026 25056 8346 26080
rect 8026 24992 8034 25056
rect 8098 24992 8114 25056
rect 8178 24992 8194 25056
rect 8258 24992 8274 25056
rect 8338 24992 8346 25056
rect 8026 23968 8346 24992
rect 8026 23904 8034 23968
rect 8098 23904 8114 23968
rect 8178 23904 8194 23968
rect 8258 23904 8274 23968
rect 8338 23904 8346 23968
rect 8026 22880 8346 23904
rect 8026 22816 8034 22880
rect 8098 22816 8114 22880
rect 8178 22816 8194 22880
rect 8258 22816 8274 22880
rect 8338 22816 8346 22880
rect 8026 21792 8346 22816
rect 8026 21728 8034 21792
rect 8098 21728 8114 21792
rect 8178 21728 8194 21792
rect 8258 21728 8274 21792
rect 8338 21728 8346 21792
rect 8026 20704 8346 21728
rect 8026 20640 8034 20704
rect 8098 20640 8114 20704
rect 8178 20640 8194 20704
rect 8258 20640 8274 20704
rect 8338 20640 8346 20704
rect 8026 19616 8346 20640
rect 8026 19552 8034 19616
rect 8098 19552 8114 19616
rect 8178 19552 8194 19616
rect 8258 19552 8274 19616
rect 8338 19552 8346 19616
rect 8026 18528 8346 19552
rect 11568 29952 11888 30512
rect 11568 29888 11576 29952
rect 11640 29888 11656 29952
rect 11720 29888 11736 29952
rect 11800 29888 11816 29952
rect 11880 29888 11888 29952
rect 11568 28864 11888 29888
rect 11568 28800 11576 28864
rect 11640 28800 11656 28864
rect 11720 28800 11736 28864
rect 11800 28800 11816 28864
rect 11880 28800 11888 28864
rect 11568 27776 11888 28800
rect 11568 27712 11576 27776
rect 11640 27712 11656 27776
rect 11720 27712 11736 27776
rect 11800 27712 11816 27776
rect 11880 27712 11888 27776
rect 11568 26688 11888 27712
rect 11568 26624 11576 26688
rect 11640 26624 11656 26688
rect 11720 26624 11736 26688
rect 11800 26624 11816 26688
rect 11880 26624 11888 26688
rect 11568 25600 11888 26624
rect 11568 25536 11576 25600
rect 11640 25536 11656 25600
rect 11720 25536 11736 25600
rect 11800 25536 11816 25600
rect 11880 25536 11888 25600
rect 11568 24512 11888 25536
rect 11568 24448 11576 24512
rect 11640 24448 11656 24512
rect 11720 24448 11736 24512
rect 11800 24448 11816 24512
rect 11880 24448 11888 24512
rect 11568 23424 11888 24448
rect 11568 23360 11576 23424
rect 11640 23360 11656 23424
rect 11720 23360 11736 23424
rect 11800 23360 11816 23424
rect 11880 23360 11888 23424
rect 11568 22336 11888 23360
rect 11568 22272 11576 22336
rect 11640 22272 11656 22336
rect 11720 22272 11736 22336
rect 11800 22272 11816 22336
rect 11880 22272 11888 22336
rect 11568 21248 11888 22272
rect 11568 21184 11576 21248
rect 11640 21184 11656 21248
rect 11720 21184 11736 21248
rect 11800 21184 11816 21248
rect 11880 21184 11888 21248
rect 11568 20160 11888 21184
rect 11568 20096 11576 20160
rect 11640 20096 11656 20160
rect 11720 20096 11736 20160
rect 11800 20096 11816 20160
rect 11880 20096 11888 20160
rect 10179 19412 10245 19413
rect 10179 19348 10180 19412
rect 10244 19348 10245 19412
rect 10179 19347 10245 19348
rect 8026 18464 8034 18528
rect 8098 18464 8114 18528
rect 8178 18464 8194 18528
rect 8258 18464 8274 18528
rect 8338 18464 8346 18528
rect 8026 17440 8346 18464
rect 8026 17376 8034 17440
rect 8098 17376 8114 17440
rect 8178 17376 8194 17440
rect 8258 17376 8274 17440
rect 8338 17376 8346 17440
rect 8026 16352 8346 17376
rect 8026 16288 8034 16352
rect 8098 16288 8114 16352
rect 8178 16288 8194 16352
rect 8258 16288 8274 16352
rect 8338 16288 8346 16352
rect 8026 15264 8346 16288
rect 8026 15200 8034 15264
rect 8098 15200 8114 15264
rect 8178 15200 8194 15264
rect 8258 15200 8274 15264
rect 8338 15200 8346 15264
rect 8026 14176 8346 15200
rect 8026 14112 8034 14176
rect 8098 14112 8114 14176
rect 8178 14112 8194 14176
rect 8258 14112 8274 14176
rect 8338 14112 8346 14176
rect 8026 13088 8346 14112
rect 8026 13024 8034 13088
rect 8098 13024 8114 13088
rect 8178 13024 8194 13088
rect 8258 13024 8274 13088
rect 8338 13024 8346 13088
rect 8026 12000 8346 13024
rect 8026 11936 8034 12000
rect 8098 11936 8114 12000
rect 8178 11936 8194 12000
rect 8258 11936 8274 12000
rect 8338 11936 8346 12000
rect 8026 10912 8346 11936
rect 8026 10848 8034 10912
rect 8098 10848 8114 10912
rect 8178 10848 8194 10912
rect 8258 10848 8274 10912
rect 8338 10848 8346 10912
rect 8026 9824 8346 10848
rect 8026 9760 8034 9824
rect 8098 9760 8114 9824
rect 8178 9760 8194 9824
rect 8258 9760 8274 9824
rect 8338 9760 8346 9824
rect 8026 8736 8346 9760
rect 10182 9485 10242 19347
rect 11568 19072 11888 20096
rect 11568 19008 11576 19072
rect 11640 19008 11656 19072
rect 11720 19008 11736 19072
rect 11800 19008 11816 19072
rect 11880 19008 11888 19072
rect 11568 17984 11888 19008
rect 11568 17920 11576 17984
rect 11640 17920 11656 17984
rect 11720 17920 11736 17984
rect 11800 17920 11816 17984
rect 11880 17920 11888 17984
rect 11568 16896 11888 17920
rect 11568 16832 11576 16896
rect 11640 16832 11656 16896
rect 11720 16832 11736 16896
rect 11800 16832 11816 16896
rect 11880 16832 11888 16896
rect 11568 15808 11888 16832
rect 11568 15744 11576 15808
rect 11640 15744 11656 15808
rect 11720 15744 11736 15808
rect 11800 15744 11816 15808
rect 11880 15744 11888 15808
rect 11568 14720 11888 15744
rect 11568 14656 11576 14720
rect 11640 14656 11656 14720
rect 11720 14656 11736 14720
rect 11800 14656 11816 14720
rect 11880 14656 11888 14720
rect 11568 13632 11888 14656
rect 11568 13568 11576 13632
rect 11640 13568 11656 13632
rect 11720 13568 11736 13632
rect 11800 13568 11816 13632
rect 11880 13568 11888 13632
rect 10547 13292 10613 13293
rect 10547 13228 10548 13292
rect 10612 13228 10613 13292
rect 10547 13227 10613 13228
rect 10179 9484 10245 9485
rect 10179 9420 10180 9484
rect 10244 9420 10245 9484
rect 10179 9419 10245 9420
rect 8026 8672 8034 8736
rect 8098 8672 8114 8736
rect 8178 8672 8194 8736
rect 8258 8672 8274 8736
rect 8338 8672 8346 8736
rect 8026 7648 8346 8672
rect 10550 8261 10610 13227
rect 11568 12544 11888 13568
rect 11568 12480 11576 12544
rect 11640 12480 11656 12544
rect 11720 12480 11736 12544
rect 11800 12480 11816 12544
rect 11880 12480 11888 12544
rect 11568 11456 11888 12480
rect 11568 11392 11576 11456
rect 11640 11392 11656 11456
rect 11720 11392 11736 11456
rect 11800 11392 11816 11456
rect 11880 11392 11888 11456
rect 11568 10368 11888 11392
rect 11568 10304 11576 10368
rect 11640 10304 11656 10368
rect 11720 10304 11736 10368
rect 11800 10304 11816 10368
rect 11880 10304 11888 10368
rect 11568 9280 11888 10304
rect 11568 9216 11576 9280
rect 11640 9216 11656 9280
rect 11720 9216 11736 9280
rect 11800 9216 11816 9280
rect 11880 9216 11888 9280
rect 10547 8260 10613 8261
rect 10547 8196 10548 8260
rect 10612 8196 10613 8260
rect 10547 8195 10613 8196
rect 8026 7584 8034 7648
rect 8098 7584 8114 7648
rect 8178 7584 8194 7648
rect 8258 7584 8274 7648
rect 8338 7584 8346 7648
rect 8026 6560 8346 7584
rect 8026 6496 8034 6560
rect 8098 6496 8114 6560
rect 8178 6496 8194 6560
rect 8258 6496 8274 6560
rect 8338 6496 8346 6560
rect 8026 5472 8346 6496
rect 8026 5408 8034 5472
rect 8098 5408 8114 5472
rect 8178 5408 8194 5472
rect 8258 5408 8274 5472
rect 8338 5408 8346 5472
rect 8026 4384 8346 5408
rect 8026 4320 8034 4384
rect 8098 4320 8114 4384
rect 8178 4320 8194 4384
rect 8258 4320 8274 4384
rect 8338 4320 8346 4384
rect 8026 3296 8346 4320
rect 8026 3232 8034 3296
rect 8098 3232 8114 3296
rect 8178 3232 8194 3296
rect 8258 3232 8274 3296
rect 8338 3232 8346 3296
rect 8026 2208 8346 3232
rect 8026 2144 8034 2208
rect 8098 2144 8114 2208
rect 8178 2144 8194 2208
rect 8258 2144 8274 2208
rect 8338 2144 8346 2208
rect 8026 2128 8346 2144
rect 11568 8192 11888 9216
rect 11568 8128 11576 8192
rect 11640 8128 11656 8192
rect 11720 8128 11736 8192
rect 11800 8128 11816 8192
rect 11880 8128 11888 8192
rect 11568 7104 11888 8128
rect 11568 7040 11576 7104
rect 11640 7040 11656 7104
rect 11720 7040 11736 7104
rect 11800 7040 11816 7104
rect 11880 7040 11888 7104
rect 11568 6016 11888 7040
rect 11568 5952 11576 6016
rect 11640 5952 11656 6016
rect 11720 5952 11736 6016
rect 11800 5952 11816 6016
rect 11880 5952 11888 6016
rect 11568 4928 11888 5952
rect 11568 4864 11576 4928
rect 11640 4864 11656 4928
rect 11720 4864 11736 4928
rect 11800 4864 11816 4928
rect 11880 4864 11888 4928
rect 11568 3840 11888 4864
rect 11568 3776 11576 3840
rect 11640 3776 11656 3840
rect 11720 3776 11736 3840
rect 11800 3776 11816 3840
rect 11880 3776 11888 3840
rect 11568 2752 11888 3776
rect 11568 2688 11576 2752
rect 11640 2688 11656 2752
rect 11720 2688 11736 2752
rect 11800 2688 11816 2752
rect 11880 2688 11888 2752
rect 11568 2128 11888 2688
rect 15109 30496 15429 30512
rect 15109 30432 15117 30496
rect 15181 30432 15197 30496
rect 15261 30432 15277 30496
rect 15341 30432 15357 30496
rect 15421 30432 15429 30496
rect 15109 29408 15429 30432
rect 15109 29344 15117 29408
rect 15181 29344 15197 29408
rect 15261 29344 15277 29408
rect 15341 29344 15357 29408
rect 15421 29344 15429 29408
rect 15109 28320 15429 29344
rect 15109 28256 15117 28320
rect 15181 28256 15197 28320
rect 15261 28256 15277 28320
rect 15341 28256 15357 28320
rect 15421 28256 15429 28320
rect 15109 27232 15429 28256
rect 15109 27168 15117 27232
rect 15181 27168 15197 27232
rect 15261 27168 15277 27232
rect 15341 27168 15357 27232
rect 15421 27168 15429 27232
rect 15109 26144 15429 27168
rect 15109 26080 15117 26144
rect 15181 26080 15197 26144
rect 15261 26080 15277 26144
rect 15341 26080 15357 26144
rect 15421 26080 15429 26144
rect 15109 25056 15429 26080
rect 15109 24992 15117 25056
rect 15181 24992 15197 25056
rect 15261 24992 15277 25056
rect 15341 24992 15357 25056
rect 15421 24992 15429 25056
rect 15109 23968 15429 24992
rect 15109 23904 15117 23968
rect 15181 23904 15197 23968
rect 15261 23904 15277 23968
rect 15341 23904 15357 23968
rect 15421 23904 15429 23968
rect 15109 22880 15429 23904
rect 15109 22816 15117 22880
rect 15181 22816 15197 22880
rect 15261 22816 15277 22880
rect 15341 22816 15357 22880
rect 15421 22816 15429 22880
rect 15109 21792 15429 22816
rect 15109 21728 15117 21792
rect 15181 21728 15197 21792
rect 15261 21728 15277 21792
rect 15341 21728 15357 21792
rect 15421 21728 15429 21792
rect 15109 20704 15429 21728
rect 18651 29952 18971 30512
rect 18651 29888 18659 29952
rect 18723 29888 18739 29952
rect 18803 29888 18819 29952
rect 18883 29888 18899 29952
rect 18963 29888 18971 29952
rect 18651 28864 18971 29888
rect 18651 28800 18659 28864
rect 18723 28800 18739 28864
rect 18803 28800 18819 28864
rect 18883 28800 18899 28864
rect 18963 28800 18971 28864
rect 18651 27776 18971 28800
rect 18651 27712 18659 27776
rect 18723 27712 18739 27776
rect 18803 27712 18819 27776
rect 18883 27712 18899 27776
rect 18963 27712 18971 27776
rect 18651 26688 18971 27712
rect 18651 26624 18659 26688
rect 18723 26624 18739 26688
rect 18803 26624 18819 26688
rect 18883 26624 18899 26688
rect 18963 26624 18971 26688
rect 18651 25600 18971 26624
rect 18651 25536 18659 25600
rect 18723 25536 18739 25600
rect 18803 25536 18819 25600
rect 18883 25536 18899 25600
rect 18963 25536 18971 25600
rect 18651 24512 18971 25536
rect 18651 24448 18659 24512
rect 18723 24448 18739 24512
rect 18803 24448 18819 24512
rect 18883 24448 18899 24512
rect 18963 24448 18971 24512
rect 18651 23424 18971 24448
rect 18651 23360 18659 23424
rect 18723 23360 18739 23424
rect 18803 23360 18819 23424
rect 18883 23360 18899 23424
rect 18963 23360 18971 23424
rect 18651 22336 18971 23360
rect 18651 22272 18659 22336
rect 18723 22272 18739 22336
rect 18803 22272 18819 22336
rect 18883 22272 18899 22336
rect 18963 22272 18971 22336
rect 18651 21248 18971 22272
rect 18651 21184 18659 21248
rect 18723 21184 18739 21248
rect 18803 21184 18819 21248
rect 18883 21184 18899 21248
rect 18963 21184 18971 21248
rect 16251 20772 16317 20773
rect 16251 20708 16252 20772
rect 16316 20708 16317 20772
rect 16251 20707 16317 20708
rect 15109 20640 15117 20704
rect 15181 20640 15197 20704
rect 15261 20640 15277 20704
rect 15341 20640 15357 20704
rect 15421 20640 15429 20704
rect 15109 19616 15429 20640
rect 15109 19552 15117 19616
rect 15181 19552 15197 19616
rect 15261 19552 15277 19616
rect 15341 19552 15357 19616
rect 15421 19552 15429 19616
rect 15109 18528 15429 19552
rect 15109 18464 15117 18528
rect 15181 18464 15197 18528
rect 15261 18464 15277 18528
rect 15341 18464 15357 18528
rect 15421 18464 15429 18528
rect 15109 17440 15429 18464
rect 15109 17376 15117 17440
rect 15181 17376 15197 17440
rect 15261 17376 15277 17440
rect 15341 17376 15357 17440
rect 15421 17376 15429 17440
rect 15109 16352 15429 17376
rect 15109 16288 15117 16352
rect 15181 16288 15197 16352
rect 15261 16288 15277 16352
rect 15341 16288 15357 16352
rect 15421 16288 15429 16352
rect 15109 15264 15429 16288
rect 15109 15200 15117 15264
rect 15181 15200 15197 15264
rect 15261 15200 15277 15264
rect 15341 15200 15357 15264
rect 15421 15200 15429 15264
rect 15109 14176 15429 15200
rect 16254 15197 16314 20707
rect 18651 20160 18971 21184
rect 18651 20096 18659 20160
rect 18723 20096 18739 20160
rect 18803 20096 18819 20160
rect 18883 20096 18899 20160
rect 18963 20096 18971 20160
rect 18651 19072 18971 20096
rect 18651 19008 18659 19072
rect 18723 19008 18739 19072
rect 18803 19008 18819 19072
rect 18883 19008 18899 19072
rect 18963 19008 18971 19072
rect 18651 17984 18971 19008
rect 18651 17920 18659 17984
rect 18723 17920 18739 17984
rect 18803 17920 18819 17984
rect 18883 17920 18899 17984
rect 18963 17920 18971 17984
rect 18651 16896 18971 17920
rect 18651 16832 18659 16896
rect 18723 16832 18739 16896
rect 18803 16832 18819 16896
rect 18883 16832 18899 16896
rect 18963 16832 18971 16896
rect 18651 15808 18971 16832
rect 18651 15744 18659 15808
rect 18723 15744 18739 15808
rect 18803 15744 18819 15808
rect 18883 15744 18899 15808
rect 18963 15744 18971 15808
rect 16251 15196 16317 15197
rect 16251 15132 16252 15196
rect 16316 15132 16317 15196
rect 16251 15131 16317 15132
rect 15109 14112 15117 14176
rect 15181 14112 15197 14176
rect 15261 14112 15277 14176
rect 15341 14112 15357 14176
rect 15421 14112 15429 14176
rect 15109 13088 15429 14112
rect 15109 13024 15117 13088
rect 15181 13024 15197 13088
rect 15261 13024 15277 13088
rect 15341 13024 15357 13088
rect 15421 13024 15429 13088
rect 15109 12000 15429 13024
rect 15109 11936 15117 12000
rect 15181 11936 15197 12000
rect 15261 11936 15277 12000
rect 15341 11936 15357 12000
rect 15421 11936 15429 12000
rect 15109 10912 15429 11936
rect 15109 10848 15117 10912
rect 15181 10848 15197 10912
rect 15261 10848 15277 10912
rect 15341 10848 15357 10912
rect 15421 10848 15429 10912
rect 15109 9824 15429 10848
rect 15109 9760 15117 9824
rect 15181 9760 15197 9824
rect 15261 9760 15277 9824
rect 15341 9760 15357 9824
rect 15421 9760 15429 9824
rect 15109 8736 15429 9760
rect 15109 8672 15117 8736
rect 15181 8672 15197 8736
rect 15261 8672 15277 8736
rect 15341 8672 15357 8736
rect 15421 8672 15429 8736
rect 15109 7648 15429 8672
rect 15109 7584 15117 7648
rect 15181 7584 15197 7648
rect 15261 7584 15277 7648
rect 15341 7584 15357 7648
rect 15421 7584 15429 7648
rect 15109 6560 15429 7584
rect 15109 6496 15117 6560
rect 15181 6496 15197 6560
rect 15261 6496 15277 6560
rect 15341 6496 15357 6560
rect 15421 6496 15429 6560
rect 15109 5472 15429 6496
rect 15109 5408 15117 5472
rect 15181 5408 15197 5472
rect 15261 5408 15277 5472
rect 15341 5408 15357 5472
rect 15421 5408 15429 5472
rect 15109 4384 15429 5408
rect 15109 4320 15117 4384
rect 15181 4320 15197 4384
rect 15261 4320 15277 4384
rect 15341 4320 15357 4384
rect 15421 4320 15429 4384
rect 15109 3296 15429 4320
rect 15109 3232 15117 3296
rect 15181 3232 15197 3296
rect 15261 3232 15277 3296
rect 15341 3232 15357 3296
rect 15421 3232 15429 3296
rect 15109 2208 15429 3232
rect 15109 2144 15117 2208
rect 15181 2144 15197 2208
rect 15261 2144 15277 2208
rect 15341 2144 15357 2208
rect 15421 2144 15429 2208
rect 15109 2128 15429 2144
rect 18651 14720 18971 15744
rect 18651 14656 18659 14720
rect 18723 14656 18739 14720
rect 18803 14656 18819 14720
rect 18883 14656 18899 14720
rect 18963 14656 18971 14720
rect 18651 13632 18971 14656
rect 18651 13568 18659 13632
rect 18723 13568 18739 13632
rect 18803 13568 18819 13632
rect 18883 13568 18899 13632
rect 18963 13568 18971 13632
rect 18651 12544 18971 13568
rect 18651 12480 18659 12544
rect 18723 12480 18739 12544
rect 18803 12480 18819 12544
rect 18883 12480 18899 12544
rect 18963 12480 18971 12544
rect 18651 11456 18971 12480
rect 18651 11392 18659 11456
rect 18723 11392 18739 11456
rect 18803 11392 18819 11456
rect 18883 11392 18899 11456
rect 18963 11392 18971 11456
rect 18651 10368 18971 11392
rect 18651 10304 18659 10368
rect 18723 10304 18739 10368
rect 18803 10304 18819 10368
rect 18883 10304 18899 10368
rect 18963 10304 18971 10368
rect 18651 9280 18971 10304
rect 18651 9216 18659 9280
rect 18723 9216 18739 9280
rect 18803 9216 18819 9280
rect 18883 9216 18899 9280
rect 18963 9216 18971 9280
rect 18651 8192 18971 9216
rect 18651 8128 18659 8192
rect 18723 8128 18739 8192
rect 18803 8128 18819 8192
rect 18883 8128 18899 8192
rect 18963 8128 18971 8192
rect 18651 7104 18971 8128
rect 18651 7040 18659 7104
rect 18723 7040 18739 7104
rect 18803 7040 18819 7104
rect 18883 7040 18899 7104
rect 18963 7040 18971 7104
rect 18651 6016 18971 7040
rect 18651 5952 18659 6016
rect 18723 5952 18739 6016
rect 18803 5952 18819 6016
rect 18883 5952 18899 6016
rect 18963 5952 18971 6016
rect 18651 4928 18971 5952
rect 18651 4864 18659 4928
rect 18723 4864 18739 4928
rect 18803 4864 18819 4928
rect 18883 4864 18899 4928
rect 18963 4864 18971 4928
rect 18651 3840 18971 4864
rect 18651 3776 18659 3840
rect 18723 3776 18739 3840
rect 18803 3776 18819 3840
rect 18883 3776 18899 3840
rect 18963 3776 18971 3840
rect 18651 2752 18971 3776
rect 18651 2688 18659 2752
rect 18723 2688 18739 2752
rect 18803 2688 18819 2752
rect 18883 2688 18899 2752
rect 18963 2688 18971 2752
rect 18651 2128 18971 2688
rect 22192 30496 22512 30512
rect 22192 30432 22200 30496
rect 22264 30432 22280 30496
rect 22344 30432 22360 30496
rect 22424 30432 22440 30496
rect 22504 30432 22512 30496
rect 22192 29408 22512 30432
rect 22192 29344 22200 29408
rect 22264 29344 22280 29408
rect 22344 29344 22360 29408
rect 22424 29344 22440 29408
rect 22504 29344 22512 29408
rect 22192 28320 22512 29344
rect 22192 28256 22200 28320
rect 22264 28256 22280 28320
rect 22344 28256 22360 28320
rect 22424 28256 22440 28320
rect 22504 28256 22512 28320
rect 22192 27232 22512 28256
rect 22192 27168 22200 27232
rect 22264 27168 22280 27232
rect 22344 27168 22360 27232
rect 22424 27168 22440 27232
rect 22504 27168 22512 27232
rect 22192 26144 22512 27168
rect 22192 26080 22200 26144
rect 22264 26080 22280 26144
rect 22344 26080 22360 26144
rect 22424 26080 22440 26144
rect 22504 26080 22512 26144
rect 22192 25056 22512 26080
rect 22192 24992 22200 25056
rect 22264 24992 22280 25056
rect 22344 24992 22360 25056
rect 22424 24992 22440 25056
rect 22504 24992 22512 25056
rect 22192 23968 22512 24992
rect 22192 23904 22200 23968
rect 22264 23904 22280 23968
rect 22344 23904 22360 23968
rect 22424 23904 22440 23968
rect 22504 23904 22512 23968
rect 22192 22880 22512 23904
rect 22192 22816 22200 22880
rect 22264 22816 22280 22880
rect 22344 22816 22360 22880
rect 22424 22816 22440 22880
rect 22504 22816 22512 22880
rect 22192 21792 22512 22816
rect 25734 29952 26054 30512
rect 25734 29888 25742 29952
rect 25806 29888 25822 29952
rect 25886 29888 25902 29952
rect 25966 29888 25982 29952
rect 26046 29888 26054 29952
rect 25734 28864 26054 29888
rect 29275 30496 29595 30512
rect 29275 30432 29283 30496
rect 29347 30432 29363 30496
rect 29427 30432 29443 30496
rect 29507 30432 29523 30496
rect 29587 30432 29595 30496
rect 29275 29408 29595 30432
rect 29275 29344 29283 29408
rect 29347 29344 29363 29408
rect 29427 29344 29443 29408
rect 29507 29344 29523 29408
rect 29587 29344 29595 29408
rect 28763 29068 28829 29069
rect 28763 29004 28764 29068
rect 28828 29004 28829 29068
rect 28763 29003 28829 29004
rect 25734 28800 25742 28864
rect 25806 28800 25822 28864
rect 25886 28800 25902 28864
rect 25966 28800 25982 28864
rect 26046 28800 26054 28864
rect 25734 27776 26054 28800
rect 25734 27712 25742 27776
rect 25806 27712 25822 27776
rect 25886 27712 25902 27776
rect 25966 27712 25982 27776
rect 26046 27712 26054 27776
rect 25734 26688 26054 27712
rect 25734 26624 25742 26688
rect 25806 26624 25822 26688
rect 25886 26624 25902 26688
rect 25966 26624 25982 26688
rect 26046 26624 26054 26688
rect 25734 25600 26054 26624
rect 25734 25536 25742 25600
rect 25806 25536 25822 25600
rect 25886 25536 25902 25600
rect 25966 25536 25982 25600
rect 26046 25536 26054 25600
rect 25734 24512 26054 25536
rect 25734 24448 25742 24512
rect 25806 24448 25822 24512
rect 25886 24448 25902 24512
rect 25966 24448 25982 24512
rect 26046 24448 26054 24512
rect 25734 23424 26054 24448
rect 25734 23360 25742 23424
rect 25806 23360 25822 23424
rect 25886 23360 25902 23424
rect 25966 23360 25982 23424
rect 26046 23360 26054 23424
rect 24347 22540 24413 22541
rect 24347 22476 24348 22540
rect 24412 22476 24413 22540
rect 24347 22475 24413 22476
rect 22192 21728 22200 21792
rect 22264 21728 22280 21792
rect 22344 21728 22360 21792
rect 22424 21728 22440 21792
rect 22504 21728 22512 21792
rect 22192 20704 22512 21728
rect 22192 20640 22200 20704
rect 22264 20640 22280 20704
rect 22344 20640 22360 20704
rect 22424 20640 22440 20704
rect 22504 20640 22512 20704
rect 22192 19616 22512 20640
rect 22192 19552 22200 19616
rect 22264 19552 22280 19616
rect 22344 19552 22360 19616
rect 22424 19552 22440 19616
rect 22504 19552 22512 19616
rect 22192 18528 22512 19552
rect 22192 18464 22200 18528
rect 22264 18464 22280 18528
rect 22344 18464 22360 18528
rect 22424 18464 22440 18528
rect 22504 18464 22512 18528
rect 22192 17440 22512 18464
rect 22192 17376 22200 17440
rect 22264 17376 22280 17440
rect 22344 17376 22360 17440
rect 22424 17376 22440 17440
rect 22504 17376 22512 17440
rect 22192 16352 22512 17376
rect 22192 16288 22200 16352
rect 22264 16288 22280 16352
rect 22344 16288 22360 16352
rect 22424 16288 22440 16352
rect 22504 16288 22512 16352
rect 22192 15264 22512 16288
rect 22192 15200 22200 15264
rect 22264 15200 22280 15264
rect 22344 15200 22360 15264
rect 22424 15200 22440 15264
rect 22504 15200 22512 15264
rect 22192 14176 22512 15200
rect 22192 14112 22200 14176
rect 22264 14112 22280 14176
rect 22344 14112 22360 14176
rect 22424 14112 22440 14176
rect 22504 14112 22512 14176
rect 22192 13088 22512 14112
rect 22192 13024 22200 13088
rect 22264 13024 22280 13088
rect 22344 13024 22360 13088
rect 22424 13024 22440 13088
rect 22504 13024 22512 13088
rect 22192 12000 22512 13024
rect 22192 11936 22200 12000
rect 22264 11936 22280 12000
rect 22344 11936 22360 12000
rect 22424 11936 22440 12000
rect 22504 11936 22512 12000
rect 22192 10912 22512 11936
rect 22192 10848 22200 10912
rect 22264 10848 22280 10912
rect 22344 10848 22360 10912
rect 22424 10848 22440 10912
rect 22504 10848 22512 10912
rect 22192 9824 22512 10848
rect 22192 9760 22200 9824
rect 22264 9760 22280 9824
rect 22344 9760 22360 9824
rect 22424 9760 22440 9824
rect 22504 9760 22512 9824
rect 22192 8736 22512 9760
rect 22192 8672 22200 8736
rect 22264 8672 22280 8736
rect 22344 8672 22360 8736
rect 22424 8672 22440 8736
rect 22504 8672 22512 8736
rect 22192 7648 22512 8672
rect 22192 7584 22200 7648
rect 22264 7584 22280 7648
rect 22344 7584 22360 7648
rect 22424 7584 22440 7648
rect 22504 7584 22512 7648
rect 22192 6560 22512 7584
rect 22192 6496 22200 6560
rect 22264 6496 22280 6560
rect 22344 6496 22360 6560
rect 22424 6496 22440 6560
rect 22504 6496 22512 6560
rect 22192 5472 22512 6496
rect 24350 5541 24410 22475
rect 25734 22336 26054 23360
rect 25734 22272 25742 22336
rect 25806 22272 25822 22336
rect 25886 22272 25902 22336
rect 25966 22272 25982 22336
rect 26046 22272 26054 22336
rect 25734 21248 26054 22272
rect 25734 21184 25742 21248
rect 25806 21184 25822 21248
rect 25886 21184 25902 21248
rect 25966 21184 25982 21248
rect 26046 21184 26054 21248
rect 25734 20160 26054 21184
rect 25734 20096 25742 20160
rect 25806 20096 25822 20160
rect 25886 20096 25902 20160
rect 25966 20096 25982 20160
rect 26046 20096 26054 20160
rect 25734 19072 26054 20096
rect 25734 19008 25742 19072
rect 25806 19008 25822 19072
rect 25886 19008 25902 19072
rect 25966 19008 25982 19072
rect 26046 19008 26054 19072
rect 25734 17984 26054 19008
rect 25734 17920 25742 17984
rect 25806 17920 25822 17984
rect 25886 17920 25902 17984
rect 25966 17920 25982 17984
rect 26046 17920 26054 17984
rect 25734 16896 26054 17920
rect 27659 17236 27725 17237
rect 27659 17172 27660 17236
rect 27724 17172 27725 17236
rect 27659 17171 27725 17172
rect 25734 16832 25742 16896
rect 25806 16832 25822 16896
rect 25886 16832 25902 16896
rect 25966 16832 25982 16896
rect 26046 16832 26054 16896
rect 25734 15808 26054 16832
rect 25734 15744 25742 15808
rect 25806 15744 25822 15808
rect 25886 15744 25902 15808
rect 25966 15744 25982 15808
rect 26046 15744 26054 15808
rect 25734 14720 26054 15744
rect 25734 14656 25742 14720
rect 25806 14656 25822 14720
rect 25886 14656 25902 14720
rect 25966 14656 25982 14720
rect 26046 14656 26054 14720
rect 25734 13632 26054 14656
rect 25734 13568 25742 13632
rect 25806 13568 25822 13632
rect 25886 13568 25902 13632
rect 25966 13568 25982 13632
rect 26046 13568 26054 13632
rect 25734 12544 26054 13568
rect 25734 12480 25742 12544
rect 25806 12480 25822 12544
rect 25886 12480 25902 12544
rect 25966 12480 25982 12544
rect 26046 12480 26054 12544
rect 25734 11456 26054 12480
rect 27662 11797 27722 17171
rect 27659 11796 27725 11797
rect 27659 11732 27660 11796
rect 27724 11732 27725 11796
rect 27659 11731 27725 11732
rect 25734 11392 25742 11456
rect 25806 11392 25822 11456
rect 25886 11392 25902 11456
rect 25966 11392 25982 11456
rect 26046 11392 26054 11456
rect 25734 10368 26054 11392
rect 25734 10304 25742 10368
rect 25806 10304 25822 10368
rect 25886 10304 25902 10368
rect 25966 10304 25982 10368
rect 26046 10304 26054 10368
rect 25734 9280 26054 10304
rect 25734 9216 25742 9280
rect 25806 9216 25822 9280
rect 25886 9216 25902 9280
rect 25966 9216 25982 9280
rect 26046 9216 26054 9280
rect 25734 8192 26054 9216
rect 25734 8128 25742 8192
rect 25806 8128 25822 8192
rect 25886 8128 25902 8192
rect 25966 8128 25982 8192
rect 26046 8128 26054 8192
rect 25734 7104 26054 8128
rect 25734 7040 25742 7104
rect 25806 7040 25822 7104
rect 25886 7040 25902 7104
rect 25966 7040 25982 7104
rect 26046 7040 26054 7104
rect 25734 6016 26054 7040
rect 28766 6765 28826 29003
rect 29275 28320 29595 29344
rect 29275 28256 29283 28320
rect 29347 28256 29363 28320
rect 29427 28256 29443 28320
rect 29507 28256 29523 28320
rect 29587 28256 29595 28320
rect 29275 27232 29595 28256
rect 29275 27168 29283 27232
rect 29347 27168 29363 27232
rect 29427 27168 29443 27232
rect 29507 27168 29523 27232
rect 29587 27168 29595 27232
rect 29275 26144 29595 27168
rect 29275 26080 29283 26144
rect 29347 26080 29363 26144
rect 29427 26080 29443 26144
rect 29507 26080 29523 26144
rect 29587 26080 29595 26144
rect 29275 25056 29595 26080
rect 29275 24992 29283 25056
rect 29347 24992 29363 25056
rect 29427 24992 29443 25056
rect 29507 24992 29523 25056
rect 29587 24992 29595 25056
rect 29275 23968 29595 24992
rect 29275 23904 29283 23968
rect 29347 23904 29363 23968
rect 29427 23904 29443 23968
rect 29507 23904 29523 23968
rect 29587 23904 29595 23968
rect 29275 22880 29595 23904
rect 29275 22816 29283 22880
rect 29347 22816 29363 22880
rect 29427 22816 29443 22880
rect 29507 22816 29523 22880
rect 29587 22816 29595 22880
rect 29275 21792 29595 22816
rect 29275 21728 29283 21792
rect 29347 21728 29363 21792
rect 29427 21728 29443 21792
rect 29507 21728 29523 21792
rect 29587 21728 29595 21792
rect 29275 20704 29595 21728
rect 29275 20640 29283 20704
rect 29347 20640 29363 20704
rect 29427 20640 29443 20704
rect 29507 20640 29523 20704
rect 29587 20640 29595 20704
rect 29275 19616 29595 20640
rect 29275 19552 29283 19616
rect 29347 19552 29363 19616
rect 29427 19552 29443 19616
rect 29507 19552 29523 19616
rect 29587 19552 29595 19616
rect 29275 18528 29595 19552
rect 29275 18464 29283 18528
rect 29347 18464 29363 18528
rect 29427 18464 29443 18528
rect 29507 18464 29523 18528
rect 29587 18464 29595 18528
rect 29275 17440 29595 18464
rect 29275 17376 29283 17440
rect 29347 17376 29363 17440
rect 29427 17376 29443 17440
rect 29507 17376 29523 17440
rect 29587 17376 29595 17440
rect 29275 16352 29595 17376
rect 29275 16288 29283 16352
rect 29347 16288 29363 16352
rect 29427 16288 29443 16352
rect 29507 16288 29523 16352
rect 29587 16288 29595 16352
rect 29275 15264 29595 16288
rect 29275 15200 29283 15264
rect 29347 15200 29363 15264
rect 29427 15200 29443 15264
rect 29507 15200 29523 15264
rect 29587 15200 29595 15264
rect 29275 14176 29595 15200
rect 29275 14112 29283 14176
rect 29347 14112 29363 14176
rect 29427 14112 29443 14176
rect 29507 14112 29523 14176
rect 29587 14112 29595 14176
rect 29275 13088 29595 14112
rect 29275 13024 29283 13088
rect 29347 13024 29363 13088
rect 29427 13024 29443 13088
rect 29507 13024 29523 13088
rect 29587 13024 29595 13088
rect 29275 12000 29595 13024
rect 29275 11936 29283 12000
rect 29347 11936 29363 12000
rect 29427 11936 29443 12000
rect 29507 11936 29523 12000
rect 29587 11936 29595 12000
rect 29275 10912 29595 11936
rect 29275 10848 29283 10912
rect 29347 10848 29363 10912
rect 29427 10848 29443 10912
rect 29507 10848 29523 10912
rect 29587 10848 29595 10912
rect 29275 9824 29595 10848
rect 29275 9760 29283 9824
rect 29347 9760 29363 9824
rect 29427 9760 29443 9824
rect 29507 9760 29523 9824
rect 29587 9760 29595 9824
rect 29275 8736 29595 9760
rect 29275 8672 29283 8736
rect 29347 8672 29363 8736
rect 29427 8672 29443 8736
rect 29507 8672 29523 8736
rect 29587 8672 29595 8736
rect 29275 7648 29595 8672
rect 29275 7584 29283 7648
rect 29347 7584 29363 7648
rect 29427 7584 29443 7648
rect 29507 7584 29523 7648
rect 29587 7584 29595 7648
rect 28763 6764 28829 6765
rect 28763 6700 28764 6764
rect 28828 6700 28829 6764
rect 28763 6699 28829 6700
rect 25734 5952 25742 6016
rect 25806 5952 25822 6016
rect 25886 5952 25902 6016
rect 25966 5952 25982 6016
rect 26046 5952 26054 6016
rect 24347 5540 24413 5541
rect 24347 5476 24348 5540
rect 24412 5476 24413 5540
rect 24347 5475 24413 5476
rect 22192 5408 22200 5472
rect 22264 5408 22280 5472
rect 22344 5408 22360 5472
rect 22424 5408 22440 5472
rect 22504 5408 22512 5472
rect 22192 4384 22512 5408
rect 22192 4320 22200 4384
rect 22264 4320 22280 4384
rect 22344 4320 22360 4384
rect 22424 4320 22440 4384
rect 22504 4320 22512 4384
rect 22192 3296 22512 4320
rect 22192 3232 22200 3296
rect 22264 3232 22280 3296
rect 22344 3232 22360 3296
rect 22424 3232 22440 3296
rect 22504 3232 22512 3296
rect 22192 2208 22512 3232
rect 22192 2144 22200 2208
rect 22264 2144 22280 2208
rect 22344 2144 22360 2208
rect 22424 2144 22440 2208
rect 22504 2144 22512 2208
rect 22192 2128 22512 2144
rect 25734 4928 26054 5952
rect 25734 4864 25742 4928
rect 25806 4864 25822 4928
rect 25886 4864 25902 4928
rect 25966 4864 25982 4928
rect 26046 4864 26054 4928
rect 25734 3840 26054 4864
rect 25734 3776 25742 3840
rect 25806 3776 25822 3840
rect 25886 3776 25902 3840
rect 25966 3776 25982 3840
rect 26046 3776 26054 3840
rect 25734 2752 26054 3776
rect 25734 2688 25742 2752
rect 25806 2688 25822 2752
rect 25886 2688 25902 2752
rect 25966 2688 25982 2752
rect 26046 2688 26054 2752
rect 25734 2128 26054 2688
rect 29275 6560 29595 7584
rect 29275 6496 29283 6560
rect 29347 6496 29363 6560
rect 29427 6496 29443 6560
rect 29507 6496 29523 6560
rect 29587 6496 29595 6560
rect 29275 5472 29595 6496
rect 29275 5408 29283 5472
rect 29347 5408 29363 5472
rect 29427 5408 29443 5472
rect 29507 5408 29523 5472
rect 29587 5408 29595 5472
rect 29275 4384 29595 5408
rect 29275 4320 29283 4384
rect 29347 4320 29363 4384
rect 29427 4320 29443 4384
rect 29507 4320 29523 4384
rect 29587 4320 29595 4384
rect 29275 3296 29595 4320
rect 29275 3232 29283 3296
rect 29347 3232 29363 3296
rect 29427 3232 29443 3296
rect 29507 3232 29523 3296
rect 29587 3232 29595 3296
rect 29275 2208 29595 3232
rect 29275 2144 29283 2208
rect 29347 2144 29363 2208
rect 29427 2144 29443 2208
rect 29507 2144 29523 2208
rect 29587 2144 29595 2208
rect 29275 2128 29595 2144
use sky130_fd_sc_hd__or4b_1  _0462_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0463_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5244 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0464_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _0465_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _0466_
timestamp 1688980957
transform 1 0 10212 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _0467_
timestamp 1688980957
transform 1 0 21252 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0468_
timestamp 1688980957
transform 1 0 17296 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0469_
timestamp 1688980957
transform 1 0 13432 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0470_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7728 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0471_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8464 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0472_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22080 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_4  _0473_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__or4bb_4  _0474_
timestamp 1688980957
transform 1 0 19044 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_8  _0475_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  _0476_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7176 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  _0477_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9936 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0478_
timestamp 1688980957
transform 1 0 10580 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  _0479_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__and2_1  _0480_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7544 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0481_
timestamp 1688980957
transform 1 0 7544 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _0482_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6716 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0483_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10396 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_4  _0484_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__nor3b_2  _0485_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7268 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0486_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12972 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0487_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13892 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand4b_4  _0488_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__or4b_1  _0489_
timestamp 1688980957
transform 1 0 22080 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0490_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23276 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_8  _0491_
timestamp 1688980957
transform 1 0 22356 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__nor3b_4  _0492_
timestamp 1688980957
transform 1 0 20148 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__a22o_1  _0493_
timestamp 1688980957
transform 1 0 15916 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _0494_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15916 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__a221o_1  _0495_
timestamp 1688980957
transform 1 0 10396 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0496_
timestamp 1688980957
transform 1 0 14076 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0497_
timestamp 1688980957
transform 1 0 16928 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_2  _0498_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15272 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a22oi_2  _0499_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16836 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0500_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8188 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nor3b_1  _0501_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0502_
timestamp 1688980957
transform 1 0 5244 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0503_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0504_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4968 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0505_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0506_
timestamp 1688980957
transform 1 0 16376 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_1  _0507_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0508_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _0509_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17756 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _0510_
timestamp 1688980957
transform 1 0 6624 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor3b_1  _0511_
timestamp 1688980957
transform 1 0 5520 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0512_
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0513_
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0514_
timestamp 1688980957
transform 1 0 6072 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _0515_
timestamp 1688980957
transform 1 0 17572 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0516_
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_2  _0517_
timestamp 1688980957
transform 1 0 17112 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0518_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_2  _0519_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _0520_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0521_
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__nor3b_1  _0522_
timestamp 1688980957
transform 1 0 6992 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0523_
timestamp 1688980957
transform 1 0 5336 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0524_
timestamp 1688980957
transform 1 0 4232 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0525_
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _0526_
timestamp 1688980957
transform 1 0 17664 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0527_
timestamp 1688980957
transform 1 0 16100 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_2  _0528_
timestamp 1688980957
transform 1 0 16836 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _0529_
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0530_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0531_
timestamp 1688980957
transform 1 0 15916 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0532_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17756 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0533_
timestamp 1688980957
transform 1 0 18400 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0534_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18952 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0535_
timestamp 1688980957
transform 1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0536_
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_4  _0537_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__o21ai_1  _0538_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19688 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_2  _0539_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0540_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19596 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0541_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20148 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0542_
timestamp 1688980957
transform 1 0 20608 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0543_
timestamp 1688980957
transform 1 0 20056 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0544_
timestamp 1688980957
transform 1 0 20516 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0545_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19872 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0546_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0547_
timestamp 1688980957
transform 1 0 20056 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0548_
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0549_
timestamp 1688980957
transform 1 0 8188 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0550_
timestamp 1688980957
transform 1 0 4416 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0551_
timestamp 1688980957
transform 1 0 4968 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0552_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4048 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0553_
timestamp 1688980957
transform 1 0 7084 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0554_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6532 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0555_
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0556_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0557_
timestamp 1688980957
transform 1 0 5704 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0558_
timestamp 1688980957
transform 1 0 4968 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0559_
timestamp 1688980957
transform 1 0 4692 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0560_
timestamp 1688980957
transform 1 0 3864 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0561_
timestamp 1688980957
transform 1 0 4232 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0562_
timestamp 1688980957
transform 1 0 3404 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0563_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0564_
timestamp 1688980957
transform 1 0 6164 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0565_
timestamp 1688980957
transform 1 0 5244 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0566_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5520 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0568_
timestamp 1688980957
transform 1 0 7360 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0569_
timestamp 1688980957
transform 1 0 7084 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0570_
timestamp 1688980957
transform 1 0 7176 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0571_
timestamp 1688980957
transform 1 0 6624 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0572_
timestamp 1688980957
transform 1 0 7636 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0573_
timestamp 1688980957
transform 1 0 8740 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0574_
timestamp 1688980957
transform 1 0 6900 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0575_
timestamp 1688980957
transform 1 0 9476 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0576_
timestamp 1688980957
transform 1 0 10304 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0577_
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0578_
timestamp 1688980957
transform 1 0 9936 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0579_
timestamp 1688980957
transform 1 0 11040 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0580_
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0581_
timestamp 1688980957
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0582_
timestamp 1688980957
transform 1 0 10488 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0583_
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0584_
timestamp 1688980957
transform 1 0 11960 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0585_
timestamp 1688980957
transform 1 0 11316 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _0586_
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0587_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12420 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0588_
timestamp 1688980957
transform 1 0 12972 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0589_
timestamp 1688980957
transform 1 0 14352 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0590_
timestamp 1688980957
transform 1 0 16008 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0591_
timestamp 1688980957
transform 1 0 15456 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0592_
timestamp 1688980957
transform 1 0 13156 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0593_
timestamp 1688980957
transform 1 0 14904 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0594_
timestamp 1688980957
transform 1 0 16008 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0595_
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0596_
timestamp 1688980957
transform 1 0 16100 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1688980957
transform 1 0 17296 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0598_
timestamp 1688980957
transform 1 0 16652 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0599_
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0600_
timestamp 1688980957
transform 1 0 18032 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0601_
timestamp 1688980957
transform 1 0 17112 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0602_
timestamp 1688980957
transform 1 0 16192 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0603_
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0604_
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0605_
timestamp 1688980957
transform 1 0 21712 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0606_
timestamp 1688980957
transform 1 0 20792 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0607_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22540 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0608_
timestamp 1688980957
transform 1 0 22172 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0609_
timestamp 1688980957
transform 1 0 22632 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0610_
timestamp 1688980957
transform 1 0 23092 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0611_
timestamp 1688980957
transform 1 0 22448 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0612_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22080 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0613_
timestamp 1688980957
transform 1 0 20608 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0614_
timestamp 1688980957
transform 1 0 20148 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0615_
timestamp 1688980957
transform 1 0 20608 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0616_
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0617_
timestamp 1688980957
transform 1 0 6992 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0618_
timestamp 1688980957
transform 1 0 15732 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0619_
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _0620_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1688980957
transform 1 0 6164 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0622_
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0623_
timestamp 1688980957
transform 1 0 5612 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0624_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0625_
timestamp 1688980957
transform 1 0 18860 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0626_
timestamp 1688980957
transform 1 0 16836 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0627_
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_4  _0628_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19044 0 -1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0629_
timestamp 1688980957
transform 1 0 11408 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0630_
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0631_
timestamp 1688980957
transform 1 0 19136 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0632_
timestamp 1688980957
transform 1 0 19320 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_4  _0633_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__a221o_1  _0634_
timestamp 1688980957
transform 1 0 10396 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0635_
timestamp 1688980957
transform 1 0 12052 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0636_
timestamp 1688980957
transform 1 0 17940 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0637_
timestamp 1688980957
transform 1 0 20240 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0638_
timestamp 1688980957
transform 1 0 19964 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _0639_
timestamp 1688980957
transform 1 0 18584 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _0640_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20792 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0641_
timestamp 1688980957
transform 1 0 7268 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0642_
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0643_
timestamp 1688980957
transform 1 0 19872 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0644_
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _0645_
timestamp 1688980957
transform 1 0 18676 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_4  _0646_
timestamp 1688980957
transform 1 0 21896 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1688980957
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0648_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20148 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0649_
timestamp 1688980957
transform 1 0 18492 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0650_
timestamp 1688980957
transform 1 0 20884 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0651_
timestamp 1688980957
transform 1 0 20332 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0652_
timestamp 1688980957
transform 1 0 25024 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0653_
timestamp 1688980957
transform 1 0 23092 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0654_
timestamp 1688980957
transform 1 0 22724 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _0655_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23276 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0656_
timestamp 1688980957
transform 1 0 23460 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0657_
timestamp 1688980957
transform 1 0 24932 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0658_
timestamp 1688980957
transform 1 0 21252 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0659_
timestamp 1688980957
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0660_
timestamp 1688980957
transform 1 0 24564 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0661_
timestamp 1688980957
transform 1 0 25208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0662_
timestamp 1688980957
transform 1 0 21712 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0663_
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0664_
timestamp 1688980957
transform 1 0 25484 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _0665_
timestamp 1688980957
transform 1 0 23460 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0666_
timestamp 1688980957
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0667_
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0668_
timestamp 1688980957
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0669_
timestamp 1688980957
transform 1 0 24840 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0670_
timestamp 1688980957
transform 1 0 23644 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0671_
timestamp 1688980957
transform 1 0 24380 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1688980957
transform 1 0 21068 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0673_
timestamp 1688980957
transform 1 0 20792 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1688980957
transform 1 0 12052 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_4  _0675_
timestamp 1688980957
transform 1 0 19780 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__nand2b_4  _0676_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11684 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_8  _0677_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11776 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_1  _0678_
timestamp 1688980957
transform 1 0 22080 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0679_
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  _0680_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23184 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _0681_
timestamp 1688980957
transform 1 0 16008 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0682_
timestamp 1688980957
transform 1 0 14996 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0683_
timestamp 1688980957
transform 1 0 15916 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0684_
timestamp 1688980957
transform 1 0 17296 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0685_
timestamp 1688980957
transform 1 0 18216 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0686_
timestamp 1688980957
transform 1 0 14904 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0687_
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0688_
timestamp 1688980957
transform 1 0 15732 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0689_
timestamp 1688980957
transform 1 0 15640 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0690_
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0691_
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0692_
timestamp 1688980957
transform 1 0 17940 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0693_
timestamp 1688980957
transform 1 0 14904 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0694_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22356 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _0695_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _0696_
timestamp 1688980957
transform 1 0 10304 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1688980957
transform 1 0 9936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_2  _0698_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12696 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0699_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10212 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _0700_
timestamp 1688980957
transform 1 0 10212 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0701_
timestamp 1688980957
transform 1 0 9384 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0702_
timestamp 1688980957
transform 1 0 8648 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0703_
timestamp 1688980957
transform 1 0 9016 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0704_
timestamp 1688980957
transform 1 0 4600 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0705_
timestamp 1688980957
transform 1 0 5612 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0706_
timestamp 1688980957
transform 1 0 8188 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0707_
timestamp 1688980957
transform 1 0 5244 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0708_
timestamp 1688980957
transform 1 0 5612 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0709_
timestamp 1688980957
transform 1 0 4508 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0710_
timestamp 1688980957
transform 1 0 11500 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0711_
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0712_
timestamp 1688980957
transform 1 0 9844 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0713_
timestamp 1688980957
transform 1 0 11408 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0714_
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _0715_
timestamp 1688980957
transform 1 0 6716 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0716_
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0717_
timestamp 1688980957
transform 1 0 10580 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0718_
timestamp 1688980957
transform 1 0 12052 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0719_
timestamp 1688980957
transform 1 0 6164 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0720_
timestamp 1688980957
transform 1 0 6348 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0721_
timestamp 1688980957
transform 1 0 7268 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0722_
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0723_
timestamp 1688980957
transform 1 0 7268 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0724_
timestamp 1688980957
transform 1 0 6808 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0725_
timestamp 1688980957
transform 1 0 12236 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0726_
timestamp 1688980957
transform 1 0 7452 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0727_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0728_
timestamp 1688980957
transform 1 0 10856 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _0729_
timestamp 1688980957
transform 1 0 11592 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _0730_
timestamp 1688980957
transform 1 0 3956 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0731_
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0732_
timestamp 1688980957
transform 1 0 12788 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0733_
timestamp 1688980957
transform 1 0 14352 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0734_
timestamp 1688980957
transform 1 0 4968 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0735_
timestamp 1688980957
transform 1 0 3312 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0736_
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0737_
timestamp 1688980957
transform 1 0 7084 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0738_
timestamp 1688980957
transform 1 0 4600 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0739_
timestamp 1688980957
transform 1 0 3772 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0740_
timestamp 1688980957
transform 1 0 14812 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0741_
timestamp 1688980957
transform 1 0 5060 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0742_
timestamp 1688980957
transform 1 0 11868 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0743_
timestamp 1688980957
transform 1 0 10948 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0744_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0745_
timestamp 1688980957
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _0746_
timestamp 1688980957
transform 1 0 3956 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0747_
timestamp 1688980957
transform 1 0 10028 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0748_
timestamp 1688980957
transform 1 0 12236 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0749_
timestamp 1688980957
transform 1 0 10304 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0750_
timestamp 1688980957
transform 1 0 3956 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0751_
timestamp 1688980957
transform 1 0 3128 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0752_
timestamp 1688980957
transform 1 0 6716 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0753_
timestamp 1688980957
transform 1 0 3312 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0754_
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0755_
timestamp 1688980957
transform 1 0 4600 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0756_
timestamp 1688980957
transform 1 0 9844 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0757_
timestamp 1688980957
transform 1 0 3956 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0758_
timestamp 1688980957
transform 1 0 9844 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0759_
timestamp 1688980957
transform 1 0 11408 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0760_
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0761_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0762_
timestamp 1688980957
transform 1 0 20332 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1688980957
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0764_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24656 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _0765_
timestamp 1688980957
transform 1 0 27232 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0766_
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0767_
timestamp 1688980957
transform 1 0 23460 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0768_
timestamp 1688980957
transform 1 0 20516 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0769_
timestamp 1688980957
transform 1 0 20056 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0770_
timestamp 1688980957
transform 1 0 20700 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0771_
timestamp 1688980957
transform 1 0 22908 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0772_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21068 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0773_
timestamp 1688980957
transform 1 0 21068 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0774_
timestamp 1688980957
transform 1 0 24104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0775_
timestamp 1688980957
transform 1 0 23460 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0776_
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _0777_
timestamp 1688980957
transform 1 0 24104 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0778_
timestamp 1688980957
transform 1 0 27508 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0779_
timestamp 1688980957
transform 1 0 27048 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0780_
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0781_
timestamp 1688980957
transform 1 0 22724 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0782_
timestamp 1688980957
transform 1 0 22908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0783_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22172 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0784_
timestamp 1688980957
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0785_
timestamp 1688980957
transform 1 0 20976 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0786_
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _0787_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22172 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0788_
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0789_
timestamp 1688980957
transform 1 0 25300 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0790_
timestamp 1688980957
transform 1 0 27048 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0791_
timestamp 1688980957
transform 1 0 26588 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0792_
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0793_
timestamp 1688980957
transform 1 0 27600 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0794_
timestamp 1688980957
transform 1 0 27416 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0795_
timestamp 1688980957
transform 1 0 27692 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0796_
timestamp 1688980957
transform 1 0 27876 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0797_
timestamp 1688980957
transform 1 0 25852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0798_
timestamp 1688980957
transform 1 0 28244 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0799_
timestamp 1688980957
transform 1 0 28336 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0800_
timestamp 1688980957
transform 1 0 27692 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0801_
timestamp 1688980957
transform 1 0 15548 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0802_
timestamp 1688980957
transform 1 0 18492 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0803_
timestamp 1688980957
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0804_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1688980957
transform 1 0 17480 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0806_
timestamp 1688980957
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0807_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0808_
timestamp 1688980957
transform 1 0 16376 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _0809_
timestamp 1688980957
transform 1 0 18492 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0810_
timestamp 1688980957
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0811_
timestamp 1688980957
transform 1 0 16560 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0812_
timestamp 1688980957
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0813_
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0814_
timestamp 1688980957
transform 1 0 18216 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0815_
timestamp 1688980957
transform 1 0 16744 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0816_
timestamp 1688980957
transform 1 0 17848 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0817_
timestamp 1688980957
transform 1 0 16928 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0818_
timestamp 1688980957
transform 1 0 17204 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0819_
timestamp 1688980957
transform 1 0 15824 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0820_
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0821_
timestamp 1688980957
transform 1 0 8372 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0822_
timestamp 1688980957
transform 1 0 14812 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0823_
timestamp 1688980957
transform 1 0 15364 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1688980957
transform 1 0 14352 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0825_
timestamp 1688980957
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0826_
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0827_
timestamp 1688980957
transform 1 0 12880 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0828_
timestamp 1688980957
transform 1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0829_
timestamp 1688980957
transform 1 0 14812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0830_
timestamp 1688980957
transform 1 0 15364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _0831_
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0832_
timestamp 1688980957
transform 1 0 2208 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1688980957
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0834_
timestamp 1688980957
transform 1 0 13800 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0835_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12788 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0836_
timestamp 1688980957
transform 1 0 13156 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1688980957
transform 1 0 12512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _0838_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12880 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_2  _0839_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0840_
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0841_
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0842_
timestamp 1688980957
transform 1 0 19688 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0843_
timestamp 1688980957
transform 1 0 19228 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _0844_
timestamp 1688980957
transform 1 0 23552 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0845_
timestamp 1688980957
transform 1 0 22448 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_2  _0846_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0847_
timestamp 1688980957
transform 1 0 21344 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0848_
timestamp 1688980957
transform 1 0 17664 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _0849_
timestamp 1688980957
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0850_
timestamp 1688980957
transform 1 0 21620 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0851_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20148 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0852_
timestamp 1688980957
transform 1 0 19964 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0853_
timestamp 1688980957
transform 1 0 20700 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _0854_
timestamp 1688980957
transform 1 0 15732 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1688980957
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0856_
timestamp 1688980957
transform 1 0 18768 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0857_
timestamp 1688980957
transform 1 0 18308 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0858_
timestamp 1688980957
transform 1 0 19044 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0859_
timestamp 1688980957
transform 1 0 18400 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0860_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0861_
timestamp 1688980957
transform 1 0 19688 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0862_
timestamp 1688980957
transform 1 0 19964 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0863_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0864_
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0865_
timestamp 1688980957
transform 1 0 19780 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0866_
timestamp 1688980957
transform 1 0 21712 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0867_
timestamp 1688980957
transform 1 0 23000 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0868_
timestamp 1688980957
transform 1 0 23828 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0869_
timestamp 1688980957
transform 1 0 22264 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0870_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1688980957
transform 1 0 24932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0872_
timestamp 1688980957
transform 1 0 25392 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0873_
timestamp 1688980957
transform 1 0 27416 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0874_
timestamp 1688980957
transform 1 0 28244 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0875_
timestamp 1688980957
transform 1 0 23184 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0876_
timestamp 1688980957
transform 1 0 23092 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0877_
timestamp 1688980957
transform 1 0 22540 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0878_
timestamp 1688980957
transform 1 0 22816 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0879_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22356 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _0880_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _0881_
timestamp 1688980957
transform 1 0 23552 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0882_
timestamp 1688980957
transform 1 0 23276 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0883_
timestamp 1688980957
transform 1 0 23460 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0884_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24196 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0885_
timestamp 1688980957
transform 1 0 21712 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0886_
timestamp 1688980957
transform 1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0887_
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0888_
timestamp 1688980957
transform 1 0 22816 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0889_
timestamp 1688980957
transform 1 0 23092 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0890_
timestamp 1688980957
transform 1 0 22540 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0891_
timestamp 1688980957
transform 1 0 21988 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0892_
timestamp 1688980957
transform 1 0 22356 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0893_
timestamp 1688980957
transform 1 0 23920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0894_
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0895_
timestamp 1688980957
transform 1 0 23368 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _0896_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23368 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0897_
timestamp 1688980957
transform 1 0 24472 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0898_
timestamp 1688980957
transform 1 0 23828 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0899_
timestamp 1688980957
transform 1 0 27508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0900_
timestamp 1688980957
transform 1 0 25852 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0901_
timestamp 1688980957
transform 1 0 24840 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _0902_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0903_
timestamp 1688980957
transform 1 0 27232 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0904_
timestamp 1688980957
transform 1 0 25576 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0905_
timestamp 1688980957
transform 1 0 26312 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0906_
timestamp 1688980957
transform 1 0 28152 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0907_
timestamp 1688980957
transform 1 0 26220 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_2  _0908_
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _0909_
timestamp 1688980957
transform 1 0 27692 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0910_
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0911_
timestamp 1688980957
transform 1 0 25484 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0912_
timestamp 1688980957
transform 1 0 25852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _0913_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26128 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _0914_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25392 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0915_
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _0916_
timestamp 1688980957
transform 1 0 14168 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0917_
timestamp 1688980957
transform 1 0 15640 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0918_
timestamp 1688980957
transform 1 0 17572 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0919_
timestamp 1688980957
transform 1 0 14812 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0920_
timestamp 1688980957
transform 1 0 16376 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0921_
timestamp 1688980957
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0922_
timestamp 1688980957
transform 1 0 2576 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0923_
timestamp 1688980957
transform 1 0 2208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0924_
timestamp 1688980957
transform 1 0 3864 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0925_
timestamp 1688980957
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0926_
timestamp 1688980957
transform 1 0 2668 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0927_
timestamp 1688980957
transform 1 0 13892 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0928_
timestamp 1688980957
transform 1 0 13524 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0929_
timestamp 1688980957
transform 1 0 14168 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1688980957
transform 1 0 12972 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0931_
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0932_
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0933_
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0934_
timestamp 1688980957
transform 1 0 14536 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0935_
timestamp 1688980957
transform 1 0 12972 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0936_
timestamp 1688980957
transform 1 0 13524 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0937_
timestamp 1688980957
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0938_
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0939_
timestamp 1688980957
transform 1 0 13064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0940_
timestamp 1688980957
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0941_
timestamp 1688980957
transform 1 0 26128 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1688980957
transform 1 0 22264 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0943_
timestamp 1688980957
transform 1 0 22540 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0944_
timestamp 1688980957
transform 1 0 22724 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0945_
timestamp 1688980957
transform 1 0 22816 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0946_
timestamp 1688980957
transform 1 0 23552 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0947_
timestamp 1688980957
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0948_
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0949_
timestamp 1688980957
transform 1 0 26128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0950_
timestamp 1688980957
transform 1 0 25668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0951_
timestamp 1688980957
transform 1 0 26680 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0952_
timestamp 1688980957
transform 1 0 26036 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0953_
timestamp 1688980957
transform 1 0 26496 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0954_
timestamp 1688980957
transform 1 0 24472 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0955_
timestamp 1688980957
transform 1 0 27692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0956_
timestamp 1688980957
transform 1 0 26864 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0957_
timestamp 1688980957
transform 1 0 28152 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0958_
timestamp 1688980957
transform 1 0 27232 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0959_
timestamp 1688980957
transform 1 0 27232 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0960_
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0961_
timestamp 1688980957
transform 1 0 26404 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1688980957
transform 1 0 27876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0963_
timestamp 1688980957
transform 1 0 27692 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0964_
timestamp 1688980957
transform 1 0 28152 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0965_
timestamp 1688980957
transform 1 0 27784 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0966_
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0967_
timestamp 1688980957
transform 1 0 26588 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0968_
timestamp 1688980957
transform 1 0 25852 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0969_
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0970_
timestamp 1688980957
transform 1 0 25116 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0971_
timestamp 1688980957
transform 1 0 23644 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0972_
timestamp 1688980957
transform 1 0 18584 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0973_
timestamp 1688980957
transform 1 0 9016 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _0974_
timestamp 1688980957
transform 1 0 9108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0975_
timestamp 1688980957
transform 1 0 11224 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0976_
timestamp 1688980957
transform 1 0 9844 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _0977_
timestamp 1688980957
transform 1 0 10580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0978_
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0979_
timestamp 1688980957
transform 1 0 10304 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0980_
timestamp 1688980957
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0981_
timestamp 1688980957
transform 1 0 10672 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0982_
timestamp 1688980957
transform 1 0 9844 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0983_
timestamp 1688980957
transform 1 0 8464 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0984_
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0985_
timestamp 1688980957
transform 1 0 21988 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0986_
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0987_
timestamp 1688980957
transform 1 0 20792 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0988_
timestamp 1688980957
transform 1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0989_
timestamp 1688980957
transform 1 0 9936 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0990_
timestamp 1688980957
transform 1 0 9200 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0991_
timestamp 1688980957
transform 1 0 10396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0992_
timestamp 1688980957
transform 1 0 9752 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0993_
timestamp 1688980957
transform 1 0 10856 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0994_
timestamp 1688980957
transform 1 0 11224 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0995_
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0996_
timestamp 1688980957
transform 1 0 19320 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0997_
timestamp 1688980957
transform 1 0 17664 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0998_
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0999_
timestamp 1688980957
transform 1 0 19780 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1000_
timestamp 1688980957
transform 1 0 18400 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1001_
timestamp 1688980957
transform 1 0 17572 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1002_
timestamp 1688980957
transform 1 0 16928 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1688980957
transform 1 0 16836 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1004_
timestamp 1688980957
transform 1 0 15640 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1005_
timestamp 1688980957
transform 1 0 15640 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1006_
timestamp 1688980957
transform 1 0 15640 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1007_
timestamp 1688980957
transform 1 0 16100 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1008_
timestamp 1688980957
transform 1 0 14904 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _1009_
timestamp 1688980957
transform 1 0 15272 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1010_
timestamp 1688980957
transform 1 0 15088 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1011_
timestamp 1688980957
transform 1 0 14720 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1012_
timestamp 1688980957
transform 1 0 14076 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1013_
timestamp 1688980957
transform 1 0 14812 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1014_
timestamp 1688980957
transform 1 0 12972 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1688980957
transform 1 0 11868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1016_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1017_
timestamp 1688980957
transform 1 0 16468 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1018_
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1019_
timestamp 1688980957
transform 1 0 1840 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1020_
timestamp 1688980957
transform 1 0 7820 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1021_
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1022_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20608 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1023_
timestamp 1688980957
transform 1 0 6992 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1024_
timestamp 1688980957
transform 1 0 3128 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1025_
timestamp 1688980957
transform 1 0 5244 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1026_
timestamp 1688980957
transform 1 0 4692 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1027_
timestamp 1688980957
transform 1 0 3220 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1028_
timestamp 1688980957
transform 1 0 3680 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1029_
timestamp 1688980957
transform 1 0 4324 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1030_
timestamp 1688980957
transform 1 0 6900 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1031_
timestamp 1688980957
transform 1 0 7636 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1032_
timestamp 1688980957
transform 1 0 7912 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1033_
timestamp 1688980957
transform 1 0 10396 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1034_
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1035_
timestamp 1688980957
transform 1 0 10764 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1036_
timestamp 1688980957
transform 1 0 12512 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1037_
timestamp 1688980957
transform 1 0 13432 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1038_
timestamp 1688980957
transform 1 0 13432 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1039_
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1040_
timestamp 1688980957
transform 1 0 16744 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1041_
timestamp 1688980957
transform 1 0 16468 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1042_
timestamp 1688980957
transform 1 0 18952 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1043_
timestamp 1688980957
transform 1 0 19872 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1044_
timestamp 1688980957
transform 1 0 22448 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1045_
timestamp 1688980957
transform 1 0 22908 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1046_
timestamp 1688980957
transform 1 0 19872 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1047_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1048_
timestamp 1688980957
transform 1 0 20516 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1049_
timestamp 1688980957
transform 1 0 22448 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1050_
timestamp 1688980957
transform 1 0 24932 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1051_
timestamp 1688980957
transform 1 0 26220 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1052_
timestamp 1688980957
transform 1 0 24932 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1053_
timestamp 1688980957
transform 1 0 14444 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1054_
timestamp 1688980957
transform 1 0 1564 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1055_
timestamp 1688980957
transform 1 0 1748 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1056_
timestamp 1688980957
transform 1 0 13248 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1057_
timestamp 1688980957
transform 1 0 13524 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1058_
timestamp 1688980957
transform 1 0 13432 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1059_
timestamp 1688980957
transform 1 0 13432 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1060_
timestamp 1688980957
transform 1 0 22908 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1061_
timestamp 1688980957
transform 1 0 24472 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1062_
timestamp 1688980957
transform 1 0 26772 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1063_
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1064_
timestamp 1688980957
transform 1 0 23460 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1065_
timestamp 1688980957
transform 1 0 24472 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1066_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1067_
timestamp 1688980957
transform 1 0 8648 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1068_
timestamp 1688980957
transform 1 0 6164 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1069_
timestamp 1688980957
transform 1 0 20056 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1070_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1071_
timestamp 1688980957
transform 1 0 8464 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1072_
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1073_
timestamp 1688980957
transform 1 0 18768 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1074_
timestamp 1688980957
transform 1 0 18400 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1075_
timestamp 1688980957
transform 1 0 16376 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1076_
timestamp 1688980957
transform 1 0 14996 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1077_
timestamp 1688980957
transform 1 0 11592 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1078_
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1079_
timestamp 1688980957
transform 1 0 9568 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1080_
timestamp 1688980957
transform 1 0 9200 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1081_
timestamp 1688980957
transform 1 0 9016 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1082_
timestamp 1688980957
transform 1 0 1840 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1083_
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1084_
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1085_
timestamp 1688980957
transform 1 0 1840 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1086_
timestamp 1688980957
transform 1 0 2300 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1087_
timestamp 1688980957
transform 1 0 1656 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1088_
timestamp 1688980957
transform 1 0 9200 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1089_
timestamp 1688980957
transform 1 0 2116 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1090_
timestamp 1688980957
transform 1 0 9200 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1091_
timestamp 1688980957
transform 1 0 12144 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1092_
timestamp 1688980957
transform 1 0 12880 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1093_
timestamp 1688980957
transform 1 0 12144 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1094_
timestamp 1688980957
transform 1 0 4048 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1095_
timestamp 1688980957
transform 1 0 1840 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1096_
timestamp 1688980957
transform 1 0 7912 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1097_
timestamp 1688980957
transform 1 0 6624 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1098_
timestamp 1688980957
transform 1 0 1840 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1099_
timestamp 1688980957
transform 1 0 1932 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1100_
timestamp 1688980957
transform 1 0 12144 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1101_
timestamp 1688980957
transform 1 0 1840 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1102_
timestamp 1688980957
transform 1 0 12144 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1103_
timestamp 1688980957
transform 1 0 12144 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1104_
timestamp 1688980957
transform 1 0 10120 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1105_
timestamp 1688980957
transform 1 0 11776 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1106_
timestamp 1688980957
transform 1 0 5244 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1107_
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1108_
timestamp 1688980957
transform 1 0 6992 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1109_
timestamp 1688980957
transform 1 0 6532 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1110_
timestamp 1688980957
transform 1 0 5428 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1111_
timestamp 1688980957
transform 1 0 6256 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1112_
timestamp 1688980957
transform 1 0 12052 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1113_
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1114_
timestamp 1688980957
transform 1 0 11592 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1115_
timestamp 1688980957
transform 1 0 9568 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1116_
timestamp 1688980957
transform 1 0 9016 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1117_
timestamp 1688980957
transform 1 0 9292 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1118_
timestamp 1688980957
transform 1 0 3680 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1119_
timestamp 1688980957
transform 1 0 3772 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1120_
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1121_
timestamp 1688980957
transform 1 0 4232 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1122_
timestamp 1688980957
transform 1 0 5152 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1123_
timestamp 1688980957
transform 1 0 3864 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1124_
timestamp 1688980957
transform 1 0 9200 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1125_
timestamp 1688980957
transform 1 0 3956 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1126_
timestamp 1688980957
transform 1 0 9200 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1127_
timestamp 1688980957
transform 1 0 14720 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1128_
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1129_
timestamp 1688980957
transform 1 0 16560 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1130_
timestamp 1688980957
transform 1 0 17296 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1131_
timestamp 1688980957
transform 1 0 14168 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1132_
timestamp 1688980957
transform 1 0 17020 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1133_
timestamp 1688980957
transform 1 0 14352 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1134_
timestamp 1688980957
transform 1 0 16284 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1135_
timestamp 1688980957
transform 1 0 16560 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1136_
timestamp 1688980957
transform 1 0 14720 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1137_
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1138_
timestamp 1688980957
transform 1 0 14444 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1139_
timestamp 1688980957
transform 1 0 19872 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1140_
timestamp 1688980957
transform 1 0 18032 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1141_
timestamp 1688980957
transform 1 0 19964 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1142_
timestamp 1688980957
transform 1 0 22816 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2300 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk
timestamp 1688980957
transform 1 0 4876 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1688980957
transform 1 0 4600 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1688980957
transform 1 0 9936 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1688980957
transform 1 0 11040 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1688980957
transform 1 0 5244 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1688980957
transform 1 0 10396 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1688980957
transform 1 0 10856 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1688980957
transform 1 0 18216 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1688980957
transform 1 0 21988 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1688980957
transform 1 0 22632 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1688980957
transform 1 0 15364 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1688980957
transform 1 0 14536 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1688980957
transform 1 0 17388 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1688980957
transform 1 0 19596 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout35
timestamp 1688980957
transform 1 0 7820 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout36
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout37
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout38
timestamp 1688980957
transform 1 0 14628 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout39
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout40
timestamp 1688980957
transform 1 0 27968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout41
timestamp 1688980957
transform 1 0 24288 0 -1 29376
box -38 -48 866 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_35
timestamp 1688980957
transform 1 0 4324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_47 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1688980957
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_72
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_119
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_131
timestamp 1688980957
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_149
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_156
timestamp 1688980957
transform 1 0 15456 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_203
timestamp 1688980957
transform 1 0 19780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_215
timestamp 1688980957
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_225 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_233
timestamp 1688980957
transform 1 0 22540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_245
timestamp 1688980957
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_265 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_275
timestamp 1688980957
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 1688980957
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_293
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_147
timestamp 1688980957
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_159
timestamp 1688980957
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_187
timestamp 1688980957
transform 1 0 18308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_199
timestamp 1688980957
transform 1 0 19412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_211
timestamp 1688980957
transform 1 0 20516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_9
timestamp 1688980957
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_135
timestamp 1688980957
transform 1 0 13524 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_158
timestamp 1688980957
transform 1 0 15640 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_174
timestamp 1688980957
transform 1 0 17112 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_261
timestamp 1688980957
transform 1 0 25116 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_11
timestamp 1688980957
transform 1 0 2116 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_147
timestamp 1688980957
transform 1 0 14628 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_155
timestamp 1688980957
transform 1 0 15364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_166
timestamp 1688980957
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_184
timestamp 1688980957
transform 1 0 18032 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_188
timestamp 1688980957
transform 1 0 18400 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_209
timestamp 1688980957
transform 1 0 20332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_221
timestamp 1688980957
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_254
timestamp 1688980957
transform 1 0 24472 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_260
timestamp 1688980957
transform 1 0 25024 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_272
timestamp 1688980957
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_113
timestamp 1688980957
transform 1 0 11500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_125
timestamp 1688980957
transform 1 0 12604 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_134
timestamp 1688980957
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_187
timestamp 1688980957
transform 1 0 18308 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 1688980957
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_214
timestamp 1688980957
transform 1 0 20792 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_226
timestamp 1688980957
transform 1 0 21896 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_238
timestamp 1688980957
transform 1 0 23000 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_250
timestamp 1688980957
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_77
timestamp 1688980957
transform 1 0 8188 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 1688980957
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_134
timestamp 1688980957
transform 1 0 13432 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_146
timestamp 1688980957
transform 1 0 14536 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_158
timestamp 1688980957
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_166
timestamp 1688980957
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_197
timestamp 1688980957
transform 1 0 19228 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_211
timestamp 1688980957
transform 1 0 20516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_296
timestamp 1688980957
transform 1 0 28336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_304
timestamp 1688980957
transform 1 0 29072 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_51
timestamp 1688980957
transform 1 0 5796 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_55
timestamp 1688980957
transform 1 0 6164 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_76
timestamp 1688980957
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_117
timestamp 1688980957
transform 1 0 11868 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_129
timestamp 1688980957
transform 1 0 12972 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_137
timestamp 1688980957
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_50
timestamp 1688980957
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_65
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_84
timestamp 1688980957
transform 1 0 8832 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_119
timestamp 1688980957
transform 1 0 12052 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_131
timestamp 1688980957
transform 1 0 13156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_157
timestamp 1688980957
transform 1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_165
timestamp 1688980957
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_176
timestamp 1688980957
transform 1 0 17296 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_188
timestamp 1688980957
transform 1 0 18400 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_200
timestamp 1688980957
transform 1 0 19504 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_218
timestamp 1688980957
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_44
timestamp 1688980957
transform 1 0 5152 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_60
timestamp 1688980957
transform 1 0 6624 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_76
timestamp 1688980957
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_93
timestamp 1688980957
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_122
timestamp 1688980957
transform 1 0 12328 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_134
timestamp 1688980957
transform 1 0 13432 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_147
timestamp 1688980957
transform 1 0 14628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_159
timestamp 1688980957
transform 1 0 15732 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_185
timestamp 1688980957
transform 1 0 18124 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_193
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_231
timestamp 1688980957
transform 1 0 22356 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_256
timestamp 1688980957
transform 1 0 24656 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_268
timestamp 1688980957
transform 1 0 25760 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_280
timestamp 1688980957
transform 1 0 26864 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_292
timestamp 1688980957
transform 1 0 27968 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_304
timestamp 1688980957
transform 1 0 29072 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_47
timestamp 1688980957
transform 1 0 5428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_99
timestamp 1688980957
transform 1 0 10212 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_122
timestamp 1688980957
transform 1 0 12328 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_128
timestamp 1688980957
transform 1 0 12880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_158
timestamp 1688980957
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1688980957
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_189
timestamp 1688980957
transform 1 0 18492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_201
timestamp 1688980957
transform 1 0 19596 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_213
timestamp 1688980957
transform 1 0 20700 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_221
timestamp 1688980957
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_257
timestamp 1688980957
transform 1 0 24748 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_290
timestamp 1688980957
transform 1 0 27784 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_298
timestamp 1688980957
transform 1 0 28520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1688980957
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_45
timestamp 1688980957
transform 1 0 5244 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_70
timestamp 1688980957
transform 1 0 7544 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1688980957
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_149
timestamp 1688980957
transform 1 0 14812 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_161
timestamp 1688980957
transform 1 0 15916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_190
timestamp 1688980957
transform 1 0 18584 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_205
timestamp 1688980957
transform 1 0 19964 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_250
timestamp 1688980957
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_263
timestamp 1688980957
transform 1 0 25300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_274
timestamp 1688980957
transform 1 0 26312 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_291
timestamp 1688980957
transform 1 0 27876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_303
timestamp 1688980957
transform 1 0 28980 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_38
timestamp 1688980957
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_64
timestamp 1688980957
transform 1 0 6992 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_75
timestamp 1688980957
transform 1 0 8004 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_87
timestamp 1688980957
transform 1 0 9108 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_99
timestamp 1688980957
transform 1 0 10212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_129
timestamp 1688980957
transform 1 0 12972 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_157
timestamp 1688980957
transform 1 0 15548 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_165
timestamp 1688980957
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_183
timestamp 1688980957
transform 1 0 17940 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_191
timestamp 1688980957
transform 1 0 18676 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_213
timestamp 1688980957
transform 1 0 20700 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_218
timestamp 1688980957
transform 1 0 21160 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_233
timestamp 1688980957
transform 1 0 22540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_241
timestamp 1688980957
transform 1 0 23276 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_251
timestamp 1688980957
transform 1 0 24196 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_263
timestamp 1688980957
transform 1 0 25300 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_291
timestamp 1688980957
transform 1 0 27876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_303
timestamp 1688980957
transform 1 0 28980 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_7
timestamp 1688980957
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_33
timestamp 1688980957
transform 1 0 4140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_42
timestamp 1688980957
transform 1 0 4968 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_76
timestamp 1688980957
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_120
timestamp 1688980957
transform 1 0 12144 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_128
timestamp 1688980957
transform 1 0 12880 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_132
timestamp 1688980957
transform 1 0 13248 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_145
timestamp 1688980957
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_154
timestamp 1688980957
transform 1 0 15272 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_166
timestamp 1688980957
transform 1 0 16376 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_178
timestamp 1688980957
transform 1 0 17480 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_182
timestamp 1688980957
transform 1 0 17848 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_190
timestamp 1688980957
transform 1 0 18584 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_205
timestamp 1688980957
transform 1 0 19964 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_217
timestamp 1688980957
transform 1 0 21068 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_223
timestamp 1688980957
transform 1 0 21620 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_239
timestamp 1688980957
transform 1 0 23092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_299
timestamp 1688980957
transform 1 0 28612 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_50
timestamp 1688980957
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_67
timestamp 1688980957
transform 1 0 7268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_79
timestamp 1688980957
transform 1 0 8372 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_155
timestamp 1688980957
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_176
timestamp 1688980957
transform 1 0 17296 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_195
timestamp 1688980957
transform 1 0 19044 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_207
timestamp 1688980957
transform 1 0 20148 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_219
timestamp 1688980957
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_278
timestamp 1688980957
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_296
timestamp 1688980957
transform 1 0 28336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_304
timestamp 1688980957
transform 1 0 29072 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_40
timestamp 1688980957
transform 1 0 4784 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_52
timestamp 1688980957
transform 1 0 5888 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_64
timestamp 1688980957
transform 1 0 6992 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_76
timestamp 1688980957
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_113
timestamp 1688980957
transform 1 0 11500 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1688980957
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_144
timestamp 1688980957
transform 1 0 14352 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_152
timestamp 1688980957
transform 1 0 15088 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_163
timestamp 1688980957
transform 1 0 16100 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_167
timestamp 1688980957
transform 1 0 16468 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_215
timestamp 1688980957
transform 1 0 20884 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_227
timestamp 1688980957
transform 1 0 21988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_233
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_242
timestamp 1688980957
transform 1 0 23368 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_250
timestamp 1688980957
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_273
timestamp 1688980957
transform 1 0 26220 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_285
timestamp 1688980957
transform 1 0 27324 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_297
timestamp 1688980957
transform 1 0 28428 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_36
timestamp 1688980957
transform 1 0 4416 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_45
timestamp 1688980957
transform 1 0 5244 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_63
timestamp 1688980957
transform 1 0 6900 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_75
timestamp 1688980957
transform 1 0 8004 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_87
timestamp 1688980957
transform 1 0 9108 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_133
timestamp 1688980957
transform 1 0 13340 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_188
timestamp 1688980957
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_222
timestamp 1688980957
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_259
timestamp 1688980957
transform 1 0 24932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_263
timestamp 1688980957
transform 1 0 25300 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_7
timestamp 1688980957
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_44
timestamp 1688980957
transform 1 0 5152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_74
timestamp 1688980957
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1688980957
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_93
timestamp 1688980957
transform 1 0 9660 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_107
timestamp 1688980957
transform 1 0 10948 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_119
timestamp 1688980957
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_131
timestamp 1688980957
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_157
timestamp 1688980957
transform 1 0 15548 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_185
timestamp 1688980957
transform 1 0 18124 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_288
timestamp 1688980957
transform 1 0 27600 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_296
timestamp 1688980957
transform 1 0 28336 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_9
timestamp 1688980957
transform 1 0 1932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_52
timestamp 1688980957
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_67
timestamp 1688980957
transform 1 0 7268 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_78
timestamp 1688980957
transform 1 0 8280 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1688980957
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_144
timestamp 1688980957
transform 1 0 14352 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_156
timestamp 1688980957
transform 1 0 15456 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_160
timestamp 1688980957
transform 1 0 15824 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_180
timestamp 1688980957
transform 1 0 17664 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_186
timestamp 1688980957
transform 1 0 18216 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_218
timestamp 1688980957
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_255
timestamp 1688980957
transform 1 0 24564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_263
timestamp 1688980957
transform 1 0 25300 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_272
timestamp 1688980957
transform 1 0 26128 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_33
timestamp 1688980957
transform 1 0 4140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_75
timestamp 1688980957
transform 1 0 8004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_119
timestamp 1688980957
transform 1 0 12052 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_156
timestamp 1688980957
transform 1 0 15456 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_160
timestamp 1688980957
transform 1 0 15824 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_174
timestamp 1688980957
transform 1 0 17112 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_186
timestamp 1688980957
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1688980957
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_206
timestamp 1688980957
transform 1 0 20056 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_218
timestamp 1688980957
transform 1 0 21160 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_230
timestamp 1688980957
transform 1 0 22264 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1688980957
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1688980957
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1688980957
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_301
timestamp 1688980957
transform 1 0 28796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_35
timestamp 1688980957
transform 1 0 4324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_76
timestamp 1688980957
transform 1 0 8096 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_108
timestamp 1688980957
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_128
timestamp 1688980957
transform 1 0 12880 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_132
timestamp 1688980957
transform 1 0 13248 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_176
timestamp 1688980957
transform 1 0 17296 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_207
timestamp 1688980957
transform 1 0 20148 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_215
timestamp 1688980957
transform 1 0 20884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_243
timestamp 1688980957
transform 1 0 23460 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_255
timestamp 1688980957
transform 1 0 24564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_267
timestamp 1688980957
transform 1 0 25668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1688980957
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_11
timestamp 1688980957
transform 1 0 2116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_66
timestamp 1688980957
transform 1 0 7176 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1688980957
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_100
timestamp 1688980957
transform 1 0 10304 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_120
timestamp 1688980957
transform 1 0 12144 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_132
timestamp 1688980957
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_189
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_203
timestamp 1688980957
transform 1 0 19780 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_215
timestamp 1688980957
transform 1 0 20884 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_223
timestamp 1688980957
transform 1 0 21620 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_227
timestamp 1688980957
transform 1 0 21988 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_247
timestamp 1688980957
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1688980957
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_269
timestamp 1688980957
transform 1 0 25852 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_281
timestamp 1688980957
transform 1 0 26956 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_293
timestamp 1688980957
transform 1 0 28060 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_28
timestamp 1688980957
transform 1 0 3680 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_40
timestamp 1688980957
transform 1 0 4784 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_52
timestamp 1688980957
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_64
timestamp 1688980957
transform 1 0 6992 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_76
timestamp 1688980957
transform 1 0 8096 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_88
timestamp 1688980957
transform 1 0 9200 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_94
timestamp 1688980957
transform 1 0 9752 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_102
timestamp 1688980957
transform 1 0 10488 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_146
timestamp 1688980957
transform 1 0 14536 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_157
timestamp 1688980957
transform 1 0 15548 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_165
timestamp 1688980957
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_187
timestamp 1688980957
transform 1 0 18308 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_212
timestamp 1688980957
transform 1 0 20608 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_216
timestamp 1688980957
transform 1 0 20976 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_233
timestamp 1688980957
transform 1 0 22540 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_253
timestamp 1688980957
transform 1 0 24380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_274
timestamp 1688980957
transform 1 0 26312 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_289
timestamp 1688980957
transform 1 0 27692 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_304
timestamp 1688980957
transform 1 0 29072 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_72
timestamp 1688980957
transform 1 0 7728 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_113
timestamp 1688980957
transform 1 0 11500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_134
timestamp 1688980957
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_150
timestamp 1688980957
transform 1 0 14904 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_171
timestamp 1688980957
transform 1 0 16836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_183
timestamp 1688980957
transform 1 0 17940 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1688980957
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_216
timestamp 1688980957
transform 1 0 20976 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_240
timestamp 1688980957
transform 1 0 23184 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp 1688980957
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_277
timestamp 1688980957
transform 1 0 26588 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_302
timestamp 1688980957
transform 1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_31
timestamp 1688980957
transform 1 0 3956 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_52
timestamp 1688980957
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_87
timestamp 1688980957
transform 1 0 9108 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_108
timestamp 1688980957
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_140
timestamp 1688980957
transform 1 0 13984 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_144
timestamp 1688980957
transform 1 0 14352 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_203
timestamp 1688980957
transform 1 0 19780 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_234
timestamp 1688980957
transform 1 0 22632 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_250
timestamp 1688980957
transform 1 0 24104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_262
timestamp 1688980957
transform 1 0 25208 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_277
timestamp 1688980957
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1688980957
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_7
timestamp 1688980957
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_33
timestamp 1688980957
transform 1 0 4140 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_54
timestamp 1688980957
transform 1 0 6072 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_80
timestamp 1688980957
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_108
timestamp 1688980957
transform 1 0 11040 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_116
timestamp 1688980957
transform 1 0 11776 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_164
timestamp 1688980957
transform 1 0 16192 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 1688980957
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_208
timestamp 1688980957
transform 1 0 20240 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_220
timestamp 1688980957
transform 1 0 21344 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_232
timestamp 1688980957
transform 1 0 22448 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_238
timestamp 1688980957
transform 1 0 23000 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_265
timestamp 1688980957
transform 1 0 25484 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_287
timestamp 1688980957
transform 1 0 27508 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_299
timestamp 1688980957
transform 1 0 28612 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_6
timestamp 1688980957
transform 1 0 1656 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_14
timestamp 1688980957
transform 1 0 2392 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_43
timestamp 1688980957
transform 1 0 5060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_47
timestamp 1688980957
transform 1 0 5428 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_72
timestamp 1688980957
transform 1 0 7728 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_90
timestamp 1688980957
transform 1 0 9384 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_94
timestamp 1688980957
transform 1 0 9752 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 1688980957
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_121
timestamp 1688980957
transform 1 0 12236 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_136
timestamp 1688980957
transform 1 0 13616 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_148
timestamp 1688980957
transform 1 0 14720 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_166
timestamp 1688980957
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1688980957
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1688980957
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1688980957
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1688980957
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_237
timestamp 1688980957
transform 1 0 22908 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_246
timestamp 1688980957
transform 1 0 23736 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_258
timestamp 1688980957
transform 1 0 24840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_266
timestamp 1688980957
transform 1 0 25576 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_270
timestamp 1688980957
transform 1 0 25944 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_278
timestamp 1688980957
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1688980957
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_23
timestamp 1688980957
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_37
timestamp 1688980957
transform 1 0 4508 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_57
timestamp 1688980957
transform 1 0 6348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_69
timestamp 1688980957
transform 1 0 7452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_81
timestamp 1688980957
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_93
timestamp 1688980957
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_102
timestamp 1688980957
transform 1 0 10488 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_111
timestamp 1688980957
transform 1 0 11316 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_123
timestamp 1688980957
transform 1 0 12420 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_135
timestamp 1688980957
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_148
timestamp 1688980957
transform 1 0 14720 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_157
timestamp 1688980957
transform 1 0 15548 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_169
timestamp 1688980957
transform 1 0 16652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_181
timestamp 1688980957
transform 1 0 17756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1688980957
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_221
timestamp 1688980957
transform 1 0 21436 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_233
timestamp 1688980957
transform 1 0 22540 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_248
timestamp 1688980957
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_262
timestamp 1688980957
transform 1 0 25208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_268
timestamp 1688980957
transform 1 0 25760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_283
timestamp 1688980957
transform 1 0 27140 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_297
timestamp 1688980957
transform 1 0 28428 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_23
timestamp 1688980957
transform 1 0 3220 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_52
timestamp 1688980957
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_89
timestamp 1688980957
transform 1 0 9292 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_119
timestamp 1688980957
transform 1 0 12052 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_148
timestamp 1688980957
transform 1 0 14720 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_158
timestamp 1688980957
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1688980957
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_177
timestamp 1688980957
transform 1 0 17388 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_198
timestamp 1688980957
transform 1 0 19320 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_210
timestamp 1688980957
transform 1 0 20424 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_234
timestamp 1688980957
transform 1 0 22632 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_300
timestamp 1688980957
transform 1 0 28704 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_304
timestamp 1688980957
transform 1 0 29072 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_43
timestamp 1688980957
transform 1 0 5060 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_72
timestamp 1688980957
transform 1 0 7728 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_91
timestamp 1688980957
transform 1 0 9476 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_170
timestamp 1688980957
transform 1 0 16744 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_204
timestamp 1688980957
transform 1 0 19872 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_227
timestamp 1688980957
transform 1 0 21988 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_239
timestamp 1688980957
transform 1 0 23092 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_249
timestamp 1688980957
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_284
timestamp 1688980957
transform 1 0 27232 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_297
timestamp 1688980957
transform 1 0 28428 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_7
timestamp 1688980957
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_48
timestamp 1688980957
transform 1 0 5520 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_78
timestamp 1688980957
transform 1 0 8280 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_121
timestamp 1688980957
transform 1 0 12236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_141
timestamp 1688980957
transform 1 0 14076 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_147
timestamp 1688980957
transform 1 0 14628 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_193
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_218
timestamp 1688980957
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_268
timestamp 1688980957
transform 1 0 25760 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_304
timestamp 1688980957
transform 1 0 29072 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_40
timestamp 1688980957
transform 1 0 4784 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_52
timestamp 1688980957
transform 1 0 5888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_62
timestamp 1688980957
transform 1 0 6808 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_93
timestamp 1688980957
transform 1 0 9660 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_118
timestamp 1688980957
transform 1 0 11960 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_128
timestamp 1688980957
transform 1 0 12880 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_171
timestamp 1688980957
transform 1 0 16836 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_184
timestamp 1688980957
transform 1 0 18032 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1688980957
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1688980957
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1688980957
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1688980957
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_9
timestamp 1688980957
transform 1 0 1932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_21
timestamp 1688980957
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_33
timestamp 1688980957
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_45
timestamp 1688980957
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_53
timestamp 1688980957
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_65
timestamp 1688980957
transform 1 0 7084 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_94
timestamp 1688980957
transform 1 0 9752 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_106
timestamp 1688980957
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_121
timestamp 1688980957
transform 1 0 12236 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_134
timestamp 1688980957
transform 1 0 13432 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_146
timestamp 1688980957
transform 1 0 14536 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_157
timestamp 1688980957
transform 1 0 15548 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1688980957
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_176
timestamp 1688980957
transform 1 0 17296 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_188
timestamp 1688980957
transform 1 0 18400 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_212
timestamp 1688980957
transform 1 0 20608 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1688980957
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1688980957
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1688980957
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_285
timestamp 1688980957
transform 1 0 27324 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_291
timestamp 1688980957
transform 1 0 27876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_303
timestamp 1688980957
transform 1 0 28980 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_7
timestamp 1688980957
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_37
timestamp 1688980957
transform 1 0 4508 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_49
timestamp 1688980957
transform 1 0 5612 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_72
timestamp 1688980957
transform 1 0 7728 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_93
timestamp 1688980957
transform 1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_110
timestamp 1688980957
transform 1 0 11224 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_118
timestamp 1688980957
transform 1 0 11960 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_126
timestamp 1688980957
transform 1 0 12696 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_136
timestamp 1688980957
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_153
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_164
timestamp 1688980957
transform 1 0 16192 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_176
timestamp 1688980957
transform 1 0 17296 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_188
timestamp 1688980957
transform 1 0 18400 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1688980957
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1688980957
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1688980957
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1688980957
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1688980957
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_277
timestamp 1688980957
transform 1 0 26588 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_281
timestamp 1688980957
transform 1 0 26956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_297
timestamp 1688980957
transform 1 0 28428 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_23
timestamp 1688980957
transform 1 0 3220 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_40
timestamp 1688980957
transform 1 0 4784 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_52
timestamp 1688980957
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_85
timestamp 1688980957
transform 1 0 8924 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_107
timestamp 1688980957
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_151
timestamp 1688980957
transform 1 0 14996 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_163
timestamp 1688980957
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_189
timestamp 1688980957
transform 1 0 18492 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_203
timestamp 1688980957
transform 1 0 19780 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_215
timestamp 1688980957
transform 1 0 20884 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_230
timestamp 1688980957
transform 1 0 22264 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_234
timestamp 1688980957
transform 1 0 22632 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_240
timestamp 1688980957
transform 1 0 23184 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_253
timestamp 1688980957
transform 1 0 24380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_265
timestamp 1688980957
transform 1 0 25484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_303
timestamp 1688980957
transform 1 0 28980 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_49
timestamp 1688980957
transform 1 0 5612 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_61
timestamp 1688980957
transform 1 0 6716 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_75
timestamp 1688980957
transform 1 0 8004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_99
timestamp 1688980957
transform 1 0 10212 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_157
timestamp 1688980957
transform 1 0 15548 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_224
timestamp 1688980957
transform 1 0 21712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_249
timestamp 1688980957
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_273
timestamp 1688980957
transform 1 0 26220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_300
timestamp 1688980957
transform 1 0 28704 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_304
timestamp 1688980957
transform 1 0 29072 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_21
timestamp 1688980957
transform 1 0 3036 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_84
timestamp 1688980957
transform 1 0 8832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_106
timestamp 1688980957
transform 1 0 10856 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_127
timestamp 1688980957
transform 1 0 12788 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_148
timestamp 1688980957
transform 1 0 14720 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_160
timestamp 1688980957
transform 1 0 15824 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_201
timestamp 1688980957
transform 1 0 19596 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_266
timestamp 1688980957
transform 1 0 25576 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_278
timestamp 1688980957
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_284
timestamp 1688980957
transform 1 0 27232 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_290
timestamp 1688980957
transform 1 0 27784 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_302
timestamp 1688980957
transform 1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_40
timestamp 1688980957
transform 1 0 4784 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_44
timestamp 1688980957
transform 1 0 5152 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_81
timestamp 1688980957
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1688980957
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_165
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_173
timestamp 1688980957
transform 1 0 17020 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_183
timestamp 1688980957
transform 1 0 17940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_205
timestamp 1688980957
transform 1 0 19964 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_215
timestamp 1688980957
transform 1 0 20884 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_271
timestamp 1688980957
transform 1 0 26036 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_283
timestamp 1688980957
transform 1 0 27140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_295
timestamp 1688980957
transform 1 0 28244 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_303
timestamp 1688980957
transform 1 0 28980 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_35
timestamp 1688980957
transform 1 0 4324 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_44
timestamp 1688980957
transform 1 0 5152 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_68
timestamp 1688980957
transform 1 0 7360 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_78
timestamp 1688980957
transform 1 0 8280 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_109
timestamp 1688980957
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_128
timestamp 1688980957
transform 1 0 12880 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_140
timestamp 1688980957
transform 1 0 13984 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_148
timestamp 1688980957
transform 1 0 14720 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_166
timestamp 1688980957
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_177
timestamp 1688980957
transform 1 0 17388 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_189
timestamp 1688980957
transform 1 0 18492 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_201
timestamp 1688980957
transform 1 0 19596 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_209
timestamp 1688980957
transform 1 0 20332 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_216
timestamp 1688980957
transform 1 0 20976 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_228
timestamp 1688980957
transform 1 0 22080 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_234
timestamp 1688980957
transform 1 0 22632 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_238
timestamp 1688980957
transform 1 0 23000 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_242
timestamp 1688980957
transform 1 0 23368 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_265
timestamp 1688980957
transform 1 0 25484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_277
timestamp 1688980957
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_293
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_35
timestamp 1688980957
transform 1 0 4324 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_44
timestamp 1688980957
transform 1 0 5152 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_52
timestamp 1688980957
transform 1 0 5888 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_64
timestamp 1688980957
transform 1 0 6992 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_76
timestamp 1688980957
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_117
timestamp 1688980957
transform 1 0 11868 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_129
timestamp 1688980957
transform 1 0 12972 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_137
timestamp 1688980957
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_163
timestamp 1688980957
transform 1 0 16100 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_175
timestamp 1688980957
transform 1 0 17204 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_182
timestamp 1688980957
transform 1 0 17848 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 1688980957
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_220
timestamp 1688980957
transform 1 0 21344 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_232
timestamp 1688980957
transform 1 0 22448 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_244
timestamp 1688980957
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_263
timestamp 1688980957
transform 1 0 25300 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_275
timestamp 1688980957
transform 1 0 26404 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_287
timestamp 1688980957
transform 1 0 27508 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_299
timestamp 1688980957
transform 1 0 28612 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_9
timestamp 1688980957
transform 1 0 1932 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_21
timestamp 1688980957
transform 1 0 3036 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_33
timestamp 1688980957
transform 1 0 4140 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_45
timestamp 1688980957
transform 1 0 5244 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_53
timestamp 1688980957
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_87
timestamp 1688980957
transform 1 0 9108 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_108
timestamp 1688980957
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_121
timestamp 1688980957
transform 1 0 12236 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_138
timestamp 1688980957
transform 1 0 13800 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_164
timestamp 1688980957
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_186
timestamp 1688980957
transform 1 0 18216 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_198
timestamp 1688980957
transform 1 0 19320 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_210
timestamp 1688980957
transform 1 0 20424 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_222
timestamp 1688980957
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 1688980957
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 1688980957
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 1688980957
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 1688980957
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1688980957
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_35
timestamp 1688980957
transform 1 0 4324 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_43
timestamp 1688980957
transform 1 0 5060 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_68
timestamp 1688980957
transform 1 0 7360 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_80
timestamp 1688980957
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_93
timestamp 1688980957
transform 1 0 9660 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_104
timestamp 1688980957
transform 1 0 10672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_112
timestamp 1688980957
transform 1 0 11408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_137
timestamp 1688980957
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_145
timestamp 1688980957
transform 1 0 14444 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_157
timestamp 1688980957
transform 1 0 15548 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 1688980957
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_207
timestamp 1688980957
transform 1 0 20148 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_219
timestamp 1688980957
transform 1 0 21252 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_231
timestamp 1688980957
transform 1 0 22356 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_243
timestamp 1688980957
transform 1 0 23460 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1688980957
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 1688980957
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 1688980957
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_301
timestamp 1688980957
transform 1 0 28796 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_21
timestamp 1688980957
transform 1 0 3036 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_47
timestamp 1688980957
transform 1 0 5428 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_72
timestamp 1688980957
transform 1 0 7728 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_100
timestamp 1688980957
transform 1 0 10304 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_136
timestamp 1688980957
transform 1 0 13616 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_148
timestamp 1688980957
transform 1 0 14720 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_166
timestamp 1688980957
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_174
timestamp 1688980957
transform 1 0 17112 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_220
timestamp 1688980957
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1688980957
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_7
timestamp 1688980957
transform 1 0 1748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_35
timestamp 1688980957
transform 1 0 4324 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_109
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_120
timestamp 1688980957
transform 1 0 12144 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_132
timestamp 1688980957
transform 1 0 13248 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_149
timestamp 1688980957
transform 1 0 14812 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_235
timestamp 1688980957
transform 1 0 22724 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_247
timestamp 1688980957
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 1688980957
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 1688980957
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_301
timestamp 1688980957
transform 1 0 28796 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_80
timestamp 1688980957
transform 1 0 8464 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_92
timestamp 1688980957
transform 1 0 9568 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_104
timestamp 1688980957
transform 1 0 10672 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_189
timestamp 1688980957
transform 1 0 18492 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_212
timestamp 1688980957
transform 1 0 20608 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1688980957
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 1688980957
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_11
timestamp 1688980957
transform 1 0 2116 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_49
timestamp 1688980957
transform 1 0 5612 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_63
timestamp 1688980957
transform 1 0 6900 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_75
timestamp 1688980957
transform 1 0 8004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_125
timestamp 1688980957
transform 1 0 12604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_137
timestamp 1688980957
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1688980957
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 1688980957
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1688980957
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_202
timestamp 1688980957
transform 1 0 19688 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_214
timestamp 1688980957
transform 1 0 20792 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_226
timestamp 1688980957
transform 1 0 21896 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_238
timestamp 1688980957
transform 1 0 23000 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_250
timestamp 1688980957
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 1688980957
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_301
timestamp 1688980957
transform 1 0 28796 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_73
timestamp 1688980957
transform 1 0 7820 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_94
timestamp 1688980957
transform 1 0 9752 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_106
timestamp 1688980957
transform 1 0 10856 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_119
timestamp 1688980957
transform 1 0 12052 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_123
timestamp 1688980957
transform 1 0 12420 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_148
timestamp 1688980957
transform 1 0 14720 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_160
timestamp 1688980957
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_173
timestamp 1688980957
transform 1 0 17020 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_180
timestamp 1688980957
transform 1 0 17664 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_192
timestamp 1688980957
transform 1 0 18768 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_204
timestamp 1688980957
transform 1 0 19872 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_212
timestamp 1688980957
transform 1 0 20608 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_219
timestamp 1688980957
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1688980957
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1688980957
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1688980957
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_293
timestamp 1688980957
transform 1 0 28060 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_9
timestamp 1688980957
transform 1 0 1932 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_25
timestamp 1688980957
transform 1 0 3404 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_33
timestamp 1688980957
transform 1 0 4140 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_42
timestamp 1688980957
transform 1 0 4968 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_54
timestamp 1688980957
transform 1 0 6072 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_66
timestamp 1688980957
transform 1 0 7176 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_77
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_91
timestamp 1688980957
transform 1 0 9476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_103
timestamp 1688980957
transform 1 0 10580 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_121
timestamp 1688980957
transform 1 0 12236 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_130
timestamp 1688980957
transform 1 0 13064 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_150
timestamp 1688980957
transform 1 0 14904 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_162
timestamp 1688980957
transform 1 0 16008 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_187
timestamp 1688980957
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1688980957
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_201
timestamp 1688980957
transform 1 0 19596 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_228
timestamp 1688980957
transform 1 0 22080 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_237
timestamp 1688980957
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 1688980957
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1688980957
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 1688980957
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_301
timestamp 1688980957
transform 1 0 28796 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_23
timestamp 1688980957
transform 1 0 3220 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_54
timestamp 1688980957
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_68
timestamp 1688980957
transform 1 0 7360 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_96
timestamp 1688980957
transform 1 0 9936 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_120
timestamp 1688980957
transform 1 0 12144 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_128
timestamp 1688980957
transform 1 0 12880 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_165
timestamp 1688980957
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_191
timestamp 1688980957
transform 1 0 18676 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_222
timestamp 1688980957
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_257
timestamp 1688980957
transform 1 0 24748 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_269
timestamp 1688980957
transform 1 0 25852 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_277
timestamp 1688980957
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_62
timestamp 1688980957
transform 1 0 6808 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_95
timestamp 1688980957
transform 1 0 9844 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_126
timestamp 1688980957
transform 1 0 12696 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_130
timestamp 1688980957
transform 1 0 13064 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_149
timestamp 1688980957
transform 1 0 14812 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_161
timestamp 1688980957
transform 1 0 15916 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_190
timestamp 1688980957
transform 1 0 18584 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_201
timestamp 1688980957
transform 1 0 19596 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_270
timestamp 1688980957
transform 1 0 25944 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_282
timestamp 1688980957
transform 1 0 27048 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_294
timestamp 1688980957
transform 1 0 28152 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_302
timestamp 1688980957
transform 1 0 28888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_87
timestamp 1688980957
transform 1 0 9108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_99
timestamp 1688980957
transform 1 0 10212 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_133
timestamp 1688980957
transform 1 0 13340 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_162
timestamp 1688980957
transform 1 0 16008 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_197
timestamp 1688980957
transform 1 0 19228 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_203
timestamp 1688980957
transform 1 0 19780 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_231
timestamp 1688980957
transform 1 0 22356 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_250
timestamp 1688980957
transform 1 0 24104 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 1688980957
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 1688980957
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1688980957
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1688980957
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_44
timestamp 1688980957
transform 1 0 5152 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_52
timestamp 1688980957
transform 1 0 5888 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_64
timestamp 1688980957
transform 1 0 6992 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_73
timestamp 1688980957
transform 1 0 7820 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_81
timestamp 1688980957
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_94
timestamp 1688980957
transform 1 0 9752 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_106
timestamp 1688980957
transform 1 0 10856 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_117
timestamp 1688980957
transform 1 0 11868 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_129
timestamp 1688980957
transform 1 0 12972 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_137
timestamp 1688980957
transform 1 0 13708 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_156
timestamp 1688980957
transform 1 0 15456 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_168
timestamp 1688980957
transform 1 0 16560 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_179
timestamp 1688980957
transform 1 0 17572 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_191
timestamp 1688980957
transform 1 0 18676 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1688980957
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_215
timestamp 1688980957
transform 1 0 20884 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_227
timestamp 1688980957
transform 1 0 21988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_239
timestamp 1688980957
transform 1 0 23092 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_248
timestamp 1688980957
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1688980957
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1688980957
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_301
timestamp 1688980957
transform 1 0 28796 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_6
timestamp 1688980957
transform 1 0 1656 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_14
timestamp 1688980957
transform 1 0 2392 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_23
timestamp 1688980957
transform 1 0 3220 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_29
timestamp 1688980957
transform 1 0 3772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_41
timestamp 1688980957
transform 1 0 4876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_53
timestamp 1688980957
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_65
timestamp 1688980957
transform 1 0 7084 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_77
timestamp 1688980957
transform 1 0 8188 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_83
timestamp 1688980957
transform 1 0 8740 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_85
timestamp 1688980957
transform 1 0 8924 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_100
timestamp 1688980957
transform 1 0 10304 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_147
timestamp 1688980957
transform 1 0 14628 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_159
timestamp 1688980957
transform 1 0 15732 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_177
timestamp 1688980957
transform 1 0 17388 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_184
timestamp 1688980957
transform 1 0 18032 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_197
timestamp 1688980957
transform 1 0 19228 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_209
timestamp 1688980957
transform 1 0 20332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_221
timestamp 1688980957
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_231
timestamp 1688980957
transform 1 0 22356 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_243
timestamp 1688980957
transform 1 0 23460 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_251
timestamp 1688980957
transform 1 0 24196 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_253
timestamp 1688980957
transform 1 0 24380 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_261
timestamp 1688980957
transform 1 0 25116 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_268
timestamp 1688980957
transform 1 0 25760 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 2668 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 10488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 17480 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 16192 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 16928 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 13248 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 7544 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 14996 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 16008 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 6440 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform 1 0 14812 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 8188 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 12512 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform 1 0 4048 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 13340 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform 1 0 5244 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform 1 0 8648 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform 1 0 7544 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform 1 0 13616 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform 1 0 7544 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform 1 0 14996 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 4416 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 13340 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform 1 0 4324 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform 1 0 4140 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 8096 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform 1 0 12880 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform 1 0 9476 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform 1 0 17204 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform 1 0 4232 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform 1 0 4416 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform 1 0 4324 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform 1 0 5612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 9936 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform 1 0 7820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform 1 0 4048 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform 1 0 5244 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform 1 0 4416 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform 1 0 10580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform 1 0 9660 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 20792 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform 1 0 15272 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform 1 0 15272 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform 1 0 3864 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform 1 0 4324 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform 1 0 9568 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform 1 0 18492 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform 1 0 25116 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform 1 0 9108 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform 1 0 8096 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform 1 0 6164 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform 1 0 5060 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform 1 0 23368 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform 1 0 25208 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform 1 0 5520 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform 1 0 26496 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform 1 0 14536 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform 1 0 25392 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform 1 0 26864 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform 1 0 10396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform 1 0 23092 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform 1 0 25024 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1688980957
transform 1 0 28336 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap33
timestamp 1688980957
transform 1 0 8280 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  max_cap34
timestamp 1688980957
transform 1 0 19412 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output4
timestamp 1688980957
transform 1 0 14904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output5
timestamp 1688980957
transform 1 0 9752 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output6
timestamp 1688980957
transform -1 0 1932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output7
timestamp 1688980957
transform 1 0 28612 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output8
timestamp 1688980957
transform 1 0 17480 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 1688980957
transform 1 0 28612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1688980957
transform 1 0 28796 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 1688980957
transform 1 0 25852 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1688980957
transform 1 0 28796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1688980957
transform 1 0 25208 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1688980957
transform 1 0 6532 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1688980957
transform 1 0 21988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1688980957
transform 1 0 28796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1688980957
transform 1 0 2668 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1688980957
transform 1 0 28612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1688980957
transform 1 0 28796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1688980957
transform 1 0 28612 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1688980957
transform 1 0 14076 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1688980957
transform 1 0 28796 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 29440 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 29440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 29440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 29440 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 29440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 29440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 29440 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 29440 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 29440 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 29440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 29440 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 29440 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 29440 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 29440 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 29440 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 29440 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 29440 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 29440 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 29440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 29440 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 29440 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 29440 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 29440 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 29440 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 29440 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 29440 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 29440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 29440 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 29440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 29440 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 29440 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 29440 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 29440 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 29440 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 29440 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 29440 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 29440 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 29440 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 29440 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 29440 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 29440 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 29440 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 29440 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 29440 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 29440 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 29440 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 29440 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 29440 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 29440 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 29440 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 29440 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 29440 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 3680 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 8832 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 13984 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 19136 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 24288 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 28998 31925 29054 32725 0 FreeSans 224 90 0 0 nrst
port 1 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 out_0[0]
port 2 nsew signal tristate
flabel metal2 s 9678 31925 9734 32725 0 FreeSans 224 90 0 0 out_0[1]
port 3 nsew signal tristate
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 out_0[2]
port 4 nsew signal tristate
flabel metal3 s 29781 10888 30581 11008 0 FreeSans 480 0 0 0 out_0[3]
port 5 nsew signal tristate
flabel metal2 s 17406 31925 17462 32725 0 FreeSans 224 90 0 0 out_0[4]
port 6 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 out_0[5]
port 7 nsew signal tristate
flabel metal3 s 29781 18368 30581 18488 0 FreeSans 480 0 0 0 out_0[6]
port 8 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 out_1[0]
port 9 nsew signal tristate
flabel metal3 s 29781 22448 30581 22568 0 FreeSans 480 0 0 0 out_1[1]
port 10 nsew signal tristate
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 out_1[2]
port 11 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 out_1[3]
port 12 nsew signal tristate
flabel metal2 s 21270 31925 21326 32725 0 FreeSans 224 90 0 0 out_1[4]
port 13 nsew signal tristate
flabel metal2 s 25134 31925 25190 32725 0 FreeSans 224 90 0 0 out_1[5]
port 14 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 out_1[6]
port 15 nsew signal tristate
flabel metal2 s 6458 31925 6514 32725 0 FreeSans 224 90 0 0 out_2[0]
port 16 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 out_2[1]
port 17 nsew signal tristate
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 out_2[2]
port 18 nsew signal tristate
flabel metal3 s 29781 2728 30581 2848 0 FreeSans 480 0 0 0 out_2[3]
port 19 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 out_2[4]
port 20 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 out_2[5]
port 21 nsew signal tristate
flabel metal2 s 2594 31925 2650 32725 0 FreeSans 224 90 0 0 out_2[6]
port 22 nsew signal tristate
flabel metal3 s 29781 6808 30581 6928 0 FreeSans 480 0 0 0 out_3[0]
port 23 nsew signal tristate
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 out_3[1]
port 24 nsew signal tristate
flabel metal3 s 29781 26528 30581 26648 0 FreeSans 480 0 0 0 out_3[2]
port 25 nsew signal tristate
flabel metal3 s 29781 30608 30581 30728 0 FreeSans 480 0 0 0 out_3[3]
port 26 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 out_3[4]
port 27 nsew signal tristate
flabel metal2 s 13542 31925 13598 32725 0 FreeSans 224 90 0 0 out_3[5]
port 28 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 out_3[6]
port 29 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 pb_0
port 30 nsew signal input
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 pb_1
port 31 nsew signal input
flabel metal3 s 29781 14288 30581 14408 0 FreeSans 480 0 0 0 time_done
port 32 nsew signal tristate
flabel metal4 s 4485 2128 4805 30512 0 FreeSans 1920 90 0 0 vccd1
port 33 nsew power bidirectional
flabel metal4 s 11568 2128 11888 30512 0 FreeSans 1920 90 0 0 vccd1
port 33 nsew power bidirectional
flabel metal4 s 18651 2128 18971 30512 0 FreeSans 1920 90 0 0 vccd1
port 33 nsew power bidirectional
flabel metal4 s 25734 2128 26054 30512 0 FreeSans 1920 90 0 0 vccd1
port 33 nsew power bidirectional
flabel metal4 s 8026 2128 8346 30512 0 FreeSans 1920 90 0 0 vssd1
port 34 nsew ground bidirectional
flabel metal4 s 15109 2128 15429 30512 0 FreeSans 1920 90 0 0 vssd1
port 34 nsew ground bidirectional
flabel metal4 s 22192 2128 22512 30512 0 FreeSans 1920 90 0 0 vssd1
port 34 nsew ground bidirectional
flabel metal4 s 29275 2128 29595 30512 0 FreeSans 1920 90 0 0 vssd1
port 34 nsew ground bidirectional
rlabel metal1 15272 29920 15272 29920 0 vccd1
rlabel via1 15349 30464 15349 30464 0 vssd1
rlabel metal1 5290 25840 5290 25840 0 CLKDIV.count\[0\]
rlabel metal1 11960 28186 11960 28186 0 CLKDIV.count\[10\]
rlabel metal1 11454 28050 11454 28050 0 CLKDIV.count\[11\]
rlabel metal1 11868 27438 11868 27438 0 CLKDIV.count\[12\]
rlabel metal1 13202 27506 13202 27506 0 CLKDIV.count\[13\]
rlabel metal1 14398 27846 14398 27846 0 CLKDIV.count\[14\]
rlabel metal2 15594 28016 15594 28016 0 CLKDIV.count\[15\]
rlabel metal2 18354 28458 18354 28458 0 CLKDIV.count\[16\]
rlabel metal1 17802 28118 17802 28118 0 CLKDIV.count\[17\]
rlabel metal1 17296 27982 17296 27982 0 CLKDIV.count\[18\]
rlabel metal1 19320 28186 19320 28186 0 CLKDIV.count\[19\]
rlabel metal2 4646 24990 4646 24990 0 CLKDIV.count\[1\]
rlabel metal1 21344 27302 21344 27302 0 CLKDIV.count\[20\]
rlabel metal1 24748 28662 24748 28662 0 CLKDIV.count\[21\]
rlabel metal1 22402 28458 22402 28458 0 CLKDIV.count\[22\]
rlabel metal2 21390 28458 21390 28458 0 CLKDIV.count\[23\]
rlabel metal2 5750 25194 5750 25194 0 CLKDIV.count\[2\]
rlabel metal1 6026 25908 6026 25908 0 CLKDIV.count\[3\]
rlabel metal1 5198 27438 5198 27438 0 CLKDIV.count\[4\]
rlabel metal2 6210 28288 6210 28288 0 CLKDIV.count\[5\]
rlabel metal1 5934 28730 5934 28730 0 CLKDIV.count\[6\]
rlabel metal1 6762 28016 6762 28016 0 CLKDIV.count\[7\]
rlabel metal1 9108 28594 9108 28594 0 CLKDIV.count\[8\]
rlabel metal1 9660 27982 9660 27982 0 CLKDIV.count\[9\]
rlabel metal1 17572 23698 17572 23698 0 CLKDIV.secpulse
rlabel metal1 16284 21862 16284 21862 0 CTR.minutes
rlabel metal1 20792 24786 20792 24786 0 CTR.time_out\[0\]
rlabel metal1 7774 6664 7774 6664 0 CTR.time_out\[10\]
rlabel metal1 15640 8534 15640 8534 0 CTR.time_out\[11\]
rlabel metal1 20286 24786 20286 24786 0 CTR.time_out\[1\]
rlabel metal2 19366 19516 19366 19516 0 CTR.time_out\[2\]
rlabel metal1 16882 25194 16882 25194 0 CTR.time_out\[3\]
rlabel metal1 11822 24072 11822 24072 0 CTR.time_out\[4\]
rlabel metal1 7038 22542 7038 22542 0 CTR.time_out\[5\]
rlabel metal1 7590 16150 7590 16150 0 CTR.time_out\[6\]
rlabel metal1 7636 11050 7636 11050 0 CTR.time_out\[7\]
rlabel metal1 14076 10574 14076 10574 0 CTR.time_out\[8\]
rlabel metal1 14076 7854 14076 7854 0 CTR.time_out\[9\]
rlabel metal1 20470 14586 20470 14586 0 FSM.next_state\[0\]
rlabel metal1 18354 12920 18354 12920 0 FSM.next_state\[1\]
rlabel metal1 20046 11322 20046 11322 0 FSM.next_state\[2\]
rlabel metal1 23138 10744 23138 10744 0 FSM.next_state\[3\]
rlabel metal1 22126 14960 22126 14960 0 FSM.state\[0\]
rlabel metal1 24288 11050 24288 11050 0 FSM.state\[1\]
rlabel metal1 23736 11730 23736 11730 0 FSM.state\[2\]
rlabel metal1 23644 11662 23644 11662 0 FSM.state\[3\]
rlabel metal1 10810 8942 10810 8942 0 MEM.addr\[0\]
rlabel metal1 10994 9010 10994 9010 0 MEM.addr\[1\]
rlabel metal2 12466 5236 12466 5236 0 MEM.addr\[2\]
rlabel metal2 16146 17442 16146 17442 0 MEM.mem1\[0\]
rlabel metal1 20010 8942 20010 8942 0 MEM.mem1\[10\]
rlabel metal1 15134 14518 15134 14518 0 MEM.mem1\[11\]
rlabel metal2 18446 21828 18446 21828 0 MEM.mem1\[1\]
rlabel metal1 18860 20978 18860 20978 0 MEM.mem1\[2\]
rlabel metal1 18906 17272 18906 17272 0 MEM.mem1\[3\]
rlabel metal1 15916 19278 15916 19278 0 MEM.mem1\[4\]
rlabel metal1 18860 18734 18860 18734 0 MEM.mem1\[5\]
rlabel metal1 15640 16014 15640 16014 0 MEM.mem1\[6\]
rlabel metal2 18078 11492 18078 11492 0 MEM.mem1\[7\]
rlabel metal2 18354 9724 18354 9724 0 MEM.mem1\[8\]
rlabel metal1 16652 13294 16652 13294 0 MEM.mem1\[9\]
rlabel viali 11546 17646 11546 17646 0 MEM.mem2\[0\]
rlabel metal1 6072 6222 6072 6222 0 MEM.mem2\[10\]
rlabel metal2 10994 15878 10994 15878 0 MEM.mem2\[11\]
rlabel metal1 10442 23290 10442 23290 0 MEM.mem2\[1\]
rlabel metal1 11500 22542 11500 22542 0 MEM.mem2\[2\]
rlabel metal1 5336 18054 5336 18054 0 MEM.mem2\[3\]
rlabel metal1 5474 21658 5474 21658 0 MEM.mem2\[4\]
rlabel metal1 7774 21318 7774 21318 0 MEM.mem2\[5\]
rlabel metal1 5888 15674 5888 15674 0 MEM.mem2\[6\]
rlabel metal1 6762 13294 6762 13294 0 MEM.mem2\[7\]
rlabel metal1 5658 6834 5658 6834 0 MEM.mem2\[8\]
rlabel metal1 10902 12750 10902 12750 0 MEM.mem2\[9\]
rlabel metal1 13662 18190 13662 18190 0 MEM.mem3\[0\]
rlabel metal1 8050 6290 8050 6290 0 MEM.mem3\[10\]
rlabel metal2 12650 15062 12650 15062 0 MEM.mem3\[11\]
rlabel metal1 11914 19278 11914 19278 0 MEM.mem3\[1\]
rlabel metal1 13984 20434 13984 20434 0 MEM.mem3\[2\]
rlabel metal1 7406 17680 7406 17680 0 MEM.mem3\[3\]
rlabel metal1 7682 20230 7682 20230 0 MEM.mem3\[4\]
rlabel metal1 8878 18938 8878 18938 0 MEM.mem3\[5\]
rlabel metal1 8234 14790 8234 14790 0 MEM.mem3\[6\]
rlabel metal1 7268 11730 7268 11730 0 MEM.mem3\[7\]
rlabel metal1 7314 6290 7314 6290 0 MEM.mem3\[8\]
rlabel metal1 13800 12818 13800 12818 0 MEM.mem3\[9\]
rlabel metal2 13938 18088 13938 18088 0 MEM.mem4\[0\]
rlabel metal1 4738 9010 4738 9010 0 MEM.mem4\[10\]
rlabel metal1 13662 15470 13662 15470 0 MEM.mem4\[11\]
rlabel metal1 12650 21590 12650 21590 0 MEM.mem4\[1\]
rlabel metal1 14490 20808 14490 20808 0 MEM.mem4\[2\]
rlabel metal1 5796 15130 5796 15130 0 MEM.mem4\[3\]
rlabel metal1 3910 19754 3910 19754 0 MEM.mem4\[4\]
rlabel metal1 9292 19278 9292 19278 0 MEM.mem4\[5\]
rlabel metal1 8556 15674 8556 15674 0 MEM.mem4\[6\]
rlabel metal1 4554 11084 4554 11084 0 MEM.mem4\[7\]
rlabel metal1 3910 9690 3910 9690 0 MEM.mem4\[8\]
rlabel metal1 14030 12206 14030 12206 0 MEM.mem4\[9\]
rlabel metal2 11362 18020 11362 18020 0 MEM.mem5\[0\]
rlabel metal1 4186 8330 4186 8330 0 MEM.mem5\[10\]
rlabel metal1 11040 15674 11040 15674 0 MEM.mem5\[11\]
rlabel metal1 10902 23494 10902 23494 0 MEM.mem5\[1\]
rlabel metal2 10810 21148 10810 21148 0 MEM.mem5\[2\]
rlabel metal1 4692 18734 4692 18734 0 MEM.mem5\[3\]
rlabel metal1 5106 22542 5106 22542 0 MEM.mem5\[4\]
rlabel metal1 7728 22202 7728 22202 0 MEM.mem5\[5\]
rlabel metal1 4462 15980 4462 15980 0 MEM.mem5\[6\]
rlabel metal1 4370 11730 4370 11730 0 MEM.mem5\[7\]
rlabel metal1 4232 7854 4232 7854 0 MEM.mem5\[8\]
rlabel metal2 10810 13566 10810 13566 0 MEM.mem5\[9\]
rlabel metal1 15548 17034 15548 17034 0 MEM.next_mem1\[0\]
rlabel metal1 18860 8398 18860 8398 0 MEM.next_mem1\[10\]
rlabel metal2 15502 14348 15502 14348 0 MEM.next_mem1\[11\]
rlabel metal1 16744 21114 16744 21114 0 MEM.next_mem1\[1\]
rlabel metal1 17526 20230 17526 20230 0 MEM.next_mem1\[2\]
rlabel metal1 18216 17306 18216 17306 0 MEM.next_mem1\[3\]
rlabel metal1 14996 18802 14996 18802 0 MEM.next_mem1\[4\]
rlabel metal1 17342 18360 17342 18360 0 MEM.next_mem1\[5\]
rlabel metal1 15502 15538 15502 15538 0 MEM.next_mem1\[6\]
rlabel metal1 16422 11050 16422 11050 0 MEM.next_mem1\[7\]
rlabel metal1 17066 9690 17066 9690 0 MEM.next_mem1\[8\]
rlabel metal1 15042 12920 15042 12920 0 MEM.next_mem1\[9\]
rlabel metal2 9890 17578 9890 17578 0 MEM.next_mem2\[0\]
rlabel metal1 5421 5882 5421 5882 0 MEM.next_mem2\[10\]
rlabel metal1 9522 15096 9522 15096 0 MEM.next_mem2\[11\]
rlabel metal2 9246 22746 9246 22746 0 MEM.next_mem2\[1\]
rlabel metal1 9660 21862 9660 21862 0 MEM.next_mem2\[2\]
rlabel metal1 5152 17306 5152 17306 0 MEM.next_mem2\[3\]
rlabel metal1 5382 23086 5382 23086 0 MEM.next_mem2\[4\]
rlabel metal1 7728 21454 7728 21454 0 MEM.next_mem2\[5\]
rlabel metal1 4554 15368 4554 15368 0 MEM.next_mem2\[6\]
rlabel metal1 5842 12274 5842 12274 0 MEM.next_mem2\[7\]
rlabel metal1 4186 6392 4186 6392 0 MEM.next_mem2\[8\]
rlabel metal1 10948 13430 10948 13430 0 MEM.next_mem2\[9\]
rlabel metal1 12466 17272 12466 17272 0 MEM.next_mem3\[0\]
rlabel metal1 6670 5304 6670 5304 0 MEM.next_mem3\[10\]
rlabel metal1 11822 14450 11822 14450 0 MEM.next_mem3\[11\]
rlabel metal1 10810 18802 10810 18802 0 MEM.next_mem3\[1\]
rlabel metal2 12098 20196 12098 20196 0 MEM.next_mem3\[2\]
rlabel metal1 5704 17578 5704 17578 0 MEM.next_mem3\[3\]
rlabel metal1 6808 20026 6808 20026 0 MEM.next_mem3\[4\]
rlabel metal1 7590 18802 7590 18802 0 MEM.next_mem3\[5\]
rlabel metal1 7268 14586 7268 14586 0 MEM.next_mem3\[6\]
rlabel metal1 6801 11322 6801 11322 0 MEM.next_mem3\[7\]
rlabel metal1 6762 5746 6762 5746 0 MEM.next_mem3\[8\]
rlabel metal2 12834 12517 12834 12517 0 MEM.next_mem3\[9\]
rlabel metal2 14674 17136 14674 17136 0 MEM.next_mem4\[0\]
rlabel metal2 5658 9248 5658 9248 0 MEM.next_mem4\[10\]
rlabel metal2 12466 15198 12466 15198 0 MEM.next_mem4\[11\]
rlabel metal1 13340 19482 13340 19482 0 MEM.next_mem4\[1\]
rlabel metal1 14628 20570 14628 20570 0 MEM.next_mem4\[2\]
rlabel metal1 4968 14926 4968 14926 0 MEM.next_mem4\[3\]
rlabel metal1 3910 19958 3910 19958 0 MEM.next_mem4\[4\]
rlabel metal1 8372 19414 8372 19414 0 MEM.next_mem4\[5\]
rlabel metal1 7268 15538 7268 15538 0 MEM.next_mem4\[6\]
rlabel metal1 4692 10778 4692 10778 0 MEM.next_mem4\[7\]
rlabel metal2 4186 9962 4186 9962 0 MEM.next_mem4\[8\]
rlabel metal1 15364 12342 15364 12342 0 MEM.next_mem4\[9\]
rlabel metal1 10028 17578 10028 17578 0 MEM.next_mem5\[0\]
rlabel metal1 4554 8364 4554 8364 0 MEM.next_mem5\[10\]
rlabel metal1 9745 15674 9745 15674 0 MEM.next_mem5\[11\]
rlabel metal1 10902 23664 10902 23664 0 MEM.next_mem5\[1\]
rlabel metal1 10626 20298 10626 20298 0 MEM.next_mem5\[2\]
rlabel metal2 4554 17442 4554 17442 0 MEM.next_mem5\[3\]
rlabel metal1 3900 21114 3900 21114 0 MEM.next_mem5\[4\]
rlabel metal2 7314 22304 7314 22304 0 MEM.next_mem5\[5\]
rlabel metal2 3358 16252 3358 16252 0 MEM.next_mem5\[6\]
rlabel metal2 4370 11492 4370 11492 0 MEM.next_mem5\[7\]
rlabel metal1 4002 7990 4002 7990 0 MEM.next_mem5\[8\]
rlabel metal1 9522 12920 9522 12920 0 MEM.next_mem5\[9\]
rlabel metal1 9246 8568 9246 8568 0 MEM.raddr\[0\]
rlabel metal1 10557 11730 10557 11730 0 MEM.raddr\[1\]
rlabel metal1 6394 9622 6394 9622 0 MEM.raddr\[2\]
rlabel metal1 21298 17850 21298 17850 0 TIM.cnt\[0\]
rlabel metal1 18170 7820 18170 7820 0 TIM.cnt\[10\]
rlabel metal1 22379 9554 22379 9554 0 TIM.cnt\[11\]
rlabel metal1 22678 17646 22678 17646 0 TIM.cnt\[1\]
rlabel metal1 19642 19720 19642 19720 0 TIM.cnt\[2\]
rlabel metal2 20286 17663 20286 17663 0 TIM.cnt\[3\]
rlabel metal2 19734 19584 19734 19584 0 TIM.cnt\[4\]
rlabel metal2 23322 17680 23322 17680 0 TIM.cnt\[5\]
rlabel metal1 18262 9928 18262 9928 0 TIM.cnt\[6\]
rlabel metal2 23322 8160 23322 8160 0 TIM.cnt\[7\]
rlabel metal2 17526 8806 17526 8806 0 TIM.cnt\[8\]
rlabel metal2 17434 7905 17434 7905 0 TIM.cnt\[9\]
rlabel metal1 7537 25466 7537 25466 0 _0000_
rlabel metal1 10948 28594 10948 28594 0 _0001_
rlabel metal1 11224 29002 11224 29002 0 _0002_
rlabel metal1 11171 26554 11171 26554 0 _0003_
rlabel metal1 12926 27506 12926 27506 0 _0004_
rlabel metal1 14352 27982 14352 27982 0 _0005_
rlabel metal1 14352 28730 14352 28730 0 _0006_
rlabel metal1 16974 29240 16974 29240 0 _0007_
rlabel metal1 17112 28594 17112 28594 0 _0008_
rlabel metal1 16790 27336 16790 27336 0 _0009_
rlabel metal1 19320 27982 19320 27982 0 _0010_
rlabel metal1 3772 24378 3772 24378 0 _0011_
rlabel metal2 22586 27744 22586 27744 0 _0012_
rlabel metal1 22954 28594 22954 28594 0 _0013_
rlabel metal2 23230 28560 23230 28560 0 _0014_
rlabel metal1 20332 29206 20332 29206 0 _0015_
rlabel metal1 5934 24072 5934 24072 0 _0016_
rlabel metal1 5053 25466 5053 25466 0 _0017_
rlabel metal1 3496 28186 3496 28186 0 _0018_
rlabel metal1 3818 28118 3818 28118 0 _0019_
rlabel metal1 4784 28458 4784 28458 0 _0020_
rlabel metal1 7038 29036 7038 29036 0 _0021_
rlabel metal1 7498 28118 7498 28118 0 _0022_
rlabel metal1 8234 27064 8234 27064 0 _0023_
rlabel metal1 8418 25942 8418 25942 0 _0024_
rlabel metal1 20654 7922 20654 7922 0 _0025_
rlabel metal1 21429 6970 21429 6970 0 _0026_
rlabel metal1 23591 6970 23591 6970 0 _0027_
rlabel metal1 25438 7446 25438 7446 0 _0028_
rlabel metal1 26542 8840 26542 8840 0 _0029_
rlabel metal1 25346 10778 25346 10778 0 _0030_
rlabel metal1 14805 22202 14805 22202 0 _0031_
rlabel metal1 2070 13498 2070 13498 0 _0032_
rlabel metal1 2392 12410 2392 12410 0 _0033_
rlabel metal1 13708 9622 13708 9622 0 _0034_
rlabel metal1 13432 7446 13432 7446 0 _0035_
rlabel metal1 13754 6392 13754 6392 0 _0036_
rlabel via1 13665 8806 13665 8806 0 _0037_
rlabel metal1 23276 17850 23276 17850 0 _0038_
rlabel metal1 24646 14586 24646 14586 0 _0039_
rlabel metal2 27094 14620 27094 14620 0 _0040_
rlabel metal1 27232 17850 27232 17850 0 _0041_
rlabel metal1 23782 17272 23782 17272 0 _0042_
rlabel metal1 24564 13838 24564 13838 0 _0043_
rlabel metal1 9246 9010 9246 9010 0 _0044_
rlabel metal1 9752 10778 9752 10778 0 _0045_
rlabel metal2 6578 9180 6578 9180 0 _0046_
rlabel metal1 20608 17306 20608 17306 0 _0047_
rlabel metal2 9338 5100 9338 5100 0 _0048_
rlabel metal1 9338 5134 9338 5134 0 _0049_
rlabel metal1 11868 5202 11868 5202 0 _0050_
rlabel metal1 17986 24650 17986 24650 0 _0051_
rlabel metal1 18584 24854 18584 24854 0 _0052_
rlabel metal1 16698 24072 16698 24072 0 _0053_
rlabel metal2 14950 25058 14950 25058 0 _0054_
rlabel metal1 11914 23800 11914 23800 0 _0055_
rlabel metal1 11868 24854 11868 24854 0 _0056_
rlabel metal1 6026 25806 6026 25806 0 _0057_
rlabel metal2 5658 25228 5658 25228 0 _0058_
rlabel metal1 7084 26010 7084 26010 0 _0059_
rlabel metal1 14444 27574 14444 27574 0 _0060_
rlabel metal1 11500 27846 11500 27846 0 _0061_
rlabel via2 13662 28611 13662 28611 0 _0062_
rlabel metal2 17986 28169 17986 28169 0 _0063_
rlabel metal1 8096 27438 8096 27438 0 _0064_
rlabel metal1 12282 28424 12282 28424 0 _0065_
rlabel metal2 19366 14212 19366 14212 0 _0066_
rlabel metal1 18998 13260 18998 13260 0 _0067_
rlabel metal1 18952 10778 18952 10778 0 _0068_
rlabel metal1 15548 13430 15548 13430 0 _0069_
rlabel metal2 10074 20366 10074 20366 0 _0070_
rlabel metal1 15456 19822 15456 19822 0 _0071_
rlabel metal1 6808 9622 6808 9622 0 _0072_
rlabel metal1 8142 13328 8142 13328 0 _0073_
rlabel metal1 7774 12410 7774 12410 0 _0074_
rlabel metal1 8464 12750 8464 12750 0 _0075_
rlabel metal1 5796 18258 5796 18258 0 _0076_
rlabel metal2 11086 14076 11086 14076 0 _0077_
rlabel metal1 14490 13294 14490 13294 0 _0078_
rlabel metal2 7314 18700 7314 18700 0 _0079_
rlabel metal1 14214 13940 14214 13940 0 _0080_
rlabel metal1 15548 13702 15548 13702 0 _0081_
rlabel metal1 22011 13294 22011 13294 0 _0082_
rlabel metal1 22908 10778 22908 10778 0 _0083_
rlabel metal1 22954 13260 22954 13260 0 _0084_
rlabel metal1 19826 19346 19826 19346 0 _0085_
rlabel metal2 15824 14382 15824 14382 0 _0086_
rlabel metal1 16330 11526 16330 11526 0 _0087_
rlabel metal1 16928 7514 16928 7514 0 _0088_
rlabel metal1 16146 13192 16146 13192 0 _0089_
rlabel metal2 14674 13158 14674 13158 0 _0090_
rlabel metal1 15594 13260 15594 13260 0 _0091_
rlabel metal1 16882 13430 16882 13430 0 _0092_
rlabel metal1 17296 6766 17296 6766 0 _0093_
rlabel metal1 5382 8466 5382 8466 0 _0094_
rlabel metal1 5474 7514 5474 7514 0 _0095_
rlabel metal1 5382 8398 5382 8398 0 _0096_
rlabel metal1 5336 8534 5336 8534 0 _0097_
rlabel metal2 5474 8840 5474 8840 0 _0098_
rlabel via1 17968 7854 17968 7854 0 _0099_
rlabel metal1 17158 7412 17158 7412 0 _0100_
rlabel metal2 17434 6970 17434 6970 0 _0101_
rlabel metal1 17342 4998 17342 4998 0 _0102_
rlabel metal1 18722 5168 18722 5168 0 _0103_
rlabel metal1 6946 7854 6946 7854 0 _0104_
rlabel metal1 5842 8058 5842 8058 0 _0105_
rlabel metal1 6762 7922 6762 7922 0 _0106_
rlabel metal1 6164 7786 6164 7786 0 _0107_
rlabel metal2 12834 7718 12834 7718 0 _0108_
rlabel metal1 17324 8466 17324 8466 0 _0109_
rlabel metal1 17112 8466 17112 8466 0 _0110_
rlabel metal2 18538 4352 18538 4352 0 _0111_
rlabel metal1 18216 5542 18216 5542 0 _0112_
rlabel metal1 17434 6358 17434 6358 0 _0113_
rlabel metal1 6946 10642 6946 10642 0 _0114_
rlabel metal1 6578 10506 6578 10506 0 _0115_
rlabel metal1 6348 10574 6348 10574 0 _0116_
rlabel metal1 5980 10710 5980 10710 0 _0117_
rlabel metal1 9614 10744 9614 10744 0 _0118_
rlabel metal1 17048 10642 17048 10642 0 _0119_
rlabel metal1 16698 10642 16698 10642 0 _0120_
rlabel metal1 18032 6766 18032 6766 0 _0121_
rlabel metal2 16974 5338 16974 5338 0 _0122_
rlabel metal1 17526 4726 17526 4726 0 _0123_
rlabel metal1 16376 4658 16376 4658 0 _0124_
rlabel metal1 18630 4556 18630 4556 0 _0125_
rlabel metal1 19366 4658 19366 4658 0 _0126_
rlabel metal1 18124 3026 18124 3026 0 _0127_
rlabel metal1 19780 4590 19780 4590 0 _0128_
rlabel metal1 17480 6426 17480 6426 0 _0129_
rlabel metal1 20516 4590 20516 4590 0 _0130_
rlabel metal1 19642 5134 19642 5134 0 _0131_
rlabel metal1 20194 5202 20194 5202 0 _0132_
rlabel metal2 20194 3740 20194 3740 0 _0133_
rlabel metal1 19918 4556 19918 4556 0 _0134_
rlabel metal2 28106 4998 28106 4998 0 _0135_
rlabel metal1 5060 24786 5060 24786 0 _0136_
rlabel metal1 4278 24242 4278 24242 0 _0137_
rlabel metal1 6486 25772 6486 25772 0 _0138_
rlabel metal1 5750 26384 5750 26384 0 _0139_
rlabel metal2 5198 24854 5198 24854 0 _0140_
rlabel metal2 5842 26078 5842 26078 0 _0141_
rlabel metal2 4278 28050 4278 28050 0 _0142_
rlabel metal1 4416 27438 4416 27438 0 _0143_
rlabel metal1 4646 27608 4646 27608 0 _0144_
rlabel metal1 6210 27948 6210 27948 0 _0145_
rlabel metal2 5842 28696 5842 28696 0 _0146_
rlabel metal2 6026 28866 6026 28866 0 _0147_
rlabel metal1 7590 28730 7590 28730 0 _0148_
rlabel metal2 7314 28288 7314 28288 0 _0149_
rlabel via1 6854 29155 6854 29155 0 _0150_
rlabel metal1 8004 28390 8004 28390 0 _0151_
rlabel metal1 8510 28594 8510 28594 0 _0152_
rlabel metal1 9936 28186 9936 28186 0 _0153_
rlabel metal1 9154 27404 9154 27404 0 _0154_
rlabel metal1 11408 28730 11408 28730 0 _0155_
rlabel metal2 11270 28628 11270 28628 0 _0156_
rlabel metal1 11362 29206 11362 29206 0 _0157_
rlabel metal1 12052 27438 12052 27438 0 _0158_
rlabel viali 11733 26894 11733 26894 0 _0159_
rlabel metal2 11914 27098 11914 27098 0 _0160_
rlabel metal1 15318 28458 15318 28458 0 _0161_
rlabel metal1 14398 26860 14398 26860 0 _0162_
rlabel metal1 14536 28662 14536 28662 0 _0163_
rlabel metal1 15134 28492 15134 28492 0 _0164_
rlabel metal2 16238 29410 16238 29410 0 _0165_
rlabel metal2 16698 28968 16698 28968 0 _0166_
rlabel metal2 16514 29410 16514 29410 0 _0167_
rlabel metal1 17204 27846 17204 27846 0 _0168_
rlabel metal1 17802 26826 17802 26826 0 _0169_
rlabel metal1 17020 27098 17020 27098 0 _0170_
rlabel metal1 19366 27438 19366 27438 0 _0171_
rlabel metal2 22678 27744 22678 27744 0 _0172_
rlabel metal1 21068 27098 21068 27098 0 _0173_
rlabel metal2 22126 27982 22126 27982 0 _0174_
rlabel metal1 22816 27506 22816 27506 0 _0175_
rlabel metal1 20378 28696 20378 28696 0 _0176_
rlabel metal1 20532 28458 20532 28458 0 _0177_
rlabel metal1 20700 28730 20700 28730 0 _0178_
rlabel metal1 6992 19822 6992 19822 0 _0179_
rlabel metal1 7682 19720 7682 19720 0 _0180_
rlabel metal1 16514 20026 16514 20026 0 _0181_
rlabel metal2 17250 19958 17250 19958 0 _0182_
rlabel metal1 21482 21420 21482 21420 0 _0183_
rlabel metal1 6486 13498 6486 13498 0 _0184_
rlabel metal2 6394 15776 6394 15776 0 _0185_
rlabel metal2 7682 17850 7682 17850 0 _0186_
rlabel metal2 19458 17935 19458 17935 0 _0187_
rlabel metal2 19274 17748 19274 17748 0 _0188_
rlabel metal2 12650 19006 12650 19006 0 _0189_
rlabel metal2 19826 18054 19826 18054 0 _0190_
rlabel metal1 20700 18122 20700 18122 0 _0191_
rlabel metal1 13754 20842 13754 20842 0 _0192_
rlabel metal1 18492 21522 18492 21522 0 _0193_
rlabel metal1 19550 21012 19550 21012 0 _0194_
rlabel metal1 20056 20978 20056 20978 0 _0195_
rlabel metal1 23874 20366 23874 20366 0 _0196_
rlabel metal1 11592 21862 11592 21862 0 _0197_
rlabel metal1 19044 20434 19044 20434 0 _0198_
rlabel metal1 18722 20502 18722 20502 0 _0199_
rlabel metal2 8694 22406 8694 22406 0 _0200_
rlabel metal2 20562 19924 20562 19924 0 _0201_
rlabel metal2 19274 20570 19274 20570 0 _0202_
rlabel metal2 22126 21029 22126 21029 0 _0203_
rlabel metal1 8786 18734 8786 18734 0 _0204_
rlabel metal2 17986 19346 17986 19346 0 _0205_
rlabel metal1 20102 18938 20102 18938 0 _0206_
rlabel metal1 19642 18938 19642 18938 0 _0207_
rlabel metal2 21298 20026 21298 20026 0 _0208_
rlabel metal1 22954 21998 22954 21998 0 _0209_
rlabel metal1 21620 21658 21620 21658 0 _0210_
rlabel metal2 20838 21828 20838 21828 0 _0211_
rlabel metal1 21022 21454 21022 21454 0 _0212_
rlabel metal1 21160 21386 21160 21386 0 _0213_
rlabel metal1 25438 22032 25438 22032 0 _0214_
rlabel metal1 24288 4182 24288 4182 0 _0215_
rlabel metal1 23000 22678 23000 22678 0 _0216_
rlabel metal1 24564 21998 24564 21998 0 _0217_
rlabel metal1 23874 21556 23874 21556 0 _0218_
rlabel metal1 25208 21862 25208 21862 0 _0219_
rlabel metal1 21574 22644 21574 22644 0 _0220_
rlabel metal1 24564 4114 24564 4114 0 _0221_
rlabel metal1 25208 3502 25208 3502 0 _0222_
rlabel metal1 24748 22066 24748 22066 0 _0223_
rlabel metal1 25622 21998 25622 21998 0 _0224_
rlabel metal1 25438 20978 25438 20978 0 _0225_
rlabel metal2 2438 4063 2438 4063 0 _0226_
rlabel metal1 2599 3502 2599 3502 0 _0227_
rlabel metal2 25254 26452 25254 26452 0 _0228_
rlabel via1 20470 18258 20470 18258 0 _0229_
rlabel metal1 11546 9622 11546 9622 0 _0230_
rlabel metal2 19780 13260 19780 13260 0 _0231_
rlabel metal1 12489 9554 12489 9554 0 _0232_
rlabel metal1 17112 12818 17112 12818 0 _0233_
rlabel metal1 22034 11322 22034 11322 0 _0234_
rlabel metal1 24150 11118 24150 11118 0 _0235_
rlabel metal1 16606 18700 16606 18700 0 _0236_
rlabel metal1 15134 13872 15134 13872 0 _0237_
rlabel metal1 19918 15436 19918 15436 0 _0238_
rlabel metal1 10350 7412 10350 7412 0 _0239_
rlabel metal1 9062 22576 9062 22576 0 _0240_
rlabel metal1 11132 6358 11132 6358 0 _0241_
rlabel metal1 12420 9894 12420 9894 0 _0242_
rlabel metal1 10580 6426 10580 6426 0 _0243_
rlabel metal2 10074 16371 10074 16371 0 _0244_
rlabel metal1 11684 6290 11684 6290 0 _0245_
rlabel metal1 7682 14382 7682 14382 0 _0246_
rlabel metal1 7314 14348 7314 14348 0 _0247_
rlabel metal1 11592 8942 11592 8942 0 _0248_
rlabel metal2 13202 19584 13202 19584 0 _0249_
rlabel metal1 13938 19346 13938 19346 0 _0250_
rlabel metal2 11086 6307 11086 6307 0 _0251_
rlabel metal2 11362 7174 11362 7174 0 _0252_
rlabel metal1 7636 22610 7636 22610 0 _0253_
rlabel metal1 6854 22474 6854 22474 0 _0254_
rlabel metal2 12650 18054 12650 18054 0 _0255_
rlabel metal1 17342 17238 17342 17238 0 _0256_
rlabel metal1 17526 17102 17526 17102 0 _0257_
rlabel metal1 23184 18394 23184 18394 0 _0258_
rlabel metal1 27370 20876 27370 20876 0 _0259_
rlabel metal1 25944 20774 25944 20774 0 _0260_
rlabel metal1 28290 20978 28290 20978 0 _0261_
rlabel metal1 23690 20468 23690 20468 0 _0262_
rlabel metal1 24104 20570 24104 20570 0 _0263_
rlabel metal1 20838 22746 20838 22746 0 _0264_
rlabel metal1 20654 22066 20654 22066 0 _0265_
rlabel metal1 21160 21930 21160 21930 0 _0266_
rlabel metal1 21482 22678 21482 22678 0 _0267_
rlabel metal2 21114 22202 21114 22202 0 _0268_
rlabel metal2 21666 22338 21666 22338 0 _0269_
rlabel metal1 23966 22644 23966 22644 0 _0270_
rlabel metal1 24656 22474 24656 22474 0 _0271_
rlabel metal1 24380 21522 24380 21522 0 _0272_
rlabel metal1 26220 20910 26220 20910 0 _0273_
rlabel metal1 27554 19686 27554 19686 0 _0274_
rlabel metal2 27554 20026 27554 20026 0 _0275_
rlabel metal1 22264 21998 22264 21998 0 _0276_
rlabel via1 22954 21947 22954 21947 0 _0277_
rlabel metal1 22678 22032 22678 22032 0 _0278_
rlabel metal1 22540 21522 22540 21522 0 _0279_
rlabel metal1 21804 20230 21804 20230 0 _0280_
rlabel metal1 21720 20570 21720 20570 0 _0281_
rlabel metal1 22402 20570 22402 20570 0 _0282_
rlabel metal1 21850 21488 21850 21488 0 _0283_
rlabel metal2 21850 21471 21850 21471 0 _0284_
rlabel metal2 27278 20570 27278 20570 0 _0285_
rlabel metal1 27048 21114 27048 21114 0 _0286_
rlabel metal1 27876 20026 27876 20026 0 _0287_
rlabel metal1 28290 19822 28290 19822 0 _0288_
rlabel viali 28567 20456 28567 20456 0 _0289_
rlabel metal1 16790 3536 16790 3536 0 _0290_
rlabel metal1 18078 5678 18078 5678 0 _0291_
rlabel metal1 18400 3162 18400 3162 0 _0292_
rlabel metal1 18170 3366 18170 3366 0 _0293_
rlabel metal1 17388 3026 17388 3026 0 _0294_
rlabel metal1 17204 2958 17204 2958 0 _0295_
rlabel metal1 16882 3468 16882 3468 0 _0296_
rlabel metal1 16008 3502 16008 3502 0 _0297_
rlabel metal2 19550 3876 19550 3876 0 _0298_
rlabel metal1 13079 4114 13079 4114 0 _0299_
rlabel metal2 16330 4318 16330 4318 0 _0300_
rlabel metal1 17079 5338 17079 5338 0 _0301_
rlabel metal1 17388 4658 17388 4658 0 _0302_
rlabel metal1 16790 7344 16790 7344 0 _0303_
rlabel metal1 17894 6800 17894 6800 0 _0304_
rlabel metal1 17618 6290 17618 6290 0 _0305_
rlabel metal2 17618 5440 17618 5440 0 _0306_
rlabel metal1 16744 4046 16744 4046 0 _0307_
rlabel metal1 13708 2414 13708 2414 0 _0308_
rlabel metal2 8418 15470 8418 15470 0 _0309_
rlabel metal1 14030 15028 14030 15028 0 _0310_
rlabel metal2 15548 16116 15548 16116 0 _0311_
rlabel metal1 15824 9894 15824 9894 0 _0312_
rlabel metal1 13524 2414 13524 2414 0 _0313_
rlabel metal1 13386 2618 13386 2618 0 _0314_
rlabel metal2 14030 3774 14030 3774 0 _0315_
rlabel metal2 14582 3400 14582 3400 0 _0316_
rlabel metal1 15134 3366 15134 3366 0 _0317_
rlabel metal2 2438 5575 2438 5575 0 _0318_
rlabel metal1 14076 3366 14076 3366 0 _0319_
rlabel metal1 12926 3706 12926 3706 0 _0320_
rlabel metal1 10304 24582 10304 24582 0 _0321_
rlabel metal1 20516 14382 20516 14382 0 _0322_
rlabel metal1 19688 15470 19688 15470 0 _0323_
rlabel metal1 19504 14994 19504 14994 0 _0324_
rlabel metal1 19458 14790 19458 14790 0 _0325_
rlabel metal1 21390 12716 21390 12716 0 _0326_
rlabel metal1 24656 16558 24656 16558 0 _0327_
rlabel metal1 20194 15538 20194 15538 0 _0328_
rlabel viali 21758 14382 21758 14382 0 _0329_
rlabel metal1 18492 14586 18492 14586 0 _0330_
rlabel metal1 21436 12954 21436 12954 0 _0331_
rlabel metal1 20378 14348 20378 14348 0 _0332_
rlabel metal1 20286 14042 20286 14042 0 _0333_
rlabel metal1 20792 14382 20792 14382 0 _0334_
rlabel metal1 16284 14994 16284 14994 0 _0335_
rlabel metal1 17572 14382 17572 14382 0 _0336_
rlabel metal1 18676 13498 18676 13498 0 _0337_
rlabel metal1 18906 13940 18906 13940 0 _0338_
rlabel metal1 19044 13906 19044 13906 0 _0339_
rlabel metal1 17940 11186 17940 11186 0 _0340_
rlabel metal1 19826 13974 19826 13974 0 _0341_
rlabel metal1 19458 14314 19458 14314 0 _0342_
rlabel metal2 19274 13770 19274 13770 0 _0343_
rlabel metal1 19872 12206 19872 12206 0 _0344_
rlabel metal2 21850 12988 21850 12988 0 _0345_
rlabel metal1 23736 12274 23736 12274 0 _0346_
rlabel metal2 22126 9418 22126 9418 0 _0347_
rlabel metal1 26266 16558 26266 16558 0 _0348_
rlabel metal2 23782 16014 23782 16014 0 _0349_
rlabel metal1 26496 16422 26496 16422 0 _0350_
rlabel metal1 27784 17510 27784 17510 0 _0351_
rlabel metal1 23276 16558 23276 16558 0 _0352_
rlabel metal1 23230 16456 23230 16456 0 _0353_
rlabel metal1 23322 14926 23322 14926 0 _0354_
rlabel metal1 22954 9146 22954 9146 0 _0355_
rlabel metal1 23414 14042 23414 14042 0 _0356_
rlabel metal1 23276 14586 23276 14586 0 _0357_
rlabel metal2 24058 16558 24058 16558 0 _0358_
rlabel metal2 23598 16320 23598 16320 0 _0359_
rlabel metal1 23276 17102 23276 17102 0 _0360_
rlabel metal2 24012 11628 24012 11628 0 _0361_
rlabel metal1 24380 6766 24380 6766 0 _0362_
rlabel metal1 21436 8466 21436 8466 0 _0363_
rlabel metal2 24058 7684 24058 7684 0 _0364_
rlabel metal2 22954 7888 22954 7888 0 _0365_
rlabel metal1 23092 8058 23092 8058 0 _0366_
rlabel metal1 22632 7514 22632 7514 0 _0367_
rlabel via1 22586 7837 22586 7837 0 _0368_
rlabel metal1 23828 8330 23828 8330 0 _0369_
rlabel metal2 23782 8126 23782 8126 0 _0370_
rlabel metal1 24702 7446 24702 7446 0 _0371_
rlabel metal2 24702 8058 24702 8058 0 _0372_
rlabel metal1 23874 7344 23874 7344 0 _0373_
rlabel metal2 27554 8160 27554 8160 0 _0374_
rlabel metal1 27324 7378 27324 7378 0 _0375_
rlabel metal1 25944 8330 25944 8330 0 _0376_
rlabel metal1 26542 7514 26542 7514 0 _0377_
rlabel metal1 25852 7854 25852 7854 0 _0378_
rlabel metal1 27462 8534 27462 8534 0 _0379_
rlabel metal2 27278 8738 27278 8738 0 _0380_
rlabel metal1 26496 9350 26496 9350 0 _0381_
rlabel metal2 25806 8704 25806 8704 0 _0382_
rlabel metal1 25668 8942 25668 8942 0 _0383_
rlabel metal1 26312 10642 26312 10642 0 _0384_
rlabel metal2 25622 10404 25622 10404 0 _0385_
rlabel metal1 25944 10642 25944 10642 0 _0386_
rlabel metal1 14628 23290 14628 23290 0 _0387_
rlabel metal1 15686 23800 15686 23800 0 _0388_
rlabel metal1 18216 24854 18216 24854 0 _0389_
rlabel metal2 15962 23018 15962 23018 0 _0390_
rlabel metal2 16744 14246 16744 14246 0 _0391_
rlabel metal1 3312 13158 3312 13158 0 _0392_
rlabel metal1 2530 13294 2530 13294 0 _0393_
rlabel metal1 2990 12274 2990 12274 0 _0394_
rlabel metal1 2898 12138 2898 12138 0 _0395_
rlabel metal1 14674 10778 14674 10778 0 _0396_
rlabel metal2 13570 10336 13570 10336 0 _0397_
rlabel metal1 14352 7854 14352 7854 0 _0398_
rlabel metal2 13110 9520 13110 9520 0 _0399_
rlabel metal1 14122 10030 14122 10030 0 _0400_
rlabel metal2 14490 7344 14490 7344 0 _0401_
rlabel metal1 13064 7378 13064 7378 0 _0402_
rlabel metal2 13938 7310 13938 7310 0 _0403_
rlabel metal1 14306 6732 14306 6732 0 _0404_
rlabel metal1 13340 8602 13340 8602 0 _0405_
rlabel metal1 23690 17544 23690 17544 0 _0406_
rlabel via1 22678 17714 22678 17714 0 _0407_
rlabel metal2 23138 17238 23138 17238 0 _0408_
rlabel metal1 23000 16762 23000 16762 0 _0409_
rlabel metal1 23506 17306 23506 17306 0 _0410_
rlabel metal2 23782 17238 23782 17238 0 _0411_
rlabel viali 26634 16559 26634 16559 0 _0412_
rlabel metal1 26818 15538 26818 15538 0 _0413_
rlabel metal1 26220 15674 26220 15674 0 _0414_
rlabel metal1 27324 16762 27324 16762 0 _0415_
rlabel metal1 26542 15504 26542 15504 0 _0416_
rlabel metal2 24702 14943 24702 14943 0 _0417_
rlabel metal1 27462 15538 27462 15538 0 _0418_
rlabel metal1 27232 15062 27232 15062 0 _0419_
rlabel metal1 27830 16558 27830 16558 0 _0420_
rlabel metal2 27278 15946 27278 15946 0 _0421_
rlabel metal2 27232 14994 27232 14994 0 _0422_
rlabel metal1 27002 17034 27002 17034 0 _0423_
rlabel metal1 27278 17000 27278 17000 0 _0424_
rlabel metal1 27370 17068 27370 17068 0 _0425_
rlabel viali 28104 16552 28104 16552 0 _0426_
rlabel metal1 27738 17170 27738 17170 0 _0427_
rlabel metal1 26818 17306 26818 17306 0 _0428_
rlabel metal1 25668 17306 25668 17306 0 _0429_
rlabel metal2 25346 17204 25346 17204 0 _0430_
rlabel metal1 9476 10098 9476 10098 0 _0431_
rlabel metal1 9200 9554 9200 9554 0 _0432_
rlabel metal1 10810 10098 10810 10098 0 _0433_
rlabel metal1 10396 10234 10396 10234 0 _0434_
rlabel metal2 10626 10098 10626 10098 0 _0435_
rlabel metal1 10166 9656 10166 9656 0 _0436_
rlabel metal1 11040 9418 11040 9418 0 _0437_
rlabel metal1 10557 9622 10557 9622 0 _0438_
rlabel metal1 8970 9452 8970 9452 0 _0439_
rlabel metal1 22356 16762 22356 16762 0 _0440_
rlabel metal2 22218 16966 22218 16966 0 _0441_
rlabel metal1 21022 17204 21022 17204 0 _0442_
rlabel metal1 10304 5746 10304 5746 0 _0443_
rlabel metal2 10074 6324 10074 6324 0 _0444_
rlabel metal1 10350 5678 10350 5678 0 _0445_
rlabel metal1 11408 4794 11408 4794 0 _0446_
rlabel metal2 17986 25568 17986 25568 0 _0447_
rlabel metal1 17894 24820 17894 24820 0 _0448_
rlabel metal2 19274 24854 19274 24854 0 _0449_
rlabel metal1 18630 25330 18630 25330 0 _0450_
rlabel metal1 16790 23834 16790 23834 0 _0451_
rlabel metal2 15686 24480 15686 24480 0 _0452_
rlabel metal1 15870 24208 15870 24208 0 _0453_
rlabel metal1 15364 23698 15364 23698 0 _0454_
rlabel metal1 15226 24752 15226 24752 0 _0455_
rlabel metal1 15134 24718 15134 24718 0 _0456_
rlabel metal2 15594 23460 15594 23460 0 _0457_
rlabel metal1 14030 23698 14030 23698 0 _0458_
rlabel metal2 15226 23358 15226 23358 0 _0459_
rlabel metal1 13386 23698 13386 23698 0 _0460_
rlabel metal2 13018 24548 13018 24548 0 _0461_
rlabel metal2 14214 12784 14214 12784 0 clk
rlabel metal1 5658 23018 5658 23018 0 clknet_0_clk
rlabel metal1 2714 5712 2714 5712 0 clknet_4_0_0_clk
rlabel metal1 20332 6834 20332 6834 0 clknet_4_10_0_clk
rlabel metal1 26956 18190 26956 18190 0 clknet_4_11_0_clk
rlabel metal1 14766 18326 14766 18326 0 clknet_4_12_0_clk
rlabel metal2 15042 24752 15042 24752 0 clknet_4_13_0_clk
rlabel metal1 17388 25262 17388 25262 0 clknet_4_14_0_clk
rlabel metal1 19918 29104 19918 29104 0 clknet_4_15_0_clk
rlabel metal1 1656 15538 1656 15538 0 clknet_4_1_0_clk
rlabel metal1 12972 6222 12972 6222 0 clknet_4_2_0_clk
rlabel metal2 9246 13838 9246 13838 0 clknet_4_3_0_clk
rlabel metal2 1886 20366 1886 20366 0 clknet_4_4_0_clk
rlabel metal2 6854 23936 6854 23936 0 clknet_4_5_0_clk
rlabel metal1 9062 21590 9062 21590 0 clknet_4_6_0_clk
rlabel metal1 11500 24786 11500 24786 0 clknet_4_7_0_clk
rlabel metal1 16698 12750 16698 12750 0 clknet_4_8_0_clk
rlabel metal1 18722 17714 18722 17714 0 clknet_4_9_0_clk
rlabel metal1 18216 15334 18216 15334 0 e1.edge_d
rlabel metal1 3496 16626 3496 16626 0 e1.intermediate
rlabel metal1 9062 15946 9062 15946 0 e1.sync
rlabel metal1 9706 24582 9706 24582 0 e2.edge_d
rlabel metal1 2944 27506 2944 27506 0 e2.intermediate
rlabel metal1 6394 24820 6394 24820 0 e2.sync
rlabel metal1 26496 29138 26496 29138 0 net1
rlabel metal1 28290 18734 28290 18734 0 net10
rlabel metal1 11224 22406 11224 22406 0 net100
rlabel metal1 9798 22542 9798 22542 0 net101
rlabel metal1 19872 27302 19872 27302 0 net102
rlabel metal1 12236 22610 12236 22610 0 net103
rlabel metal1 5014 16490 5014 16490 0 net104
rlabel metal1 14582 27030 14582 27030 0 net105
rlabel metal1 16008 28050 16008 28050 0 net106
rlabel metal1 3358 20502 3358 20502 0 net107
rlabel metal1 12006 12954 12006 12954 0 net108
rlabel metal1 15686 28594 15686 28594 0 net109
rlabel metal1 25622 2414 25622 2414 0 net11
rlabel metal1 4600 7854 4600 7854 0 net110
rlabel metal1 12650 27506 12650 27506 0 net111
rlabel metal1 3358 17102 3358 17102 0 net112
rlabel metal1 9844 27506 9844 27506 0 net113
rlabel metal1 7774 25874 7774 25874 0 net114
rlabel metal2 19182 29478 19182 29478 0 net115
rlabel metal1 10994 29138 10994 29138 0 net116
rlabel metal1 24058 13770 24058 13770 0 net117
rlabel metal1 16330 22610 16330 22610 0 net118
rlabel metal2 9798 28968 9798 28968 0 net119
rlabel metal1 27370 21862 27370 21862 0 net12
rlabel metal1 6946 28594 6946 28594 0 net120
rlabel metal1 5934 26316 5934 26316 0 net121
rlabel metal1 3266 28628 3266 28628 0 net122
rlabel metal1 22678 29172 22678 29172 0 net123
rlabel metal1 23644 27438 23644 27438 0 net124
rlabel metal2 6946 25262 6946 25262 0 net125
rlabel metal1 7268 24174 7268 24174 0 net126
rlabel metal1 26726 7922 26726 7922 0 net127
rlabel metal2 26174 9180 26174 9180 0 net128
rlabel metal1 25438 17714 25438 17714 0 net129
rlabel metal1 1886 3502 1886 3502 0 net13
rlabel metal1 14490 8806 14490 8806 0 net130
rlabel metal2 22218 27608 22218 27608 0 net131
rlabel metal1 25622 14994 25622 14994 0 net132
rlabel metal2 26082 10846 26082 10846 0 net133
rlabel metal1 22770 7446 22770 7446 0 net134
rlabel metal1 10534 5270 10534 5270 0 net135
rlabel metal1 23966 7446 23966 7446 0 net136
rlabel metal1 25300 18054 25300 18054 0 net137
rlabel metal1 1886 2414 1886 2414 0 net14
rlabel metal2 21942 30022 21942 30022 0 net15
rlabel metal1 24886 22746 24886 22746 0 net16
rlabel metal2 1518 23375 1518 23375 0 net17
rlabel metal1 6394 30226 6394 30226 0 net18
rlabel metal1 15548 3706 15548 3706 0 net19
rlabel metal1 1564 16218 1564 16218 0 net2
rlabel metal1 1886 26554 1886 26554 0 net20
rlabel metal1 17963 2890 17963 2890 0 net21
rlabel metal1 5405 2414 5405 2414 0 net22
rlabel metal1 7314 2414 7314 2414 0 net23
rlabel metal2 3542 26220 3542 26220 0 net24
rlabel metal1 24702 6426 24702 6426 0 net25
rlabel metal1 14582 2346 14582 2346 0 net26
rlabel metal1 28566 26962 28566 26962 0 net27
rlabel metal2 20102 6579 20102 6579 0 net28
rlabel metal2 1518 12835 1518 12835 0 net29
rlabel metal1 1656 29206 1656 29206 0 net3
rlabel metal1 18814 4454 18814 4454 0 net30
rlabel metal1 20516 6426 20516 6426 0 net31
rlabel metal2 23874 14144 23874 14144 0 net32
rlabel metal2 13294 13226 13294 13226 0 net33
rlabel metal1 19780 14314 19780 14314 0 net34
rlabel metal2 7130 5440 7130 5440 0 net35
rlabel metal1 13018 14423 13018 14423 0 net36
rlabel metal1 3719 24854 3719 24854 0 net37
rlabel metal1 9437 24786 9437 24786 0 net38
rlabel metal1 20194 17748 20194 17748 0 net39
rlabel metal1 16560 2482 16560 2482 0 net4
rlabel metal2 15778 15266 15778 15266 0 net40
rlabel metal2 9062 28832 9062 28832 0 net41
rlabel metal1 2806 16184 2806 16184 0 net42
rlabel metal1 2484 25126 2484 25126 0 net43
rlabel metal1 7958 24718 7958 24718 0 net44
rlabel metal1 13478 15912 13478 15912 0 net45
rlabel metal1 17434 18768 17434 18768 0 net46
rlabel metal1 18216 17170 18216 17170 0 net47
rlabel metal1 14950 19380 14950 19380 0 net48
rlabel metal1 16698 9588 16698 9588 0 net49
rlabel metal2 9890 25823 9890 25823 0 net5
rlabel metal1 17342 20502 17342 20502 0 net50
rlabel metal1 16652 12818 16652 12818 0 net51
rlabel metal1 15824 11118 15824 11118 0 net52
rlabel metal1 11914 15538 11914 15538 0 net53
rlabel metal1 7360 11118 7360 11118 0 net54
rlabel metal1 15732 16082 15732 16082 0 net55
rlabel metal2 6854 6562 6854 6562 0 net56
rlabel metal1 15042 17238 15042 17238 0 net57
rlabel metal1 5934 12920 5934 12920 0 net58
rlabel metal1 7314 19414 7314 19414 0 net59
rlabel via2 2254 11747 2254 11747 0 net6
rlabel metal1 10120 18258 10120 18258 0 net60
rlabel metal1 9890 13940 9890 13940 0 net61
rlabel metal1 7130 14314 7130 14314 0 net62
rlabel metal1 14398 20400 14398 20400 0 net63
rlabel metal1 17986 8874 17986 8874 0 net64
rlabel metal1 6394 19856 6394 19856 0 net65
rlabel metal1 11592 14994 11592 14994 0 net66
rlabel metal1 3818 10540 3818 10540 0 net67
rlabel metal1 12282 12852 12282 12852 0 net68
rlabel metal1 14812 12206 14812 12206 0 net69
rlabel metal1 28336 19686 28336 19686 0 net7
rlabel metal1 9246 20026 9246 20026 0 net70
rlabel metal1 9890 16116 9890 16116 0 net71
rlabel metal2 14122 16762 14122 16762 0 net72
rlabel metal1 5060 6698 5060 6698 0 net73
rlabel metal1 7222 16082 7222 16082 0 net74
rlabel metal1 6762 22644 6762 22644 0 net75
rlabel via2 12098 19805 12098 19805 0 net76
rlabel metal1 6256 18734 6256 18734 0 net77
rlabel metal1 14904 13906 14904 13906 0 net78
rlabel metal1 4692 10642 4692 10642 0 net79
rlabel metal2 17664 26180 17664 26180 0 net8
rlabel metal1 13386 18394 13386 18394 0 net80
rlabel metal1 5060 9554 5060 9554 0 net81
rlabel metal1 3818 11152 3818 11152 0 net82
rlabel metal1 6670 6426 6670 6426 0 net83
rlabel metal2 7498 6596 7498 6596 0 net84
rlabel metal1 12880 19346 12880 19346 0 net85
rlabel metal1 10258 20434 10258 20434 0 net86
rlabel metal1 15962 20944 15962 20944 0 net87
rlabel metal1 4002 8500 4002 8500 0 net88
rlabel metal1 4646 22406 4646 22406 0 net89
rlabel metal1 28658 2414 28658 2414 0 net9
rlabel metal1 4922 17136 4922 17136 0 net90
rlabel metal1 5934 16762 5934 16762 0 net91
rlabel metal1 10626 19754 10626 19754 0 net92
rlabel metal1 9338 22678 9338 22678 0 net93
rlabel metal2 8510 21726 8510 21726 0 net94
rlabel metal2 4002 17884 4002 17884 0 net95
rlabel metal1 5934 21590 5934 21590 0 net96
rlabel metal1 4600 21454 4600 21454 0 net97
rlabel metal1 10718 16490 10718 16490 0 net98
rlabel metal2 9706 18326 9706 18326 0 net99
rlabel metal1 28382 30260 28382 30260 0 nrst
rlabel metal2 14858 959 14858 959 0 out_0[0]
rlabel metal1 9982 30294 9982 30294 0 out_0[1]
rlabel metal3 820 11628 820 11628 0 out_0[2]
rlabel via2 29118 11067 29118 11067 0 out_0[3]
rlabel metal1 17618 30090 17618 30090 0 out_0[4]
rlabel metal2 29670 1554 29670 1554 0 out_0[5]
rlabel metal1 29256 18938 29256 18938 0 out_0[6]
rlabel metal2 25806 823 25806 823 0 out_1[0]
rlabel via2 29026 22491 29026 22491 0 out_1[1]
rlabel metal3 820 3468 820 3468 0 out_1[2]
rlabel metal2 46 1520 46 1520 0 out_1[3]
rlabel metal2 21298 31154 21298 31154 0 out_1[4]
rlabel metal1 25576 30294 25576 30294 0 out_1[5]
rlabel metal3 751 23188 751 23188 0 out_1[6]
rlabel metal2 6762 31195 6762 31195 0 out_2[0]
rlabel metal2 21942 959 21942 959 0 out_2[1]
rlabel metal3 820 27268 820 27268 0 out_2[2]
rlabel via2 29026 2805 29026 2805 0 out_2[3]
rlabel metal2 3266 1520 3266 1520 0 out_2[4]
rlabel metal2 7130 1520 7130 1520 0 out_2[5]
rlabel metal1 2898 30090 2898 30090 0 out_2[6]
rlabel metal3 29494 6868 29494 6868 0 out_3[0]
rlabel metal2 10994 1095 10994 1095 0 out_3[1]
rlabel metal2 29026 26673 29026 26673 0 out_3[2]
rlabel metal1 28980 30158 28980 30158 0 out_3[3]
rlabel metal3 751 19788 751 19788 0 out_3[4]
rlabel metal1 14122 30090 14122 30090 0 out_3[5]
rlabel metal2 18722 823 18722 823 0 out_3[6]
rlabel metal3 820 15708 820 15708 0 pb_0
rlabel metal3 751 31348 751 31348 0 pb_1
rlabel metal3 29448 14348 29448 14348 0 time_done
<< properties >>
string FIXED_BBOX 0 0 30581 32725
<< end >>
