* NGSPICE file created from top_asic.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

.subckt top_asic VGND VPWR clk mode_out[0] mode_out[1] pb[0] pb[10] pb[11] pb[12]
+ pb[13] pb[14] pb[1] pb[2] pb[3] pb[4] pb[5] pb[6] pb[7] pb[8] pb[9] reset sigout
XANTENNA__09523__A2 _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06883_ genblk1\[6\].osc.clkdiv_C.cnt\[11\] _01484_ _01728_ _01734_ _01736_ VGND
+ VGND VPWR VPWR _01737_ sky130_fd_sc_hd__a2111o_1
X_09671_ _00006_ _04151_ net1174 VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__a21oi_1
X_08622_ _03251_ _03308_ _03327_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__nor3_1
X_08553_ genblk2\[6\].wave_shpr.div.fin_quo\[0\] genblk2\[6\].wave_shpr.div.fin_quo\[1\]
+ _02734_ _02261_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout162_A net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07504_ net18 net17 VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__nor2b_2
XANTENNA__11094__A1 _05055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08484_ _03188_ _03189_ _03190_ _02885_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07435_ _02173_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__buf_1
XFILLER_0_9_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11789__B genblk1\[9\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07366_ _02091_ _02120_ _02121_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__and3_1
X_09105_ genblk2\[0\].wave_shpr.div.acc\[10\] genblk2\[0\].wave_shpr.div.b1\[10\]
+ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__or2b_1
XFILLER_0_73_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06317_ genblk1\[0\].osc.clkdiv_C.cnt\[3\] _01274_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__and2_1
XANTENNA__10185__S _04507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07297_ _02062_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09036_ _03702_ _01432_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__nand2_8
XFILLER_0_130_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06248_ _01209_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold340 genblk2\[0\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__dlygate4sd3_1
X_06179_ net765 VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__inv_2
XANTENNA__10913__S _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold351 genblk2\[0\].wave_shpr.div.quo\[10\] VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 genblk2\[2\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold373 genblk2\[4\].wave_shpr.div.acc\[19\] VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 genblk2\[4\].wave_shpr.div.quo\[11\] VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07222__B1 _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09275__A _03804_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold395 genblk2\[7\].wave_shpr.div.quo\[14\] VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08610__C _02789_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09938_ genblk2\[2\].wave_shpr.div.acc\[21\] _04342_ _04343_ VGND VGND VPWR VPWR
+ _04344_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout75_A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09514__A2 _04043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09869_ genblk2\[2\].wave_shpr.div.acc\[4\] _04291_ _04214_ VGND VGND VPWR VPWR _04292_
+ sky130_fd_sc_hd__mux2_1
Xhold1040 genblk2\[6\].wave_shpr.div.b1\[6\] VGND VGND VPWR VPWR net1258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 genblk1\[11\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR net1269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 genblk2\[8\].wave_shpr.div.b1\[8\] VGND VGND VPWR VPWR net1280 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ genblk2\[0\].wave_shpr.div.i\[1\] genblk2\[0\].wave_shpr.div.i\[0\] genblk2\[0\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__a21o_1
Xhold1073 genblk2\[0\].wave_shpr.div.b1\[14\] VGND VGND VPWR VPWR net1291 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ clknet_leaf_119_clk _00211_ net146 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1084 genblk2\[10\].wave_shpr.div.b1\[17\] VGND VGND VPWR VPWR net1302 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 genblk2\[9\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net1313 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _05590_ _05562_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__or2b_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _05464_ genblk1\[9\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__and2_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13501_ clknet_leaf_86_clk net230 net180 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10713_ _02183_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__clkbuf_4
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _05565_ _05583_ _05584_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13432_ clknet_leaf_82_clk _00751_ net201 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12034__B1 _05816_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10644_ _03704_ net747 _04647_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__a21o_1
XANTENNA__07896__C _02365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_895 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10575_ _04769_ _04801_ _04802_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__a21o_1
X_13363_ clknet_leaf_3_clk _00682_ net53 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09450__A1 genblk2\[1\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12314_ _03942_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13294_ clknet_leaf_87_clk _00615_ net179 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12245_ genblk2\[11\].wave_shpr.div.fin_quo\[0\] _05982_ _00005_ VGND VGND VPWR VPWR
+ _05983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10899__A1 _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12176_ genblk2\[10\].wave_shpr.div.i\[1\] genblk2\[10\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _05918_ sky130_fd_sc_hd__nand2_1
X_11127_ _05181_ _05185_ _05186_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__a21o_1
XANTENNA__07417__B _02153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11058_ _04967_ _05013_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10009_ genblk2\[3\].wave_shpr.div.b1\[13\] genblk2\[3\].wave_shpr.div.acc\[13\]
+ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__and2b_1
XFILLER_0_64_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10520__B1 _04655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07220_ _01365_ _01189_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__or2_4
XFILLER_0_116_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12025__B1 _05817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07151_ _01928_ net34 _01944_ _01945_ _01950_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_42_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09079__B _01210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07082_ genblk1\[8\].osc.clkdiv_C.cnt\[5\] genblk1\[8\].osc.clkdiv_C.cnt\[4\] _01892_
+ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__and3_1
XANTENNA__06255__B2 genblk1\[0\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10339__B1 _03717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12193__B_N genblk2\[11\].wave_shpr.div.b1\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout105 net106 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_4
Xfanout116 net118 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_4
Xfanout127 net16 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_4
Xfanout138 net145 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_4
Xfanout149 net150 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
X_07984_ genblk2\[7\].wave_shpr.div.fin_quo\[6\] VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__inv_2
XANTENNA__06231__B _01192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09723_ genblk2\[2\].wave_shpr.div.b1\[15\] genblk2\[2\].wave_shpr.div.acc\[15\]
+ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__and2b_1
XANTENNA__09823__A _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06935_ net1180 _01775_ _01778_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[10\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__11303__A2 _05279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09654_ genblk2\[1\].wave_shpr.div.acc\[22\] _04139_ genblk2\[1\].wave_shpr.div.acc\[23\]
+ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__o21bai_1
XANTENNA__09542__B genblk1\[1\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06866_ net1115 _01719_ _01722_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06885__C _01439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08605_ genblk2\[3\].wave_shpr.div.fin_quo\[2\] _02467_ VGND VGND VPWR VPWR _03312_
+ sky130_fd_sc_hd__nand2_1
X_06797_ genblk1\[5\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__inv_2
X_09585_ genblk2\[1\].wave_shpr.div.b1\[6\] genblk2\[1\].wave_shpr.div.acc\[6\] VGND
+ VGND VPWR VPWR _04090_ sky130_fd_sc_hd__xor2_1
XFILLER_0_145_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ _03240_ _03242_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10814__A1 _04855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08467_ _03048_ _03049_ _03050_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07997__B _01360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07418_ _02160_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08398_ genblk1\[2\].osc.clkdiv_C.cnt\[15\] _01349_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07349_ genblk1\[11\].osc.clkdiv_C.cnt\[5\] genblk1\[11\].osc.clkdiv_C.cnt\[4\] _02101_
+ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__and3_1
X_10360_ _04648_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06125__C _01096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11790__A2 _02203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09019_ genblk2\[9\].wave_shpr.div.i\[1\] genblk2\[9\].wave_shpr.div.i\[0\] genblk2\[9\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__a21o_1
X_10291_ _04572_ _04601_ _04602_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__a21o_1
X_12030_ genblk2\[10\].wave_shpr.div.quo\[8\] _05813_ _05817_ net320 VGND VGND VPWR
+ VPWR _00957_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold170 _00388_ VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 PWM.counter\[7\] VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 genblk2\[0\].wave_shpr.div.quo\[17\] VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11542__A2 _05441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12932_ clknet_leaf_31_clk _00261_ net103 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ clknet_leaf_129_clk _00194_ net66 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _05582_ _05566_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__or2b_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ clknet_leaf_93_clk _00127_ net148 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ net746 _05623_ _05624_ _05613_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__a22o_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08474__A2 _02308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11676_ genblk2\[9\].wave_shpr.div.acc\[4\] genblk2\[9\].wave_shpr.div.b1\[4\] VGND
+ VGND VPWR VPWR _05568_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13415_ clknet_leaf_120_clk net488 net141 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10627_ _04840_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06237__A1 genblk1\[0\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13346_ clknet_leaf_6_clk _00667_ net49 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10558_ _04780_ _04784_ _04785_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13277_ clknet_leaf_12_clk _00598_ net54 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12334__A _03689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10489_ _04614_ _04566_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__nor2_1
X_12228_ _05930_ _05964_ _05965_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07147__B _01946_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12159_ genblk2\[10\].wave_shpr.div.acc\[21\] _05904_ VGND VGND VPWR VPWR _05907_
+ sky130_fd_sc_hd__xor2_1
X_06720_ _01600_ _01606_ _01607_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__and3_1
XANTENNA__07163__A genblk1\[9\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06651_ net1193 _01543_ _01546_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__o21a_1
X_09370_ net821 _03841_ _03839_ _03939_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__a22o_1
X_06582_ _01489_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__buf_8
XFILLER_0_59_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08321_ _02310_ _03027_ _02314_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10728__S _04821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09662__A1 _04042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08252_ _02738_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07610__B _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07673__B1 _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06507__A _01200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07203_ genblk1\[9\].osc.clkdiv_C.cnt\[16\] _01985_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08183_ _02850_ _02888_ _02889_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout125_A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07134_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01311_ _01923_ genblk1\[9\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09818__A _04250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11559__S _05417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07065_ genblk1\[8\].osc.clkdiv_C.cnt\[0\] _01211_ _01882_ VGND VGND VPWR VPWR _01883_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_113_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07967_ genblk1\[7\].osc.clkdiv_C.cnt\[12\] _01214_ _02673_ VGND VGND VPWR VPWR _02674_
+ sky130_fd_sc_hd__a21bo_1
XANTENNA__06896__B _01439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09706_ _04167_ _04184_ _04185_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__a21o_1
X_06918_ _01761_ _01767_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__nor2_1
X_07898_ genblk1\[8\].osc.clkdiv_C.cnt\[14\] _01309_ _01576_ genblk1\[8\].osc.clkdiv_C.cnt\[15\]
+ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__a2bb2o_1
X_09637_ _04006_ _04129_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06849_ _01693_ _01710_ _01711_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07900__A1 genblk1\[8\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09568_ _03974_ _03969_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout38_A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08519_ _02216_ _02552_ genblk2\[11\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR
+ _03226_ sky130_fd_sc_hd__and3_1
X_09499_ _04040_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11530_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__and2_1
XANTENNA__11460__A1 _01819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06417__A _01360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11461_ _05427_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06136__B net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13200_ clknet_leaf_115_clk _00523_ net134 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10412_ _04672_ genblk1\[4\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__and2_1
X_11392_ genblk2\[8\].wave_shpr.div.acc\[7\] genblk2\[8\].wave_shpr.div.b1\[7\] VGND
+ VGND VPWR VPWR _05368_ sky130_fd_sc_hd__or2b_1
XFILLER_0_61_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13131_ clknet_leaf_4_clk _00456_ net46 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10343_ _04638_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10274_ _04431_ genblk2\[4\].wave_shpr.div.acc\[1\] _04585_ VGND VGND VPWR VPWR _04586_
+ sky130_fd_sc_hd__a21o_1
X_13062_ clknet_leaf_29_clk net635 net95 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11515__A2 _05448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07719__B2 genblk1\[1\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12013_ _03726_ _05810_ _03735_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_136_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12915_ clknet_leaf_36_clk _00246_ net105 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ clknet_leaf_68_clk _00177_ net211 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07711__A net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ clknet_leaf_43_clk _00110_ net124 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11233__A _05245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ genblk2\[9\].wave_shpr.div.fin_quo\[3\] genblk2\[9\].wave_shpr.div.quo\[2\]
+ _00023_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11659_ _03690_ _05551_ _05552_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__nor3_1
XFILLER_0_126_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11203__A1 _03726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold906 genblk2\[11\].wave_shpr.div.i\[1\] VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 genblk2\[10\].wave_shpr.div.acc\[19\] VGND VGND VPWR VPWR net1135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13329_ clknet_leaf_25_clk _00650_ net91 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold928 genblk1\[6\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR net1146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 PWM.final_sample_in\[6\] VGND VGND VPWR VPWR net1157 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12064__A _03833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08870_ sig_norm.b1\[2\] VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__inv_2
X_07821_ genblk2\[1\].wave_shpr.div.fin_quo\[4\] _02521_ _02523_ _02527_ VGND VGND
+ VPWR VPWR _02528_ sky130_fd_sc_hd__a22o_1
XANTENNA__06394__B1 _01337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07605__B net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07752_ genblk1\[1\].osc.clkdiv_C.cnt\[16\] _01577_ genblk1\[1\].osc.clkdiv_C.cnt\[17\]
+ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__a21oi_4
X_06703_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01592_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__nand2_1
X_07683_ _01174_ genblk1\[10\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR _02390_
+ sky130_fd_sc_hd__nand2_1
X_09422_ genblk2\[1\].wave_shpr.div.b1\[8\] genblk2\[1\].wave_shpr.div.acc\[8\] VGND
+ VGND VPWR VPWR _03986_ sky130_fd_sc_hd__and2b_1
X_06634_ genblk1\[3\].osc.clkdiv_C.cnt\[6\] _01533_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09353_ net1175 _03903_ _03910_ _03928_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06565_ _01451_ _01476_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08304_ _02969_ _03003_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11442__A1 _05417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09284_ genblk2\[0\].wave_shpr.div.acc\[3\] _03875_ _03804_ VGND VGND VPWR VPWR _03876_
+ sky130_fd_sc_hd__mux2_1
X_06496_ genblk1\[2\].osc.clkdiv_C.cnt\[14\] genblk1\[2\].osc.clkdiv_C.cnt\[1\] _01327_
+ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08235_ _02592_ _02940_ _02941_ _02467_ genblk2\[3\].wave_shpr.div.fin_quo\[6\] VGND
+ VGND VPWR VPWR _02942_ sky130_fd_sc_hd__a32o_1
XFILLER_0_15_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08166_ genblk1\[3\].osc.clkdiv_C.cnt\[8\] _01423_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11745__A2 _05623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11289__S _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07117_ _01918_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[16\] sky130_fd_sc_hd__clkbuf_1
X_08097_ _02800_ _02801_ _02802_ _02803_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__or4b_1
XFILLER_0_101_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_868 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10953__B1 _05055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07048_ _01174_ _01182_ _01336_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09571__B1 _04047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08999_ _03679_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10961_ net620 _05062_ _05064_ genblk2\[6\].wave_shpr.div.quo\[12\] _05065_ VGND
+ VGND VPWR VPWR _00640_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12700_ clknet_leaf_89_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[13\] net172 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_2
X_13680_ clknet_leaf_63_clk _00993_ net190 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10484__A2 _04715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10892_ genblk2\[6\].wave_shpr.div.fin_quo\[6\] genblk2\[6\].wave_shpr.div.quo\[5\]
+ _00017_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__mux2_1
XANTENNA__07531__A _01155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12631_ clknet_leaf_18_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[16\] net112 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10236__A2 _04457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12562_ clknet_leaf_30_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[1\] net96 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__06147__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11513_ genblk2\[8\].wave_shpr.div.quo\[10\] _05448_ _05449_ net329 _05452_ VGND
+ VGND VPWR VPWR _00805_ sky130_fd_sc_hd__a221o_1
X_12493_ clknet_leaf_107_clk _00055_ net152 VGND VGND VPWR VPWR sig_norm.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11444_ genblk2\[8\].wave_shpr.div.fin_quo\[1\] net1331 _00021_ VGND VGND VPWR VPWR
+ _05419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11375_ _05353_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10944__B1 _05056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13114_ clknet_leaf_115_clk _00439_ net135 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10326_ genblk2\[4\].wave_shpr.div.fin_quo\[7\] net1263 _00013_ VGND VGND VPWR VPWR
+ _04631_ sky130_fd_sc_hd__mux2_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ clknet_leaf_128_clk _00372_ net67 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ genblk2\[4\].wave_shpr.div.acc\[13\] genblk2\[4\].wave_shpr.div.b1\[13\]
+ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__or2b_1
XFILLER_0_147_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10188_ _04403_ _04366_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__or2b_1
XANTENNA__10132__A _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10475__A2 _04715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12829_ clknet_leaf_64_clk _00162_ net189 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12059__A _03833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07160__B genblk1\[9\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06350_ _01268_ _01296_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06281_ genblk1\[0\].osc.clkdiv_C.cnt\[16\] _01242_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08020_ _02700_ _02702_ _02701_ _02726_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__and4_1
XFILLER_0_115_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold703 genblk2\[6\].wave_shpr.div.acc\[14\] VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 genblk2\[8\].wave_shpr.div.acc\[6\] VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold725 _00413_ VGND VGND VPWR VPWR net943 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 genblk2\[10\].wave_shpr.div.acc\[8\] VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold747 genblk2\[1\].wave_shpr.div.acc\[3\] VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 genblk2\[3\].wave_shpr.div.acc\[2\] VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06377__A_N _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09971_ genblk2\[3\].wave_shpr.div.acc\[11\] genblk2\[3\].wave_shpr.div.b1\[11\]
+ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__or2b_1
XFILLER_0_40_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold769 genblk2\[9\].wave_shpr.div.acc\[17\] VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__dlygate4sd3_1
X_08922_ net678 _03588_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09553__B1 _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08853_ _03501_ _03502_ _03500_ _03503_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07804_ genblk2\[0\].wave_shpr.div.fin_quo\[0\] genblk2\[0\].wave_shpr.div.fin_quo\[1\]
+ genblk2\[0\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__or3_1
X_08784_ _03474_ _03479_ _03490_ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__a21o_1
XANTENNA__09831__A _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07735_ genblk1\[1\].osc.clkdiv_C.cnt\[5\] _02433_ _01305_ genblk1\[1\].osc.clkdiv_C.cnt\[4\]
+ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__o22a_1
XANTENNA__09856__A1 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11572__S _05417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09550__B genblk1\[1\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07666_ _02368_ _02372_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _01190_ VGND VGND VPWR
+ VPWR _02373_ sky130_fd_sc_hd__a2bb2o_1
X_09405_ genblk2\[1\].wave_shpr.div.acc\[2\] genblk2\[1\].wave_shpr.div.b1\[2\] VGND
+ VGND VPWR VPWR _03969_ sky130_fd_sc_hd__or2b_1
X_06617_ _01522_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07597_ _02265_ genblk2\[9\].wave_shpr.div.fin_quo\[5\] _02303_ VGND VGND VPWR VPWR
+ _02304_ sky130_fd_sc_hd__or3b_1
XFILLER_0_48_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09336_ genblk2\[0\].wave_shpr.div.acc\[15\] _03915_ _03889_ VGND VGND VPWR VPWR
+ _03916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06548_ _01452_ _01464_ _01465_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_118_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10916__S _05042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09267_ _03838_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__inv_2
X_06479_ genblk1\[1\].osc.clkdiv_C.cnt\[16\] _01405_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__and2_1
X_08218_ _02900_ _02922_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__and2b_1
XFILLER_0_133_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09198_ _02005_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08149_ genblk1\[3\].osc.clkdiv_C.cnt\[2\] _01513_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10926__B1 _04647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11160_ genblk2\[7\].wave_shpr.div.acc\[23\] genblk2\[7\].wave_shpr.div.acc\[25\]
+ genblk2\[7\].wave_shpr.div.acc\[24\] genblk2\[7\].wave_shpr.div.acc\[26\] VGND VGND
+ VPWR VPWR _05220_ sky130_fd_sc_hd__or4_2
X_10111_ net634 _04461_ _04462_ genblk2\[3\].wave_shpr.div.quo\[13\] _04466_ VGND
+ VGND VPWR VPWR _00389_ sky130_fd_sc_hd__a221o_1
X_11091_ _05155_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10042_ _04430_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__clkbuf_1
Xhold30 _00975_ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 genblk2\[2\].wave_shpr.div.quo\[24\] VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 _00130_ VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold63 genblk2\[4\].wave_shpr.div.i\[4\] VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 genblk2\[1\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold85 _00721_ VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 _00647_ VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__dlygate4sd3_1
X_11993_ _05801_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13732_ clknet_leaf_45_clk _01043_ net121 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10944_ genblk2\[6\].wave_shpr.div.quo\[5\] _05052_ _05056_ net720 VGND VGND VPWR
+ VPWR _00632_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13663_ clknet_leaf_44_clk _00976_ net121 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10875_ genblk2\[6\].wave_shpr.div.acc\[19\] _05018_ VGND VGND VPWR VPWR _05019_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_38_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12614_ clknet_leaf_23_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[17\] net109 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13594_ clknet_leaf_72_clk _00909_ net216 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12545_ clknet_leaf_60_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[2\] net187 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_132_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_132_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__10090__B1 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12476_ clknet_leaf_106_clk _00038_ net151 VGND VGND VPWR VPWR sig_norm.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_5 _04242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11427_ _05361_ _05401_ _05402_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09783__B1 _04241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11358_ genblk2\[7\].wave_shpr.div.acc\[23\] _05219_ VGND VGND VPWR VPWR _05342_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10309_ genblk2\[4\].wave_shpr.div.acc\[23\] _04620_ VGND VGND VPWR VPWR _04621_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11289_ genblk2\[7\].wave_shpr.div.acc\[5\] _05290_ _05222_ VGND VGND VPWR VPWR _05291_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12342__A _03689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ clknet_leaf_113_clk _00355_ net131 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10696__A2 _02183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08966__S _01155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07520_ _02230_ PWM.final_sample_in\[5\] PWM.final_sample_in\[4\] _01163_ _02239_
+ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__o221a_1
X_07451_ genblk2\[6\].wave_shpr.div.i\[2\] genblk2\[6\].wave_shpr.div.i\[3\] genblk2\[6\].wave_shpr.div.i\[0\]
+ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_146_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06402_ genblk1\[1\].osc.clkdiv_C.cnt\[1\] _01340_ _01197_ _01341_ _01345_ VGND VGND
+ VPWR VPWR _01346_ sky130_fd_sc_hd__a221o_1
X_07382_ _02091_ _02131_ _02133_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__and3_1
X_09121_ genblk2\[0\].wave_shpr.div.b1\[3\] genblk2\[0\].wave_shpr.div.acc\[3\] VGND
+ VGND VPWR VPWR _03769_ sky130_fd_sc_hd__and2b_1
X_06333_ genblk1\[0\].osc.clkdiv_C.cnt\[9\] _01284_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__and2_1
XANTENNA__10736__S _04821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_123_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_123_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08274__B1 _02525_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06264_ _01225_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__buf_6
X_09052_ _03689_ _01242_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__nand2_2
XFILLER_0_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06515__A _01440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08003_ genblk1\[6\].osc.clkdiv_C.cnt\[12\] _01666_ _02709_ VGND VGND VPWR VPWR _02710_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_5_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06195_ net996 _01159_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__nor2_1
Xhold500 genblk1\[1\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold511 genblk2\[5\].wave_shpr.div.quo\[4\] VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold522 genblk2\[10\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__buf_1
Xhold533 genblk2\[8\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold544 genblk2\[11\].wave_shpr.div.acc\[9\] VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 _00579_ VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 genblk2\[4\].wave_shpr.div.acc\[15\] VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold577 genblk2\[8\].wave_shpr.div.quo\[4\] VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold588 genblk2\[6\].wave_shpr.div.acc\[9\] VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09954_ genblk2\[2\].wave_shpr.div.i\[1\] genblk2\[2\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _04354_ sky130_fd_sc_hd__nand2_1
Xhold599 genblk2\[9\].wave_shpr.div.i\[4\] VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__dlygate4sd3_1
X_08905_ _03596_ _03607_ _02248_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__a21oi_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _04188_ _04303_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10136__A1 _03819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _02509_ _02572_ _02518_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__o21ai_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08767_ _02798_ _03466_ _03468_ _03473_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__a31o_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11636__A1 _05449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07718_ _01360_ _01302_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__nand2_4
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ _03403_ _03357_ _03173_ _03402_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_67_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07649_ genblk2\[11\].wave_shpr.div.fin_quo\[5\] _02355_ VGND VGND VPWR VPWR _02356_
+ sky130_fd_sc_hd__nor2_1
X_10660_ net729 _04853_ _04857_ net745 VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09319_ net889 _03870_ _03877_ _03902_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10591_ genblk2\[5\].wave_shpr.div.acc\[23\] genblk2\[5\].wave_shpr.div.acc\[25\]
+ genblk2\[5\].wave_shpr.div.acc\[24\] genblk2\[5\].wave_shpr.div.acc\[26\] VGND VGND
+ VPWR VPWR _04819_ sky130_fd_sc_hd__or4_2
Xclkbuf_leaf_114_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_114_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_118_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_863 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12330_ _03689_ genblk1\[11\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR _06023_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06291__A2 _01240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12261_ genblk2\[1\].wave_shpr.div.b1\[0\] _01329_ _05802_ VGND VGND VPWR VPWR _05991_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11212_ _05245_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__clkbuf_4
X_12192_ genblk2\[11\].wave_shpr.div.acc\[12\] genblk2\[11\].wave_shpr.div.b1\[12\]
+ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__or2b_1
XANTENNA__08640__A _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11143_ genblk2\[7\].wave_shpr.div.b1\[11\] genblk2\[7\].wave_shpr.div.acc\[11\]
+ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09517__B1 _04047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11074_ net1001 _05119_ _05126_ _05144_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10025_ _02170_ genblk2\[3\].wave_shpr.div.busy _02172_ VGND VGND VPWR VPWR _04421_
+ sky130_fd_sc_hd__and3_2
XANTENNA__09471__A _01418_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10410__A _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11976_ genblk2\[10\].wave_shpr.div.fin_quo\[5\] genblk2\[10\].wave_shpr.div.quo\[4\]
+ _00003_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__mux2_1
X_13715_ clknet_leaf_21_clk _01026_ net97 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10927_ genblk2\[7\].wave_shpr.div.b1\[15\] _01365_ _05042_ VGND VGND VPWR VPWR _05048_
+ sky130_fd_sc_hd__mux2_1
X_13646_ clknet_leaf_48_clk _00959_ net114 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10858_ genblk2\[6\].wave_shpr.div.b1\[10\] genblk2\[6\].wave_shpr.div.acc\[10\]
+ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07059__A1 genblk1\[8\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07059__B2 genblk1\[8\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_105_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_105_clk sky130_fd_sc_hd__clkbuf_16
X_13577_ clknet_leaf_76_clk _00892_ net207 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10789_ net1345 _04941_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__nand2_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11241__A _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12528_ clknet_leaf_43_clk _00080_ net124 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12459_ clknet_leaf_104_clk _00032_ net153 VGND VGND VPWR VPWR PWM.final_sample_in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09220__A2 _03836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09508__B1 _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07166__A genblk1\[9\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07782__A2 _01241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06951_ genblk1\[6\].osc.clkdiv_C.cnt\[16\] _01787_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__or2_1
XANTENNA__11315__B1 _05283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10669__A2 _04858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09670_ _04045_ _04150_ _04152_ _04048_ net757 VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__a32o_1
X_06882_ genblk1\[6\].osc.clkdiv_C.cnt\[9\] _01732_ _01735_ genblk1\[6\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13338__RESET_B net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08621_ _03251_ _03308_ _03327_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__o21a_1
X_08552_ genblk2\[6\].wave_shpr.div.fin_quo\[0\] _02734_ genblk2\[6\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07503_ _02223_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__clkbuf_4
X_08483_ genblk2\[3\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07434_ _02171_ genblk2\[3\].wave_shpr.div.busy _02172_ VGND VGND VPWR VPWR _02173_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_91_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08247__B1 _02223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07365_ genblk1\[11\].osc.clkdiv_C.cnt\[7\] genblk1\[11\].osc.clkdiv_C.cnt\[6\] _02108_
+ genblk1\[11\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09104_ genblk2\[0\].wave_shpr.div.acc\[11\] genblk2\[0\].wave_shpr.div.b1\[11\]
+ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__or2b_1
XFILLER_0_17_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06316_ _01269_ _01274_ _01275_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07296_ _02028_ _02060_ _02061_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09035_ _02171_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__buf_6
X_06247_ _01208_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__buf_4
XANTENNA__09556__A _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold330 genblk2\[7\].wave_shpr.div.quo\[16\] VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__dlygate4sd3_1
X_06178_ _01144_ _01145_ _01147_ _01149_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__or4bb_4
Xhold341 _00126_ VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 _00134_ VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11297__S _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold363 _00335_ VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold374 genblk1\[0\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _00470_ VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 genblk2\[3\].wave_shpr.div.b1\[9\] VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07773__A2 _01556_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09937_ genblk2\[2\].wave_shpr.div.acc\[21\] genblk2\[2\].wave_shpr.div.acc\[20\]
+ _04210_ net22 VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__or4_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _04290_ _04180_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__xnor2_1
Xhold1030 genblk2\[6\].wave_shpr.div.b1\[12\] VGND VGND VPWR VPWR net1248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 genblk2\[9\].wave_shpr.div.fin_quo\[7\] VGND VGND VPWR VPWR net1259 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout68_A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1052 genblk2\[1\].wave_shpr.div.b1\[14\] VGND VGND VPWR VPWR net1270 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ _03461_ _03463_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__nor2_1
Xhold1063 genblk2\[4\].wave_shpr.div.b1\[13\] VGND VGND VPWR VPWR net1281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 genblk2\[10\].wave_shpr.div.b1\[11\] VGND VGND VPWR VPWR net1292 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ _04250_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__clkbuf_4
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 genblk2\[5\].wave_shpr.div.b1\[9\] VGND VGND VPWR VPWR net1303 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1096 genblk2\[0\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net1314 sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ net974 _05652_ _05653_ _05674_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__a22o_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11085__A2 _05057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _03693_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__clkbuf_4
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ clknet_leaf_87_clk _00817_ net179 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ net910 _04853_ _04857_ _04885_ VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__a22o_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ genblk2\[9\].wave_shpr.div.b1\[6\] genblk2\[9\].wave_shpr.div.acc\[6\] VGND
+ VGND VPWR VPWR _05584_ sky130_fd_sc_hd__and2b_1
XANTENNA__08635__A genblk2\[8\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13431_ clknet_leaf_82_clk _00750_ net201 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10643_ _04849_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12034__B2 genblk2\[10\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10045__B1 _03717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13362_ clknet_leaf_6_clk _00681_ net47 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10574_ genblk2\[5\].wave_shpr.div.b1\[11\] genblk2\[5\].wave_shpr.div.acc\[11\]
+ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10596__A1 genblk2\[5\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12313_ genblk2\[11\].wave_shpr.div.quo\[11\] _03947_ _03944_ net467 _06013_ VGND
+ VGND VPWR VPWR _01044_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13293_ clknet_leaf_87_clk _00614_ net179 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12337__A2 _03942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12244_ _05981_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__buf_4
XFILLER_0_121_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12175_ genblk2\[10\].wave_shpr.div.i\[1\] genblk2\[10\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _05917_ sky130_fd_sc_hd__or2_1
XANTENNA__10405__A _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11000__S _05023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11126_ genblk2\[7\].wave_shpr.div.b1\[2\] genblk2\[7\].wave_shpr.div.acc\[2\] VGND
+ VGND VPWR VPWR _05186_ sky130_fd_sc_hd__and2b_1
X_11057_ net1093 _05119_ _05126_ _05132_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__a22o_1
X_10008_ _04366_ _04402_ _04403_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11959_ _05731_ _05779_ _05780_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__a21o_1
XANTENNA__08477__B1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13629_ clknet_leaf_38_clk _00942_ net116 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_27_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07150_ genblk1\[9\].osc.clkdiv_C.cnt\[12\] _01799_ _01948_ _01949_ VGND VGND VPWR
+ VPWR _01950_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11784__B1 _03693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07081_ net1162 _01892_ _01894_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__06255__A2 _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10339__A1 _03732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12006__S _05802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout106 net107 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_2
XANTENNA__06512__B _01437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout117 net118 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
Xfanout128 net129 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11551__A3 _05417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07983_ _02683_ _02689_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__nand2_1
Xfanout139 net140 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06963__B1 _01238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09722_ _04159_ _04200_ _04201_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__a21o_1
X_06934_ net28 _01777_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__nor2_1
X_09653_ genblk2\[1\].wave_shpr.div.acc\[22\] _04139_ genblk2\[1\].wave_shpr.div.acc\[23\]
+ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__or3b_1
X_06865_ net27 _01721_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__nor2_1
X_08604_ _02261_ _03309_ _03310_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__or3b_1
X_09584_ net1260 _04076_ _04080_ _04089_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06796_ genblk1\[5\].osc.clkdiv_C.cnt\[13\] _01666_ _01667_ genblk1\[5\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08535_ _02314_ _03241_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10985__A _05074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08466_ _03170_ _03171_ _03172_ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__nand3_4
XFILLER_0_77_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07140__B1 _01328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07417_ _02157_ _02153_ genblk2\[1\].wave_shpr.div.busy VGND VGND VPWR VPWR _02160_
+ sky130_fd_sc_hd__and3b_2
XFILLER_0_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08397_ genblk1\[2\].osc.clkdiv_C.cnt\[14\] _01209_ _02425_ genblk1\[2\].osc.clkdiv_C.cnt\[13\]
+ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__a22o_1
X_07348_ _02107_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07279_ genblk1\[10\].osc.clkdiv_C.cnt\[10\] _02048_ _02050_ _02028_ VGND VGND VPWR
+ VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o211a_1
XFILLER_0_21_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10924__S _05042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09286__A _03838_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07994__A2 _01732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07132__A2_N _01578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09018_ genblk2\[9\].wave_shpr.div.busy net1039 genblk2\[9\].wave_shpr.div.i\[0\]
+ _03688_ _03690_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_60_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10290_ genblk2\[4\].wave_shpr.div.b1\[10\] genblk2\[4\].wave_shpr.div.acc\[10\]
+ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__and2b_1
XFILLER_0_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09196__A1 _03712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold160 genblk2\[5\].wave_shpr.div.quo\[16\] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 genblk2\[8\].wave_shpr.div.b1\[2\] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 genblk2\[7\].wave_shpr.div.quo\[18\] VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06422__B _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold193 _00141_ VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__dlygate4sd3_1
X_12931_ clknet_leaf_31_clk _00260_ net102 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_12862_ clknet_leaf_126_clk _00193_ net61 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ net999 _05652_ _05653_ _05661_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__a22o_1
XANTENNA__08459__B1 _02261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12793_ clknet_leaf_93_clk net559 net148 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _03693_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_139_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11675_ genblk2\[9\].wave_shpr.div.b1\[4\] genblk2\[9\].wave_shpr.div.acc\[4\] VGND
+ VGND VPWR VPWR _05567_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09959__B1 _04253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13414_ clknet_leaf_120_clk _00733_ net141 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10626_ net1258 net37 _04834_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13345_ clknet_leaf_6_clk _00666_ net49 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06237__A2 _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10557_ genblk2\[5\].wave_shpr.div.b1\[2\] genblk2\[5\].wave_shpr.div.acc\[2\] VGND
+ VGND VPWR VPWR _04785_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13276_ clknet_leaf_12_clk _00597_ net54 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_110_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10488_ net881 _04715_ _04722_ _04731_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11518__B1 _05449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12227_ genblk2\[11\].wave_shpr.div.b1\[12\] genblk2\[11\].wave_shpr.div.acc\[12\]
+ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__and2b_1
XANTENNA__08934__A1 _01099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12158_ net1087 _05876_ _05883_ _05906_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__a22o_1
X_11109_ genblk2\[7\].wave_shpr.div.acc\[12\] genblk2\[7\].wave_shpr.div.b1\[12\]
+ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__or2b_1
X_12089_ _05754_ _05743_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__nor2_1
X_06650_ _01523_ _01545_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06581_ _01187_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08320_ _03025_ _03026_ genblk2\[9\].wave_shpr.div.fin_quo\[4\] _02362_ VGND VGND
+ VPWR VPWR _03027_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_86_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07122__B1 _01328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08251_ _02946_ _02951_ _02957_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06507__B _01432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07202_ genblk1\[9\].osc.clkdiv_C.cnt\[15\] _01983_ _01986_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o21a_1
X_08182_ _02850_ _02888_ _02224_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11757__B1 _03694_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07133_ genblk1\[9\].osc.clkdiv_C.cnt\[7\] _01513_ _01929_ _01931_ _01932_ VGND VGND
+ VPWR VPWR _01933_ sky130_fd_sc_hd__a221o_1
XANTENNA__11221__A2 _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout118_A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07064_ _01874_ _01876_ _01877_ _01881_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__or4b_1
XFILLER_0_113_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09178__A1 _01342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08386__C1 _01441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07966_ genblk1\[7\].osc.clkdiv_C.cnt\[12\] _01214_ _01675_ genblk1\[7\].osc.clkdiv_C.cnt\[13\]
+ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__o22a_1
X_09705_ genblk2\[2\].wave_shpr.div.b1\[6\] genblk2\[2\].wave_shpr.div.acc\[6\] VGND
+ VGND VPWR VPWR _04185_ sky130_fd_sc_hd__and2b_1
XANTENNA__09045__S _03708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06917_ genblk1\[6\].osc.clkdiv_C.cnt\[4\] _01765_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__xnor2_1
X_07897_ _02603_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_94_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08153__A2 _01500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09636_ genblk2\[1\].wave_shpr.div.acc\[25\] genblk2\[1\].wave_shpr.div.acc\[26\]
+ _04009_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__nor3_2
X_06848_ genblk1\[5\].osc.clkdiv_C.cnt\[9\] _01708_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__nor2_1
XANTENNA__07900__A2 _01172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09567_ _04042_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__clkbuf_4
X_06779_ genblk1\[4\].osc.clkdiv_C.cnt\[16\] _01652_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__or2_1
X_08518_ _03136_ _03224_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__nor2_1
X_09498_ net1282 _01327_ _04039_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08449_ genblk2\[8\].wave_shpr.div.fin_quo\[3\] net30 _02639_ _02316_ VGND VGND VPWR
+ VPWR _03156_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07664__B2 _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11460_ genblk2\[9\].wave_shpr.div.b1\[1\] _01819_ _05237_ VGND VGND VPWR VPWR _05427_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11748__B1 _05624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10411_ net665 _04651_ _04663_ genblk2\[4\].wave_shpr.div.quo\[21\] _04674_ VGND
+ VGND VPWR VPWR _00481_ sky130_fd_sc_hd__a221o_1
XFILLER_0_150_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11391_ genblk2\[8\].wave_shpr.div.acc\[8\] genblk2\[8\].wave_shpr.div.b1\[8\] VGND
+ VGND VPWR VPWR _05367_ sky130_fd_sc_hd__or2b_1
XFILLER_0_104_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13130_ clknet_leaf_3_clk _00455_ net46 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07967__A2 _01214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07529__A _01099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10342_ genblk2\[5\].wave_shpr.div.b1\[8\] _01326_ _04637_ VGND VGND VPWR VPWR _04638_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13061_ clknet_leaf_29_clk net388 net95 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10273_ genblk2\[4\].wave_shpr.div.b1\[0\] _04583_ _04584_ VGND VGND VPWR VPWR _04585_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__12173__A0 _05815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13094__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07719__A2 _01309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12012_ net1086 VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_85_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_16
X_12914_ clknet_leaf_36_clk net367 net106 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap6 _01692_ VGND VGND VPWR VPWR net1355 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ clknet_leaf_68_clk _00176_ net194 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10239__A0 _04455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11514__A _04676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07711__B net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ clknet_leaf_43_clk _00109_ net124 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11727_ _05616_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__clkbuf_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11658_ genblk2\[8\].wave_shpr.div.i\[3\] _02197_ _05549_ VGND VGND VPWR VPWR _05552_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10609_ _04829_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11203__A2 _01869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11589_ genblk2\[8\].wave_shpr.div.acc\[9\] _05502_ _05493_ VGND VGND VPWR VPWR _05503_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold907 genblk2\[11\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07439__A _02147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13328_ clknet_leaf_25_clk _00649_ net86 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold918 genblk1\[9\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR net1136 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08080__A1 _01200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold929 genblk2\[8\].wave_shpr.div.b1\[12\] VGND VGND VPWR VPWR net1147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13259_ clknet_leaf_2_clk _00582_ net43 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07820_ _02526_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__06489__S _01210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06394__B2 genblk1\[1\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07751_ _02428_ _02450_ _02452_ _02457_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__a31o_4
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_76_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_16
X_06702_ _01171_ _01591_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__nand2_4
XFILLER_0_126_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06146__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07682_ genblk1\[10\].osc.clkdiv_C.cnt\[13\] _01246_ _02386_ VGND VGND VPWR VPWR
+ _02389_ sky130_fd_sc_hd__a21oi_1
X_09421_ _03964_ _03983_ _03984_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__a21o_1
X_06633_ genblk1\[3\].osc.clkdiv_C.cnt\[6\] _01533_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__and2_1
XANTENNA__06697__A2 _01436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09352_ genblk2\[0\].wave_shpr.div.acc\[19\] _03924_ _03927_ VGND VGND VPWR VPWR
+ _03928_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06564_ genblk1\[2\].osc.clkdiv_C.cnt\[14\] _01474_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08303_ _03007_ _03005_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__xnor2_1
X_09283_ _03768_ _03874_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__xnor2_1
X_06495_ genblk1\[2\].osc.clkdiv_C.cnt\[14\] genblk1\[2\].osc.clkdiv_C.cnt\[1\] _01327_
+ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__nor3_1
XFILLER_0_145_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08234_ _02885_ _02887_ genblk2\[3\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR
+ _02941_ sky130_fd_sc_hd__o21bai_1
XANTENNA__09829__A _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10474__S _04704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08165_ genblk1\[3\].osc.clkdiv_C.cnt\[10\] _01508_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__or2_1
XANTENNA__09548__B genblk1\[1\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07116_ _01886_ _01916_ _01917_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__and3b_1
X_08096_ _01174_ genblk1\[4\].osc.clkdiv_C.cnt\[15\] _01359_ VGND VGND VPWR VPWR _02803_
+ sky130_fd_sc_hd__or3_1
XANTENNA__06253__A _01213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07047_ _01336_ _01223_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__or2_2
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08998_ net1103 sig_norm.quo\[0\] _01154_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__mux2_1
XANTENNA__06700__B _01589_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07949_ _01172_ _02011_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_67_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08126__A2 _01340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10960_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout50_A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09619_ net1019 _04109_ _04113_ _04116_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__a22o_1
X_10891_ _05029_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12630_ clknet_leaf_18_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[15\] net82 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12561_ clknet_leaf_29_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[0\] net96 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__10338__B1_N _03733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06147__B net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11512_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12492_ clknet_leaf_107_clk _00054_ net153 VGND VGND VPWR VPWR sig_norm.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11443_ _05418_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11374_ genblk2\[7\].wave_shpr.div.i\[1\] genblk2\[7\].wave_shpr.div.i\[0\] genblk2\[7\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13113_ clknet_leaf_115_clk _00438_ net134 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10325_ _04630_ VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ clknet_leaf_128_clk _00371_ net67 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10256_ genblk2\[4\].wave_shpr.div.acc\[14\] genblk2\[4\].wave_shpr.div.b1\[14\]
+ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__or2b_1
XANTENNA__11509__A _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12104__S _05865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10187_ _04451_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_58_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07325__B1 _01925_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08522__C1 _02364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06679__A2 _01363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10880__A0 genblk2\[6\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07441__B _02153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12828_ clknet_leaf_62_clk _00161_ net190 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07160__C genblk1\[9\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ clknet_leaf_58_clk _00000_ net192 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06280_ _01241_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11188__A1 _01507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold704 genblk2\[8\].wave_shpr.div.acc\[9\] VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 genblk2\[0\].wave_shpr.div.acc\[22\] VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 genblk2\[10\].wave_shpr.div.acc\[15\] VGND VGND VPWR VPWR net944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold737 genblk2\[11\].wave_shpr.div.acc\[22\] VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold748 genblk2\[3\].wave_shpr.div.acc\[8\] VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ genblk2\[3\].wave_shpr.div.acc\[12\] genblk2\[3\].wave_shpr.div.b1\[12\]
+ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__or2b_1
XANTENNA__06603__A2 _01487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold759 genblk2\[10\].wave_shpr.div.acc\[5\] VGND VGND VPWR VPWR net977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08921_ net678 _02260_ _03619_ _03574_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__a22o_1
X_08852_ _03546_ _03551_ _03557_ _03558_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__a211oi_2
XANTENNA__07564__B1 _01732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07803_ net31 VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__buf_2
XFILLER_0_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08783_ _03478_ _03477_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_49_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout185_A net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07734_ _02435_ _02436_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__nor2_1
X_07665_ _02369_ _02370_ _02371_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__a21oi_1
X_09404_ genblk2\[1\].wave_shpr.div.acc\[3\] genblk2\[1\].wave_shpr.div.b1\[3\] VGND
+ VGND VPWR VPWR _03968_ sky130_fd_sc_hd__or2b_1
X_06616_ net1101 _01523_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
X_07596_ net32 VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__buf_2
XANTENNA__06248__A _01209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09335_ _03792_ _03914_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06547_ genblk1\[2\].osc.clkdiv_C.cnt\[7\] _01461_ genblk1\[2\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09266_ net578 _03835_ _03838_ genblk2\[0\].wave_shpr.div.quo\[24\] _03862_ VGND
+ VGND VPWR VPWR _00148_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06478_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] _01403_ _01406_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08217_ _02899_ _02923_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__or2b_1
XFILLER_0_132_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09197_ _03826_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11179__A1 _03831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08044__A1 _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08148_ genblk1\[3\].osc.clkdiv_C.cnt\[1\] _01496_ _01513_ genblk1\[3\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__a22o_1
XANTENNA__10926__A1 _03704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08079_ genblk1\[5\].osc.clkdiv_C.cnt\[11\] _01355_ _02760_ _02782_ _02785_ VGND
+ VGND VPWR VPWR _02786_ sky130_fd_sc_hd__o221a_1
XFILLER_0_30_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10110_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout98_A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11090_ _05054_ _05051_ genblk2\[6\].wave_shpr.div.i\[0\] VGND VGND VPWR VPWR _05155_
+ sky130_fd_sc_hd__mux2_1
X_10041_ genblk2\[3\].wave_shpr.div.fin_quo\[7\] genblk2\[3\].wave_shpr.div.quo\[6\]
+ _04422_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__mux2_1
Xhold20 _00810_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 genblk2\[5\].wave_shpr.div.quo\[14\] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 _00316_ VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 genblk2\[6\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 genblk2\[2\].wave_shpr.div.i\[4\] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 _00214_ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 genblk2\[9\].wave_shpr.div.quo\[15\] VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 genblk2\[2\].wave_shpr.div.quo\[15\] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ genblk2\[11\].wave_shpr.div.b1\[5\] _01855_ _05433_ VGND VGND VPWR VPWR _05801_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12300__B1 _06010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10943_ genblk2\[6\].wave_shpr.div.quo\[4\] _05052_ _05056_ net271 VGND VGND VPWR
+ VPWR _00631_ sky130_fd_sc_hd__a22o_1
X_13731_ clknet_leaf_45_clk net356 net121 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10874_ genblk2\[6\].wave_shpr.div.acc\[18\] _05017_ VGND VGND VPWR VPWR _05018_
+ sky130_fd_sc_hd__or2_1
X_13662_ clknet_leaf_45_clk net248 net121 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06158__A net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12613_ clknet_leaf_23_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[16\] net94 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_2
X_13593_ clknet_leaf_72_clk _00908_ net216 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12544_ clknet_leaf_60_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[1\] net192 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12475_ clknet_leaf_116_clk FSM.next_mode\[1\] net150 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_151_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10408__A _04672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11426_ genblk2\[8\].wave_shpr.div.b1\[14\] genblk2\[8\].wave_shpr.div.acc\[14\]
+ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_6 _04242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09232__B1 _03839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09783__A1 _03732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11357_ net873 _05251_ _05315_ _05341_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_830 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10308_ genblk2\[4\].wave_shpr.div.acc\[22\] _04619_ VGND VGND VPWR VPWR _04620_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07717__A net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11288_ _05289_ _05190_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__xnor2_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ clknet_leaf_113_clk _00354_ net131 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11239__A _05074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10239_ _04455_ _04451_ genblk2\[3\].wave_shpr.div.i\[0\] VGND VGND VPWR VPWR _04556_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07450_ _02184_ VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06521__B2 _01436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06401_ _01342_ genblk1\[1\].osc.clkdiv_C.cnt\[8\] _01344_ genblk1\[1\].osc.clkdiv_C.cnt\[13\]
+ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07381_ _02132_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09120_ _03761_ genblk2\[0\].wave_shpr.div.acc\[2\] _03767_ VGND VGND VPWR VPWR _03768_
+ sky130_fd_sc_hd__a21o_1
X_06332_ _01269_ _01284_ _01285_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__09379__A _03942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09051_ _03702_ _01257_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__nand2_1
X_06263_ _01175_ _01194_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08002_ genblk1\[6\].osc.clkdiv_C.cnt\[13\] _01675_ _01666_ genblk1\[6\].osc.clkdiv_C.cnt\[12\]
+ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__o22a_1
XFILLER_0_130_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06194_ PWM.counter\[3\] _01159_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold501 genblk2\[2\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09223__B1 _03840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold512 genblk2\[3\].wave_shpr.div.b1\[16\] VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09774__A1 _03831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold523 genblk2\[11\].wave_shpr.div.i\[2\] VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 genblk2\[1\].wave_shpr.div.acc\[0\] VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_13_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold545 genblk2\[4\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold556 genblk2\[1\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10384__A2 _04657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold567 genblk2\[11\].wave_shpr.div.acc\[11\] VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 genblk2\[3\].wave_shpr.div.acc\[9\] VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ genblk2\[2\].wave_shpr.div.i\[1\] genblk2\[2\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _04353_ sky130_fd_sc_hd__or2_1
Xhold589 genblk2\[9\].wave_shpr.div.acc\[11\] VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08904_ _03584_ _03592_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__xnor2_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _04189_ _04165_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__or2b_1
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ net8 _02744_ _03541_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__and3_1
XANTENNA__10988__A _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11884__A2 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08766_ _03470_ _03472_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__and2_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07717_ net7 _02364_ _02365_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__nand3_2
XANTENNA__10199__S _04507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ _03173_ _03402_ _03403_ _03357_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07648_ genblk2\[11\].wave_shpr.div.fin_quo\[4\] _02354_ VGND VGND VPWR VPWR _02355_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_95_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10927__S _05042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07579_ _02283_ _02284_ _02285_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__or3b_1
X_09318_ genblk2\[0\].wave_shpr.div.acc\[11\] _03901_ _03889_ VGND VGND VPWR VPWR
+ _03902_ sky130_fd_sc_hd__mux2_1
X_10590_ genblk2\[5\].wave_shpr.div.acc\[22\] _04817_ VGND VGND VPWR VPWR _04818_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09249_ _03707_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12260_ _05990_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11211_ _02193_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__clkbuf_4
X_12191_ genblk2\[11\].wave_shpr.div.acc\[13\] genblk2\[11\].wave_shpr.div.b1\[13\]
+ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__or2b_1
XFILLER_0_120_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11142_ _05171_ _05200_ _05201_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__a21o_1
XANTENNA__07240__A2 _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09517__A1 genblk2\[1\].wave_shpr.div.quo\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09517__B2 net292 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11073_ genblk2\[6\].wave_shpr.div.acc\[20\] _05142_ VGND VGND VPWR VPWR _05144_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__10127__A2 _04451_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10024_ _04419_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11975_ _05792_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08087__B _02789_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13714_ clknet_leaf_31_clk _01025_ net102 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10926_ _03704_ net484 _04647_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10857_ _04974_ _04999_ _05000_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__a21o_1
X_13645_ clknet_leaf_48_clk net433 net114 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10788_ genblk2\[5\].wave_shpr.div.acc\[20\] _04941_ VGND VGND VPWR VPWR _04943_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_54_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13576_ clknet_leaf_84_clk net1210 net202 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12527_ clknet_leaf_67_clk _00079_ net193 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10138__A _04480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12458_ clknet_leaf_104_clk _00031_ net155 VGND VGND VPWR VPWR PWM.final_sample_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11409_ _05370_ _05383_ _05384_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__a21o_1
X_12389_ _05960_ _06063_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07767__B1 _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09508__A1 genblk2\[1\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06950_ genblk1\[6\].osc.clkdiv_C.cnt\[15\] _01785_ _01788_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09508__B2 _04045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06881_ _01189_ _01678_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__or2_2
XFILLER_0_118_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08620_ _03313_ _03326_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08551_ _03256_ _03257_ VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__or2_2
X_07502_ _02222_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08482_ genblk2\[3\].wave_shpr.div.fin_quo\[1\] VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07433_ genblk2\[3\].wave_shpr.div.i\[1\] _02166_ genblk2\[3\].wave_shpr.div.i\[4\]
+ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_58_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout148_A net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07364_ _02119_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09103_ genblk2\[0\].wave_shpr.div.acc\[12\] genblk2\[0\].wave_shpr.div.b1\[12\]
+ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__or2b_1
X_06315_ genblk1\[0\].osc.clkdiv_C.cnt\[1\] genblk1\[0\].osc.clkdiv_C.cnt\[0\] genblk1\[0\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07295_ genblk1\[10\].osc.clkdiv_C.cnt\[16\] _02058_ VGND VGND VPWR VPWR _02061_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09034_ _03700_ _03703_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09837__A _04269_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06246_ _01207_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__buf_4
XFILLER_0_115_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold320 genblk2\[3\].wave_shpr.div.quo\[9\] VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__dlygate4sd3_1
X_06177_ _01140_ _01148_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold331 _00728_ VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold342 genblk2\[6\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09048__S _03708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold353 genblk2\[11\].wave_shpr.div.quo\[16\] VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold364 genblk2\[6\].wave_shpr.div.quo\[17\] VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 genblk2\[8\].wave_shpr.div.b1\[4\] VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold386 genblk2\[0\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 genblk2\[8\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07773__A3 _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09936_ genblk2\[2\].wave_shpr.div.acc\[20\] _04210_ net1351 VGND VGND VPWR VPWR
+ _04342_ sky130_fd_sc_hd__or3_1
XANTENNA__09572__A _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _04181_ _04169_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__or2b_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1020 genblk2\[0\].wave_shpr.div.b1\[3\] VGND VGND VPWR VPWR net1238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 genblk2\[10\].wave_shpr.div.b1\[3\] VGND VGND VPWR VPWR net1249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1042 genblk2\[1\].wave_shpr.div.acc\[6\] VGND VGND VPWR VPWR net1260 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ _03508_ _03519_ _03523_ _03524_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__o31a_1
Xhold1053 genblk2\[2\].wave_shpr.div.b1\[13\] VGND VGND VPWR VPWR net1271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1064 genblk2\[2\].wave_shpr.div.b1\[14\] VGND VGND VPWR VPWR net1282 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ net1054 _04248_ _04214_ _04251_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__a22o_1
Xhold1075 genblk2\[7\].wave_shpr.div.b1\[5\] VGND VGND VPWR VPWR net1293 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 genblk2\[2\].wave_shpr.div.b1\[10\] VGND VGND VPWR VPWR net1304 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 genblk2\[5\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net1315 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ genblk2\[8\].wave_shpr.div.fin_quo\[0\] _02309_ _02636_ VGND VGND VPWR VPWR
+ _03456_ sky130_fd_sc_hd__a21oi_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _02203_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__clkbuf_4
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08486__B2 _02592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07820__A _02526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10711_ genblk2\[5\].wave_shpr.div.acc\[1\] _04884_ _04821_ VGND VGND VPWR VPWR _04885_
+ sky130_fd_sc_hd__mux2_1
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _05566_ _05581_ _05582_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10642_ genblk2\[6\].wave_shpr.div.b1\[13\] _04645_ _04848_ VGND VGND VPWR VPWR _04849_
+ sky130_fd_sc_hd__mux2_1
X_13430_ clknet_leaf_82_clk net853 net201 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12034__A2 _05818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10045__A1 _03714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13361_ clknet_leaf_6_clk _00680_ net47 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10573_ _04770_ _04799_ _04800_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12312_ _05835_ genblk1\[11\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13292_ clknet_leaf_88_clk _00613_ net177 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12243_ genblk2\[11\].wave_shpr.div.acc\[25\] genblk2\[11\].wave_shpr.div.acc\[24\]
+ genblk2\[11\].wave_shpr.div.acc\[26\] _05980_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__or4_2
XFILLER_0_20_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12174_ _05916_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__clkbuf_1
X_11125_ _05033_ genblk2\[7\].wave_shpr.div.acc\[1\] _05184_ VGND VGND VPWR VPWR _05185_
+ sky130_fd_sc_hd__a21o_1
X_11056_ genblk2\[6\].wave_shpr.div.acc\[15\] _05131_ _05105_ VGND VGND VPWR VPWR
+ _05132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10007_ genblk2\[3\].wave_shpr.div.b1\[12\] genblk2\[3\].wave_shpr.div.acc\[12\]
+ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__and2b_1
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12112__S _05865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08098__A _01440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10520__A2 _04657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11958_ genblk2\[10\].wave_shpr.div.b1\[17\] genblk2\[10\].wave_shpr.div.acc\[17\]
+ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09674__B1 _03819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07730__A _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10909_ net1202 _04432_ _04848_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__mux2_1
X_11889_ genblk2\[9\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__inv_2
X_13628_ clknet_leaf_65_clk _00941_ net197 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12025__A2 _05813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13559_ clknet_leaf_85_clk _00874_ net184 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_07080_ genblk1\[8\].osc.clkdiv_C.cnt\[4\] _01892_ _01886_ VGND VGND VPWR VPWR _01894_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout107 net127 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_2
Xfanout118 net126 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__buf_2
XFILLER_0_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout129 net131 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
X_07982_ genblk2\[7\].wave_shpr.div.fin_quo\[4\] _02688_ VGND VGND VPWR VPWR _02689_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06963__A1 _01229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09721_ genblk2\[2\].wave_shpr.div.b1\[14\] genblk2\[2\].wave_shpr.div.acc\[14\]
+ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__and2b_1
X_06933_ genblk1\[6\].osc.clkdiv_C.cnt\[10\] genblk1\[6\].osc.clkdiv_C.cnt\[9\] _01773_
+ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__and3_1
X_09652_ net803 _04048_ _04113_ _04140_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__a22o_1
X_06864_ genblk1\[5\].osc.clkdiv_C.cnt\[15\] genblk1\[5\].osc.clkdiv_C.cnt\[14\] _01717_
+ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__and3_1
XANTENNA__10511__A2 _04657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08603_ _03188_ _02885_ _03189_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__o21ai_1
X_09583_ genblk2\[1\].wave_shpr.div.acc\[5\] _04088_ _04011_ VGND VGND VPWR VPWR _04089_
+ sky130_fd_sc_hd__mux2_1
X_06795_ _01325_ _01254_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__or2_2
X_08534_ genblk2\[9\].wave_shpr.div.fin_quo\[0\] _02526_ _02308_ genblk2\[9\].wave_shpr.div.fin_quo\[1\]
+ _02310_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__a221o_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08465_ _03153_ _03152_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07140__B2 genblk1\[9\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07416_ _02159_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08396_ genblk1\[2\].osc.clkdiv_C.cnt\[15\] _01349_ _01209_ genblk1\[2\].osc.clkdiv_C.cnt\[14\]
+ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_70_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10027__A1 _04420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11224__B1 _05250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07347_ _02092_ _02105_ _02106_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09567__A _04042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07278_ genblk1\[10\].osc.clkdiv_C.cnt\[10\] _02048_ VGND VGND VPWR VPWR _02050_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09017_ _03689_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__buf_8
XFILLER_0_131_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06229_ freq_div.state\[2\] VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06703__B _01592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold150 smpl_rt_clkdiv.clkDiv_inst.cnt\[3\] VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 genblk2\[0\].wave_shpr.div.quo\[7\] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 genblk2\[9\].wave_shpr.div.b1\[15\] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 genblk2\[3\].wave_shpr.div.quo\[7\] VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold194 genblk2\[11\].wave_shpr.div.quo\[24\] VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__dlygate4sd3_1
X_09919_ _04329_ _04204_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08156__B1 _01576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12930_ clknet_leaf_116_clk _00009_ net150 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ clknet_leaf_129_clk _00192_ net64 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ genblk2\[9\].wave_shpr.div.acc\[4\] _05660_ _05613_ VGND VGND VPWR VPWR _05661_
+ sky130_fd_sc_hd__mux2_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ clknet_leaf_91_clk _00125_ net148 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11743_ _02203_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__clkbuf_4
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11674_ genblk2\[9\].wave_shpr.div.acc\[5\] genblk2\[9\].wave_shpr.div.b1\[5\] VGND
+ VGND VPWR VPWR _05566_ sky130_fd_sc_hd__or2b_1
XANTENNA__07682__A2 _01246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09959__A1 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11215__B1 _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13413_ clknet_leaf_120_clk net528 net142 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10625_ _04839_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06890__B1 _01739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10556_ _04633_ genblk2\[5\].wave_shpr.div.acc\[1\] _04783_ VGND VGND VPWR VPWR _04784_
+ sky130_fd_sc_hd__a21o_1
X_13344_ clknet_leaf_7_clk _00665_ net49 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10487_ genblk2\[4\].wave_shpr.div.acc\[15\] _04730_ _04704_ VGND VGND VPWR VPWR
+ _04731_ sky130_fd_sc_hd__mux2_1
X_13275_ clknet_leaf_12_clk _00596_ net54 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_121_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12226_ _05931_ _05962_ _05963_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12157_ _05904_ _05905_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__or2_1
X_11108_ genblk2\[7\].wave_shpr.div.acc\[13\] genblk2\[7\].wave_shpr.div.b1\[13\]
+ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__or2b_1
X_12088_ net868 _05844_ _05850_ _05853_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__a22o_1
XANTENNA__08147__B1 _01519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11039_ net838 _05086_ _05093_ _05118_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06580_ genblk1\[3\].osc.clkdiv_C.cnt\[12\] _01344_ genblk1\[3\].osc.clkdiv_C.cnt\[13\]
+ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07122__B2 genblk1\[9\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08250_ _02955_ _02956_ _02604_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07673__A2 _02001_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07201_ _01952_ _01985_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08181_ genblk2\[3\].wave_shpr.div.fin_quo\[5\] _02885_ _02887_ VGND VGND VPWR VPWR
+ _02888_ sky130_fd_sc_hd__or3b_1
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07132_ genblk1\[9\].osc.clkdiv_C.cnt\[16\] _01578_ _01349_ genblk1\[9\].osc.clkdiv_C.cnt\[15\]
+ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09387__A _03726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07063_ _01441_ _01878_ genblk1\[8\].osc.clkdiv_C.cnt\[2\] _01880_ VGND VGND VPWR
+ VPWR _01881_ sky130_fd_sc_hd__a31o_1
XFILLER_0_113_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10980__A2 _05051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07965_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01577_ _01675_ genblk1\[7\].osc.clkdiv_C.cnt\[13\]
+ _02671_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__a221o_1
X_09704_ _04168_ _04182_ _04183_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__a21o_1
XANTENNA__10061__A _03701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06916_ _01761_ _01765_ _01766_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
X_07896_ net14 net136 _02365_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__and3_1
X_09635_ net664 _04109_ _04113_ _04128_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06847_ genblk1\[5\].osc.clkdiv_C.cnt\[9\] _01708_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__and2_1
X_06778_ _01650_ _01648_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__nor2_1
X_09566_ net990 _04043_ _04047_ _04075_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__a22o_1
X_08517_ _03219_ _03223_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09497_ _03701_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07113__A1 genblk1\[8\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08185__B _02539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08448_ _02638_ _02639_ genblk2\[8\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR
+ _03155_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07664__A2 _02336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08379_ genblk1\[2\].osc.clkdiv_C.cnt\[6\] _01433_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__nand2_1
X_10410_ _04058_ _01644_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11390_ genblk2\[8\].wave_shpr.div.acc\[9\] genblk2\[8\].wave_shpr.div.b1\[9\] VGND
+ VGND VPWR VPWR _05366_ sky130_fd_sc_hd__or2b_1
XANTENNA__09810__B1 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10341_ _03701_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__buf_4
XFILLER_0_131_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13060_ clknet_leaf_21_clk _00387_ net95 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10272_ genblk2\[4\].wave_shpr.div.b1\[1\] genblk2\[4\].wave_shpr.div.acc\[1\] VGND
+ VGND VPWR VPWR _04584_ sky130_fd_sc_hd__xor2_1
X_12011_ _03687_ net424 _03717_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__a21bo_1
X_12913_ clknet_leaf_34_clk _00244_ net106 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap7 _01760_ VGND VGND VPWR VPWR net1356 sky130_fd_sc_hd__buf_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ clknet_leaf_116_clk _00007_ net150 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10239__A1 _04451_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ clknet_leaf_41_clk _00108_ net123 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07104__A1 genblk1\[8\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08095__B _01196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06608__B _01210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11726_ genblk2\[9\].wave_shpr.div.fin_quo\[2\] net1313 _00023_ VGND VGND VPWR VPWR
+ _05616_ sky130_fd_sc_hd__mux2_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11657_ _00020_ _05549_ net1164 VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10608_ genblk2\[5\].wave_shpr.div.fin_quo\[7\] net1344 _00015_ VGND VGND VPWR VPWR
+ _04829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09801__B1 _04252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11588_ _05391_ _05501_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold908 sig_norm.quo\[1\] VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__dlygate4sd3_1
X_13327_ clknet_leaf_25_clk net568 net86 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold919 genblk2\[2\].wave_shpr.div.acc\[2\] VGND VGND VPWR VPWR net1137 sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ genblk2\[5\].wave_shpr.div.acc\[13\] genblk2\[5\].wave_shpr.div.b1\[13\]
+ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13258_ clknet_leaf_2_clk _00581_ net51 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12209_ genblk2\[11\].wave_shpr.div.b1\[3\] genblk2\[11\].wave_shpr.div.acc\[3\]
+ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__and2b_1
X_13189_ clknet_leaf_122_clk _00512_ net78 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06394__A2 _01210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07750_ _02428_ _02453_ _02452_ _02456_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__a31o_1
X_06701_ _01173_ _01175_ _01191_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__or3b_4
X_07681_ _02387_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06632_ _01523_ _01533_ _01534_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
X_09420_ genblk2\[1\].wave_shpr.div.b1\[7\] genblk2\[1\].wave_shpr.div.acc\[7\] VGND
+ VGND VPWR VPWR _03984_ sky130_fd_sc_hd__and2b_1
XFILLER_0_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09351_ _03800_ net23 VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__nor2_1
X_06563_ net1166 _01472_ _01475_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09096__A1 _01490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08302_ _02602_ _02924_ _02927_ _03008_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09282_ _03769_ _03760_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__or2b_1
XFILLER_0_145_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06494_ _01242_ _01223_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__nor2_2
XFILLER_0_74_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08233_ _02887_ _02885_ genblk2\[3\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR
+ _02940_ sky130_fd_sc_hd__or3b_1
XFILLER_0_144_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08164_ _01181_ genblk1\[3\].osc.clkdiv_C.cnt\[9\] _01182_ VGND VGND VPWR VPWR _02871_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07115_ genblk1\[8\].osc.clkdiv_C.cnt\[16\] _01914_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08095_ _01650_ _01196_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06253__B _01214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10953__A2 _05057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09845__A _04269_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07046_ genblk1\[8\].osc.clkdiv_C.cnt\[13\] _01328_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09056__S _03708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08997_ _03678_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__clkbuf_1
X_07948_ genblk1\[7\].osc.clkdiv_C.cnt\[7\] _01947_ _02652_ _02653_ _02654_ VGND VGND
+ VPWR VPWR _02655_ sky130_fd_sc_hd__o221a_1
X_07879_ _02548_ _02561_ _02585_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__or3_2
XANTENNA__06970__A2_N _01805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09618_ genblk2\[1\].wave_shpr.div.acc\[13\] _04115_ _04095_ VGND VGND VPWR VPWR
+ _04116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout43_A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10890_ genblk2\[6\].wave_shpr.div.fin_quo\[5\] net720 _00017_ VGND VGND VPWR VPWR
+ _05029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09549_ genblk2\[1\].wave_shpr.div.quo\[21\] _04052_ _04053_ net257 _04065_ VGND
+ VGND VPWR VPWR _00228_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12560_ clknet_leaf_57_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[17\] net181 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11511_ net329 _05448_ _05449_ net450 _05451_ VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12491_ clknet_leaf_107_clk _00053_ net158 VGND VGND VPWR VPWR sig_norm.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11442_ genblk2\[8\].wave_shpr.div.fin_quo\[0\] _05417_ _00021_ VGND VGND VPWR VPWR
+ _05418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08598__B1 _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11373_ genblk2\[7\].wave_shpr.div.i\[1\] genblk2\[7\].wave_shpr.div.i\[0\] genblk2\[7\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__a21o_1
XANTENNA_hold976_A genblk1\[9\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10944__A2 _05052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13112_ clknet_leaf_115_clk _00437_ net134 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10324_ genblk2\[4\].wave_shpr.div.fin_quo\[6\] genblk2\[4\].wave_shpr.div.quo\[5\]
+ _00013_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13043_ clknet_leaf_128_clk _00370_ net66 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10255_ genblk2\[4\].wave_shpr.div.acc\[15\] genblk2\[4\].wave_shpr.div.b1\[15\]
+ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__or2b_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09562__A2 _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10186_ net942 _04486_ _04490_ _04517_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__a22o_1
XANTENNA__08522__B1 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12827_ clknet_leaf_62_clk _00160_ net190 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10880__A1 _05023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12758_ clknet_leaf_52_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[17\] net110 VGND
+ VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07628__A2 _01256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10632__A1 _01923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11709_ _05557_ _05599_ _05600_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12689_ clknet_leaf_53_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[2\] net174 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold705 genblk2\[7\].wave_shpr.div.acc\[20\] VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold716 genblk2\[0\].wave_shpr.div.acc\[10\] VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 genblk2\[10\].wave_shpr.div.acc\[14\] VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold738 genblk2\[0\].wave_shpr.div.acc\[9\] VGND VGND VPWR VPWR net956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold749 genblk2\[9\].wave_shpr.div.acc\[13\] VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08920_ _03588_ _03602_ _03618_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__o21ai_1
X_08851_ _03555_ _03556_ _03552_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09553__A2 _04042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07802_ _02221_ net31 VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__nor2_2
X_08782_ _03487_ _03488_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__nand2_1
XANTENNA__09604__S _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11648__A0 _05444_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07733_ _02430_ _02431_ _02432_ _02434_ _02439_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07664_ genblk1\[10\].osc.clkdiv_C.cnt\[6\] _02336_ _01794_ genblk1\[10\].osc.clkdiv_C.cnt\[5\]
+ _01182_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__a32o_1
XFILLER_0_95_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09403_ genblk2\[1\].wave_shpr.div.acc\[4\] genblk2\[1\].wave_shpr.div.b1\[4\] VGND
+ VGND VPWR VPWR _03967_ sky130_fd_sc_hd__and2b_1
X_06615_ _01522_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07595_ _02266_ _02277_ _02301_ genblk1\[9\].osc.clkdiv_C.cnt\[17\] genblk1\[9\].osc.clkdiv_C.cnt\[16\]
+ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09334_ _03793_ _03748_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06546_ genblk1\[2\].osc.clkdiv_C.cnt\[8\] genblk1\[2\].osc.clkdiv_C.cnt\[7\] _01461_
+ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07619__A2 _01595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06477_ net29 _01405_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__nor2_1
X_09265_ _03853_ genblk1\[0\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08216_ _02900_ _02922_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09196_ net1224 _03712_ _03822_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08147_ genblk1\[3\].osc.clkdiv_C.cnt\[1\] _01496_ _01519_ genblk1\[3\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08078_ genblk1\[5\].osc.clkdiv_C.cnt\[10\] _01667_ _02757_ VGND VGND VPWR VPWR _02785_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_101_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07029_ genblk1\[7\].osc.clkdiv_C.cnt\[16\] _01847_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__or2_1
X_10040_ _04429_ VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold10 modein.delay_octave_up_in\[0\] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 genblk2\[11\].wave_shpr.div.quo\[20\] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 _00558_ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 genblk2\[2\].wave_shpr.div.quo\[21\] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 _00631_ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 genblk2\[6\].wave_shpr.div.acc_next\[0\] VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 genblk2\[5\].wave_shpr.div.quo\[13\] VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__B1 _05417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold87 _00881_ VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 _00307_ VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11991_ _05800_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__clkbuf_1
X_13730_ clknet_leaf_74_clk _01041_ net212 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10942_ net271 _05052_ _05056_ net671 VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13661_ clknet_leaf_47_clk _00974_ net120 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10873_ _04966_ _05015_ _05016_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__a21o_1
X_12612_ clknet_leaf_23_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[15\] net94 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_4
X_13592_ clknet_leaf_72_clk _00907_ net216 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06818__B1 _01675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12543_ clknet_leaf_60_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[0\] net187 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__09480__A1 _04028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10090__A2 _04452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12474_ clknet_leaf_116_clk FSM.next_mode\[0\] net150 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11425_ _05362_ _05399_ _05400_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 _04242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11356_ genblk2\[7\].wave_shpr.div.acc\[22\] _05218_ _05340_ VGND VGND VPWR VPWR
+ _05341_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_842 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10307_ genblk2\[4\].wave_shpr.div.acc\[21\] genblk2\[4\].wave_shpr.div.acc\[20\]
+ _04617_ _04618_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__or4_1
XANTENNA__07717__B _02364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11287_ _05191_ _05176_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__or2b_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ clknet_leaf_113_clk _00353_ net134 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10238_ net375 _04457_ _04454_ _04555_ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__a22o_1
X_10169_ net966 _04486_ _04490_ _04504_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06349__A genblk1\[0\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06400_ _01343_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07380_ genblk1\[11\].osc.clkdiv_C.cnt\[12\] _02130_ VGND VGND VPWR VPWR _02132_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_128_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06331_ genblk1\[0\].osc.clkdiv_C.cnt\[7\] _01281_ genblk1\[0\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09050_ _03708_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__buf_8
XFILLER_0_32_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06262_ _01220_ _01221_ _01223_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__a21oi_4
XANTENNA_clkbuf_leaf_59_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08001_ genblk1\[6\].osc.clkdiv_C.cnt\[15\] _01577_ _01675_ genblk1\[6\].osc.clkdiv_C.cnt\[13\]
+ _02707_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06193_ _01159_ net832 VGND VGND VPWR VPWR PWM.next_counter\[2\] sky130_fd_sc_hd__nor2_1
XFILLER_0_53_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_102_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold502 genblk2\[6\].wave_shpr.div.quo\[4\] VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold513 genblk2\[11\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold524 genblk2\[6\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06812__A _01189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold535 _00234_ VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold546 genblk2\[1\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__buf_1
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold557 genblk2\[0\].wave_shpr.div.i\[2\] VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 genblk2\[0\].wave_shpr.div.acc\[17\] VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09952_ _04352_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__clkbuf_1
Xhold579 genblk2\[7\].wave_shpr.div.acc\[10\] VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08903_ _03574_ _03604_ _03606_ _01157_ net1065 VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ net903 _04282_ _04289_ _04302_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__a22o_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ genblk2\[2\].wave_shpr.div.fin_quo\[0\] _02468_ _03114_ VGND VGND VPWR VPWR
+ _03541_ sky130_fd_sc_hd__a21o_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08765_ _03471_ _03468_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09561__C _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ _02315_ _02421_ _02422_ VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12294__B1 _03733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08696_ _03355_ _03353_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07647_ genblk2\[11\].wave_shpr.div.fin_quo\[3\] _02353_ VGND VGND VPWR VPWR _02354_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_138_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07578_ genblk1\[9\].osc.clkdiv_C.cnt\[7\] _01234_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09317_ _03784_ _03900_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06529_ _01452_ _01453_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[1\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06706__B _01595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09248_ net410 _03845_ _03847_ net522 _03852_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09179_ _03816_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__clkbuf_1
X_11210_ _05244_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__clkbuf_1
X_12190_ genblk2\[11\].wave_shpr.div.acc\[14\] genblk2\[11\].wave_shpr.div.b1\[14\]
+ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__or2b_1
XFILLER_0_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11141_ genblk2\[7\].wave_shpr.div.b1\[10\] genblk2\[7\].wave_shpr.div.acc\[10\]
+ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11072_ net1138 _05119_ _05126_ _05143_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__a22o_1
XANTENNA__09517__A2 _04043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10023_ _04417_ _04418_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__or2_1
XANTENNA__07553__A _01157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11974_ genblk2\[10\].wave_shpr.div.fin_quo\[4\] net1323 _00003_ VGND VGND VPWR VPWR
+ _05792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13713_ clknet_leaf_31_clk _01024_ net99 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10925_ _05047_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06503__A2 _01411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13644_ clknet_leaf_69_clk net321 net211 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_10856_ genblk2\[6\].wave_shpr.div.b1\[9\] genblk2\[6\].wave_shpr.div.acc\[9\] VGND
+ VGND VPWR VPWR _05000_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ clknet_leaf_84_clk net307 net183 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10787_ net982 _04918_ _04922_ _04942_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__a22o_1
XANTENNA__10419__A _04654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12526_ clknet_leaf_66_clk _00078_ net197 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09205__A1 _03704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12457_ clknet_leaf_106_clk _00030_ net155 VGND VGND VPWR VPWR PWM.final_sample_in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11408_ genblk2\[8\].wave_shpr.div.b1\[5\] genblk2\[8\].wave_shpr.div.acc\[5\] VGND
+ VGND VPWR VPWR _05384_ sky130_fd_sc_hd__and2b_1
XANTENNA__07728__A _01342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12388_ _05961_ _05932_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__or2b_1
XANTENNA__07767__A1 genblk1\[0\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07767__B2 genblk1\[0\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11339_ _05214_ _05328_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09508__A2 _04043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11315__A2 _05279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13009_ clknet_leaf_133_clk _00338_ net59 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_06880_ _01729_ _01684_ _01730_ genblk1\[6\].osc.clkdiv_C.cnt\[4\] _01733_ VGND VGND
+ VPWR VPWR _01734_ sky130_fd_sc_hd__a221o_1
X_08550_ _03245_ _03235_ VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07501_ net17 net18 VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__nand2b_4
X_08481_ genblk2\[3\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__inv_2
X_07432_ _02170_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__buf_8
XANTENNA__12028__B1 _05817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07363_ genblk1\[11\].osc.clkdiv_C.cnt\[8\] genblk1\[11\].osc.clkdiv_C.cnt\[7\] _02112_
+ VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09102_ genblk2\[0\].wave_shpr.div.acc\[13\] genblk2\[0\].wave_shpr.div.b1\[13\]
+ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__or2b_1
XFILLER_0_73_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06314_ genblk1\[0\].osc.clkdiv_C.cnt\[2\] genblk1\[0\].osc.clkdiv_C.cnt\[1\] genblk1\[0\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07294_ genblk1\[10\].osc.clkdiv_C.cnt\[16\] _02058_ VGND VGND VPWR VPWR _02060_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_33_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06245_ freq_div.state\[0\] freq_div.state\[2\] freq_div.state\[1\] VGND VGND VPWR
+ VPWR _01207_ sky130_fd_sc_hd__or3b_1
X_09033_ net817 _02202_ _03698_ _03702_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout210_A net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06176_ _01139_ _01133_ _01137_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__and3_1
Xhold310 _00732_ VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 _00384_ VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 genblk2\[7\].wave_shpr.div.quo\[15\] VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold343 genblk2\[3\].wave_shpr.div.quo\[24\] VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold354 genblk2\[5\].wave_shpr.div.quo\[10\] VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 genblk2\[10\].wave_shpr.div.quo\[12\] VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 genblk2\[6\].wave_shpr.div.quo\[15\] VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 genblk2\[2\].wave_shpr.div.acc\[19\] VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 genblk2\[6\].wave_shpr.div.quo\[21\] VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__dlygate4sd3_1
X_09935_ net1034 _04315_ _04322_ _04341_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08707__B1 _02224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12911__RESET_B net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _04250_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__clkbuf_4
Xhold1010 genblk2\[1\].wave_shpr.div.acc\[25\] VGND VGND VPWR VPWR net1228 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10514__B1 _04655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1021 genblk2\[9\].wave_shpr.div.b1\[17\] VGND VGND VPWR VPWR net1239 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09380__B1 _03947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08817_ _03518_ _03521_ _03517_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__a21o_1
Xhold1032 genblk2\[7\].wave_shpr.div.b1\[3\] VGND VGND VPWR VPWR net1250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 sig_norm.quo\[10\] VGND VGND VPWR VPWR net1261 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ _04250_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__clkbuf_4
Xhold1054 genblk2\[1\].wave_shpr.div.b1\[5\] VGND VGND VPWR VPWR net1272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1065 genblk2\[5\].wave_shpr.div.b1\[10\] VGND VGND VPWR VPWR net1283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 genblk2\[9\].wave_shpr.div.b1\[2\] VGND VGND VPWR VPWR net1294 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 genblk2\[0\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR net1305 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ net14 _02744_ _02365_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__nand3_1
Xhold1098 genblk2\[1\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net1316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08486__A2 _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08679_ _02584_ _03385_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__xnor2_2
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _04783_ _04883_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__nor2_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ genblk2\[9\].wave_shpr.div.b1\[5\] genblk2\[9\].wave_shpr.div.acc\[5\] VGND
+ VGND VPWR VPWR _05582_ sky130_fd_sc_hd__and2b_1
XFILLER_0_95_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10641_ _03707_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13360_ clknet_leaf_116_clk _00019_ net139 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10572_ genblk2\[5\].wave_shpr.div.b1\[10\] genblk2\[5\].wave_shpr.div.acc\[10\]
+ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12311_ net467 _03947_ _03944_ net479 _06012_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13291_ clknet_leaf_88_clk _00612_ net177 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12242_ genblk2\[11\].wave_shpr.div.acc\[23\] _05979_ VGND VGND VPWR VPWR _05980_
+ sky130_fd_sc_hd__or2_2
XANTENNA__06452__A genblk1\[1\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12173_ _05815_ _05812_ genblk2\[10\].wave_shpr.div.i\[0\] VGND VGND VPWR VPWR _05916_
+ sky130_fd_sc_hd__mux2_1
X_11124_ genblk2\[7\].wave_shpr.div.b1\[0\] _05182_ _05183_ VGND VGND VPWR VPWR _05184_
+ sky130_fd_sc_hd__a21oi_1
X_11055_ _05011_ _05130_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__xnor2_1
X_10006_ _04367_ _04400_ _04401_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__a21o_1
XANTENNA__11517__B genblk1\[8\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11009__S _05023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08098__B _01576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11957_ _05732_ _05777_ _05778_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_98_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10908_ _05038_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07730__B genblk1\[1\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11888_ _03694_ _05611_ _05717_ _03696_ net1026 VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__a32o_1
XFILLER_0_39_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13627_ clknet_leaf_66_clk _00940_ net197 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10839_ genblk2\[6\].wave_shpr.div.acc\[0\] genblk2\[6\].wave_shpr.div.b1\[0\] VGND
+ VGND VPWR VPWR _04983_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13558_ clknet_leaf_78_clk _00873_ net208 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11784__A2 _02203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12509_ clknet_leaf_84_clk _00071_ net202 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13489_ clknet_leaf_88_clk net470 net177 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08401__A2 _01591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout108 net109 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09673__A _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07981_ _02684_ _02687_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__nand2_1
Xfanout119 net122 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_4
X_09720_ _04160_ _04198_ _04199_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__a21o_1
X_06932_ _01761_ _01775_ _01776_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__10612__A _01738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07905__B _01870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09651_ genblk2\[1\].wave_shpr.div.acc\[22\] _04139_ VGND VGND VPWR VPWR _04140_
+ sky130_fd_sc_hd__xnor2_1
X_06863_ genblk1\[5\].osc.clkdiv_C.cnt\[14\] _01717_ _01720_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__o21a_1
X_08602_ _03188_ _03189_ _02885_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__nor3_1
XFILLER_0_78_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09582_ _04087_ _03979_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__xnor2_1
X_06794_ _01440_ _01171_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__nand2_4
XFILLER_0_54_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07921__A genblk1\[8\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08533_ _03237_ _03239_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13599__RESET_B net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06693__A2_N _01313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08464_ _03163_ _03164_ _03169_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07140__A2 _01334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07415_ _02155_ _02158_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__nor2_1
X_08395_ genblk1\[2\].osc.clkdiv_C.cnt\[10\] _01420_ _03099_ _03100_ _03101_ VGND
+ VGND VPWR VPWR _03102_ sky130_fd_sc_hd__o221a_1
XANTENNA__13181__RESET_B net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09848__A _03702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07346_ genblk1\[11\].osc.clkdiv_C.cnt\[4\] _02101_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07277_ _02027_ _02048_ _02049_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_115_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09016_ _02155_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__buf_4
XANTENNA__09059__S _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06228_ _01186_ _01189_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__nor2_4
XFILLER_0_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06159_ _01114_ _01116_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__nand2_1
Xhold140 genblk2\[11\].wave_shpr.div.quo\[7\] VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 genblk2\[2\].wave_shpr.div.b1\[15\] VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 smpl_rt_clkdiv.clkDiv_inst.cnt\[4\] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 genblk2\[8\].wave_shpr.div.b1\[15\] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 genblk2\[11\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _01058_ VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__dlygate4sd3_1
X_09918_ _04205_ _04157_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__or2b_1
XANTENNA_fanout73_A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09849_ genblk2\[2\].wave_shpr.div.acc\[0\] _00008_ _04275_ net914 _04276_ VGND VGND
+ VPWR VPWR _00317_ sky130_fd_sc_hd__o221a_1
X_12860_ clknet_leaf_129_clk _00191_ net64 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08927__A _01099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _05569_ _05580_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__xor2_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ clknet_leaf_91_clk _00124_ net146 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _02248_ _01144_ _05622_ net1088 VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ genblk2\[9\].wave_shpr.div.acc\[6\] genblk2\[9\].wave_shpr.div.b1\[6\] VGND
+ VGND VPWR VPWR _05565_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13412_ clknet_leaf_120_clk net232 net142 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10624_ genblk2\[6\].wave_shpr.div.b1\[5\] _04838_ _04834_ VGND VGND VPWR VPWR _04839_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11215__B2 _05248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13343_ clknet_leaf_7_clk _00664_ net49 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10555_ genblk2\[5\].wave_shpr.div.b1\[0\] _04781_ _04782_ VGND VGND VPWR VPWR _04783_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12184__A _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13274_ clknet_leaf_118_clk _00017_ net138 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
X_10486_ _04611_ _04729_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__xnor2_1
X_12225_ genblk2\[11\].wave_shpr.div.b1\[11\] genblk2\[11\].wave_shpr.div.acc\[11\]
+ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12156_ genblk2\[10\].wave_shpr.div.acc\[19\] _05900_ genblk2\[10\].wave_shpr.div.acc\[20\]
+ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__o21a_1
X_11107_ genblk2\[7\].wave_shpr.div.acc\[14\] genblk2\[7\].wave_shpr.div.b1\[14\]
+ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__or2b_1
XFILLER_0_75_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12087_ genblk2\[10\].wave_shpr.div.acc\[3\] _05852_ _05787_ VGND VGND VPWR VPWR
+ _05853_ sky130_fd_sc_hd__mux2_1
X_11038_ genblk2\[6\].wave_shpr.div.acc\[11\] _05117_ _05105_ VGND VGND VPWR VPWR
+ _05118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12989_ clknet_leaf_132_clk _00318_ net64 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07122__A2 _01334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07200_ genblk1\[9\].osc.clkdiv_C.cnt\[15\] genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01981_
+ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__and3_1
XANTENNA__11206__A1 _03831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08180_ genblk2\[3\].wave_shpr.div.fin_quo\[4\] _02886_ VGND VGND VPWR VPWR _02887_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11757__A2 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07131_ _01930_ _01250_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07062_ genblk1\[8\].osc.clkdiv_C.cnt\[6\] _01249_ _01879_ _01490_ genblk1\[8\].osc.clkdiv_C.cnt\[7\]
+ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_70_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10717__B1 _04857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08386__A1 _01200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07916__A genblk1\[8\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07964_ _02670_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09703_ genblk2\[2\].wave_shpr.div.b1\[5\] genblk2\[2\].wave_shpr.div.acc\[5\] VGND
+ VGND VPWR VPWR _04183_ sky130_fd_sc_hd__and2b_1
XANTENNA__08138__B2 _02527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06915_ genblk1\[6\].osc.clkdiv_C.cnt\[3\] _01763_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07895_ _02423_ _02601_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__nand2_1
X_09634_ genblk2\[1\].wave_shpr.div.acc\[17\] _04127_ _04010_ VGND VGND VPWR VPWR
+ _04128_ sky130_fd_sc_hd__mux2_1
XANTENNA__10496__A2 _04715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06846_ _01693_ _01708_ _01709_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_78_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09565_ genblk2\[1\].wave_shpr.div.acc\[1\] _04074_ _04011_ VGND VGND VPWR VPWR _04075_
+ sky130_fd_sc_hd__mux2_1
X_06777_ _01650_ _01648_ _01651_ _01600_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08516_ _03220_ _03221_ _03219_ _03222_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__a211oi_2
X_09496_ _04038_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08447_ _03152_ _03153_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__or2b_1
XFILLER_0_135_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07664__A3 _01794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08378_ _03071_ _03074_ _03084_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11748__A2 _05623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07329_ genblk1\[11\].osc.clkdiv_C.cnt\[0\] _02092_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__and2b_1
XFILLER_0_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10340_ _03714_ net1097 _04432_ _03727_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10271_ genblk2\[4\].wave_shpr.div.acc\[0\] VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__inv_2
XANTENNA__10708__B1 _04858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12010_ _03732_ net384 _03733_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__o21a_1
X_12912_ clknet_leaf_34_clk _00243_ net107 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ clknet_leaf_30_clk _00006_ net104 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ clknet_leaf_44_clk _00107_ net120 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11725_ _05615_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__clkbuf_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11656_ _05449_ _05548_ _05550_ _05448_ net726 VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__a32o_1
Xfanout90 net91 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_4
X_10607_ _04828_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11587_ _05392_ _05366_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10947__B1 _05056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13326_ clknet_leaf_25_clk net314 net86 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10538_ genblk2\[5\].wave_shpr.div.acc\[14\] genblk2\[5\].wave_shpr.div.b1\[14\]
+ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__or2b_1
XANTENNA__10411__A2 _04651_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold909 genblk2\[11\].wave_shpr.div.acc\[2\] VGND VGND VPWR VPWR net1127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13257_ clknet_leaf_3_clk _00580_ net46 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09014__C1 _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10469_ _04603_ _04716_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12208_ _05940_ genblk2\[11\].wave_shpr.div.acc\[2\] _05945_ VGND VGND VPWR VPWR
+ _05946_ sky130_fd_sc_hd__a21o_1
X_13188_ clknet_leaf_118_clk _00015_ net139 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
X_12139_ net870 _05876_ _05883_ _05892_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__a22o_1
X_06700_ _01588_ _01589_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__nor2_1
X_07680_ _01181_ genblk1\[10\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR _02387_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06631_ genblk1\[3\].osc.clkdiv_C.cnt\[4\] _01530_ genblk1\[3\].osc.clkdiv_C.cnt\[5\]
+ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09350_ net688 _03903_ _03910_ _03926_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__a22o_1
X_06562_ _01451_ _01474_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__nor2_1
X_08301_ _03005_ _03007_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__or2b_1
X_09281_ net854 _03870_ _03840_ _03873_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06493_ _01197_ _01417_ _01418_ genblk1\[2\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR
+ VPWR _01419_ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08232_ _02225_ _02885_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__and2_2
XFILLER_0_142_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08163_ genblk1\[3\].osc.clkdiv_C.cnt\[13\] _01498_ _02869_ VGND VGND VPWR VPWR _02870_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10938__B1 _05023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07114_ genblk1\[8\].osc.clkdiv_C.cnt\[16\] _01914_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08094_ genblk1\[4\].osc.clkdiv_C.cnt\[14\] _01359_ _01498_ genblk1\[4\].osc.clkdiv_C.cnt\[13\]
+ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07045_ genblk1\[8\].osc.clkdiv_C.cnt\[8\] _01430_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08996_ net1134 _03596_ _01154_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07947_ genblk1\[7\].osc.clkdiv_C.cnt\[6\] _01574_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__or2_1
X_07878_ _02562_ _02584_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__nor2_1
XANTENNA__09072__S _03722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09617_ _03995_ _04114_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06829_ genblk1\[5\].osc.clkdiv_C.cnt\[1\] genblk1\[5\].osc.clkdiv_C.cnt\[0\] genblk1\[5\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__a21oi_1
X_09548_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09479_ _01433_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__inv_2
XANTENNA__08834__A2 _02468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11510_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12490_ clknet_leaf_109_clk _00052_ net158 VGND VGND VPWR VPWR sig_norm.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11441_ _05416_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12496__RESET_B net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11372_ _05248_ _05350_ _05351_ _05251_ net1113 VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__a32o_1
X_13111_ clknet_leaf_115_clk _00436_ net134 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10323_ _04629_ VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07898__A2_N _01309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13042_ clknet_leaf_128_clk _00369_ net67 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10254_ _04449_ genblk2\[4\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR _04566_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06460__A genblk1\[1\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10185_ genblk2\[3\].wave_shpr.div.acc\[11\] _04516_ _04507_ VGND VGND VPWR VPWR
+ _04517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11017__S _05023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12826_ clknet_leaf_62_clk _00159_ net190 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output17_A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ clknet_leaf_52_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[16\] net110 VGND
+ VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_135_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_135_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10093__B1 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11708_ genblk2\[9\].wave_shpr.div.b1\[14\] genblk2\[9\].wave_shpr.div.acc\[14\]
+ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12688_ clknet_leaf_53_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[1\] net112 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11639_ net704 _05507_ _05417_ _05539_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold706 genblk2\[7\].wave_shpr.div.acc\[17\] VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold717 genblk2\[9\].wave_shpr.div.acc\[20\] VGND VGND VPWR VPWR net935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13309_ clknet_leaf_117_clk _00630_ net137 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold728 genblk2\[8\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR net946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold739 genblk2\[10\].wave_shpr.div.acc\[12\] VGND VGND VPWR VPWR net957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08850_ _03552_ _03555_ _03556_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__and3_1
XANTENNA__07564__A2 _01227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07801_ genblk1\[0\].osc.clkdiv_C.cnt\[16\] _01577_ _02501_ _02507_ genblk1\[0\].osc.clkdiv_C.cnt\[17\]
+ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__a221oi_2
X_08781_ _02583_ _03486_ _02582_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_46_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11648__A1 _05441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07732_ genblk1\[1\].osc.clkdiv_C.cnt\[5\] _02433_ _02435_ _02436_ _02438_ VGND VGND
+ VPWR VPWR _02439_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07663_ _01360_ _01224_ _01241_ genblk1\[10\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR
+ VPWR _02370_ sky130_fd_sc_hd__a211o_1
X_09402_ genblk2\[1\].wave_shpr.div.acc\[5\] genblk2\[1\].wave_shpr.div.b1\[5\] VGND
+ VGND VPWR VPWR _03966_ sky130_fd_sc_hd__and2b_1
XFILLER_0_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06614_ genblk1\[3\].osc.clkdiv_C.cnt\[8\] _01483_ _01484_ genblk1\[3\].osc.clkdiv_C.cnt\[0\]
+ _01521_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07594_ _02276_ _02296_ _02300_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__or3_1
X_09333_ net840 _03903_ _03910_ _03913_ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__a22o_1
X_06545_ _01452_ _01463_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_126_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_126_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_62_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09264_ genblk2\[0\].wave_shpr.div.quo\[24\] _03835_ _03838_ net454 _03861_ VGND
+ VGND VPWR VPWR _00147_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06476_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] genblk1\[1\].osc.clkdiv_C.cnt\[14\] _01401_
+ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08215_ _02918_ _02921_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09195_ _03825_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08146_ _02851_ _02852_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08077_ _02755_ _02760_ _02781_ _02783_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07028_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01846_ _01848_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__06280__A _01241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold11 genblk2\[8\].wave_shpr.div.quo\[22\] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 _01054_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 genblk2\[4\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__buf_1
X_08979_ net372 _01157_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__nand2_1
Xhold44 _00313_ VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 genblk2\[0\].wave_shpr.div.i\[4\] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 _00653_ VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 _00557_ VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 genblk2\[9\].wave_shpr.div.quo\[24\] VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ genblk2\[11\].wave_shpr.div.b1\[4\] _04230_ _05433_ VGND VGND VPWR VPWR _05800_
+ sky130_fd_sc_hd__mux2_1
Xhold99 genblk2\[7\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12300__A2 _06009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10941_ net671 _05052_ _05056_ net756 VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13660_ clknet_leaf_47_clk net447 net120 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10872_ genblk2\[6\].wave_shpr.div.b1\[17\] genblk2\[6\].wave_shpr.div.acc\[17\]
+ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12611_ clknet_leaf_23_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[14\] net94 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_117_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_117_clk sky130_fd_sc_hd__clkbuf_16
X_13591_ clknet_leaf_72_clk _00906_ net216 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12542_ clknet_leaf_100_clk net287 net164 VGND VGND VPWR VPWR PWM.pwm_out sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12473_ clknet_leaf_32_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[7\] net99 VGND VGND
+ VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.cnt\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09766__A _01302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11424_ genblk2\[8\].wave_shpr.div.b1\[13\] genblk2\[8\].wave_shpr.div.acc\[13\]
+ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__and2b_1
XFILLER_0_22_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09232__A2 _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11355_ _05219_ _05220_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__and2b_1
XFILLER_0_120_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10306_ genblk2\[4\].wave_shpr.div.acc\[19\] genblk2\[4\].wave_shpr.div.acc\[18\]
+ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11286_ net1030 _05279_ _05283_ _05288_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__a22o_1
XANTENNA__07717__C _02365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13025_ clknet_leaf_113_clk _00352_ net134 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12011__B1_N _03717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10237_ genblk2\[3\].wave_shpr.div.acc\[25\] _04553_ VGND VGND VPWR VPWR _04555_
+ sky130_fd_sc_hd__xnor2_1
X_10168_ genblk2\[3\].wave_shpr.div.acc\[7\] _04503_ _04420_ VGND VGND VPWR VPWR _04504_
+ sky130_fd_sc_hd__mux2_1
X_10099_ _04269_ genblk1\[3\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12809_ clknet_leaf_60_clk _00142_ net187 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_108_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_108_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08564__B _02521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06330_ genblk1\[0\].osc.clkdiv_C.cnt\[8\] genblk1\[0\].osc.clkdiv_C.cnt\[7\] _01281_
+ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__and3_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06365__A _01171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06261_ _01222_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__buf_4
X_08000_ _02706_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06192_ net642 PWM.counter\[0\] net831 VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09223__A2 _03836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold503 _00632_ VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 genblk2\[4\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08431__B1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold525 genblk2\[8\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07908__B _01870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold536 genblk2\[7\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 sig_norm.i\[2\] VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06812__B _01678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09951_ _04250_ _04247_ genblk2\[2\].wave_shpr.div.i\[0\] VGND VGND VPWR VPWR _04352_
+ sky130_fd_sc_hd__mux2_1
Xhold558 genblk2\[11\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold569 genblk2\[4\].wave_shpr.div.acc\[23\] VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08902_ _03583_ _03605_ _03596_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ genblk2\[2\].wave_shpr.div.acc\[7\] _04300_ _04301_ VGND VGND VPWR VPWR _04302_
+ sky130_fd_sc_hd__mux2_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _03538_ _03539_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__nor2_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout190_A net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08764_ _02798_ _03466_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__nand2_1
XANTENNA__07643__B genblk1\[11\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07715_ _02367_ _02420_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__nor2_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12294__A1 _03732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08695_ _03170_ _03171_ _03172_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07646_ genblk2\[11\].wave_shpr.div.fin_quo\[2\] _02352_ VGND VGND VPWR VPWR _02353_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_48_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07577_ genblk1\[9\].osc.clkdiv_C.cnt\[6\] _01512_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09316_ _03785_ _03752_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06528_ genblk1\[2\].osc.clkdiv_C.cnt\[1\] genblk1\[2\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01453_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09247_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06459_ genblk1\[1\].osc.clkdiv_C.cnt\[9\] _01392_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09178_ net1171 _01342_ _03722_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08129_ _02808_ _02815_ _02821_ _02835_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__or4_2
XFILLER_0_114_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11140_ _05172_ _05198_ _05199_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11071_ net622 _05139_ _05142_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__a21o_1
X_10022_ genblk2\[3\].wave_shpr.div.acc\[23\] genblk2\[3\].wave_shpr.div.acc\[25\]
+ genblk2\[3\].wave_shpr.div.acc\[24\] genblk2\[3\].wave_shpr.div.acc\[26\] VGND VGND
+ VPWR VPWR _04418_ sky130_fd_sc_hd__or4_2
XFILLER_0_99_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11973_ _05791_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10924_ genblk2\[7\].wave_shpr.div.b1\[13\] _02374_ _05042_ VGND VGND VPWR VPWR _05047_
+ sky130_fd_sc_hd__mux2_1
X_13712_ clknet_leaf_31_clk _01023_ net100 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07161__B1 genblk1\[9\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10855_ _04975_ _04997_ _04998_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13643_ clknet_leaf_68_clk _00956_ net211 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13574_ clknet_leaf_85_clk _00889_ net183 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10786_ genblk2\[5\].wave_shpr.div.acc\[19\] _04816_ _04941_ VGND VGND VPWR VPWR
+ _04942_ sky130_fd_sc_hd__a21bo_1
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11796__B1 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12525_ clknet_leaf_67_clk _00077_ net194 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08661__B1 _02525_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12456_ clknet_leaf_20_clk net225 net108 VGND VGND VPWR VPWR modein.delay_octave_down_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11407_ _05371_ _05381_ _05382_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12387_ net816 _06039_ _06040_ _06062_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07728__B genblk1\[1\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07767__A2 _01309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11338_ _05215_ _05164_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__or2b_1
XFILLER_0_120_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11269_ _05248_ _05274_ _05275_ _05251_ net1070 VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__a32o_1
X_13008_ clknet_leaf_133_clk _00337_ net59 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07463__B _02153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07500_ _02220_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__buf_4
X_08480_ _03182_ _03186_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07431_ _02152_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__buf_6
XANTENNA__12028__A1 genblk2\[10\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06807__B _01678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07362_ _02118_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09101_ genblk2\[0\].wave_shpr.div.acc\[14\] genblk2\[0\].wave_shpr.div.b1\[14\]
+ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__or2b_1
XFILLER_0_84_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06313_ _01273_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07293_ net1143 _02057_ _02059_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09032_ _03701_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__buf_8
XFILLER_0_115_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06244_ genblk1\[0\].osc.clkdiv_C.cnt\[2\] _01190_ _01204_ _01205_ VGND VGND VPWR
+ VPWR _01206_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold300 genblk2\[10\].wave_shpr.div.quo\[18\] VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__dlygate4sd3_1
X_06175_ _01137_ _01146_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__nand2_1
Xhold311 genblk2\[3\].wave_shpr.div.quo\[22\] VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold322 genblk2\[7\].wave_shpr.div.acc_next\[0\] VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold333 genblk2\[5\].wave_shpr.div.quo\[15\] VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13316__RESET_B net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold344 _00400_ VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 genblk2\[2\].wave_shpr.div.quo\[16\] VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 genblk2\[0\].wave_shpr.div.quo\[12\] VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 genblk2\[6\].wave_shpr.div.quo\[16\] VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold388 _00336_ VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ genblk2\[2\].wave_shpr.div.acc\[20\] _04339_ VGND VGND VPWR VPWR _04341_
+ sky130_fd_sc_hd__xor2_1
Xhold399 genblk2\[8\].wave_shpr.div.quo\[18\] VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__dlygate4sd3_1
X_09865_ net975 _04282_ _04252_ _04288_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__a22o_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1000 genblk2\[0\].wave_shpr.div.fin_quo\[7\] VGND VGND VPWR VPWR net1218 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 genblk1\[5\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR net1229 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 sig_norm.acc\[4\] VGND VGND VPWR VPWR net1240 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09380__A1 _03944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1033 genblk2\[10\].wave_shpr.div.b1\[13\] VGND VGND VPWR VPWR net1251 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ _03521_ _03522_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__nand2_1
Xhold1044 genblk2\[4\].wave_shpr.div.b1\[14\] VGND VGND VPWR VPWR net1262 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ _04249_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__buf_4
Xhold1055 genblk2\[10\].wave_shpr.div.b1\[4\] VGND VGND VPWR VPWR net1273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 genblk2\[10\].wave_shpr.div.b1\[9\] VGND VGND VPWR VPWR net1284 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ _02742_ _03453_ _02745_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__o21ai_2
XANTENNA_clkbuf_leaf_90_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1077 genblk2\[1\].wave_shpr.div.b1\[2\] VGND VGND VPWR VPWR net1295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 _00173_ VGND VGND VPWR VPWR net1306 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1099 genblk2\[9\].wave_shpr.div.quo\[4\] VGND VGND VPWR VPWR net1317 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _02561_ _02562_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__or2_1
XANTENNA__10135__B_N _04455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ _01174_ _01177_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__nand2_4
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10640_ _04847_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10571_ _04771_ _04797_ _04798_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12310_ _05835_ genblk1\[11\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__and2_1
X_13290_ clknet_leaf_88_clk _00611_ net177 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12241_ genblk2\[11\].wave_shpr.div.acc\[22\] genblk2\[11\].wave_shpr.div.acc\[21\]
+ genblk2\[11\].wave_shpr.div.acc\[20\] _05978_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12172_ net1081 _05818_ _05816_ _05915_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__a22o_1
XANTENNA__06957__B1 _01732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11123_ genblk2\[7\].wave_shpr.div.b1\[1\] genblk2\[7\].wave_shpr.div.acc\[1\] VGND
+ VGND VPWR VPWR _05183_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11054_ _05012_ _04968_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__or2b_1
X_10005_ genblk2\[3\].wave_shpr.div.b1\[11\] genblk2\[3\].wave_shpr.div.acc\[11\]
+ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__and2b_1
XANTENNA_clkbuf_leaf_58_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_101_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11956_ _03832_ genblk2\[10\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR _05778_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07134__B1 _01923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10907_ net1293 _05037_ _04848_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11887_ _05715_ _05716_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13626_ clknet_leaf_67_clk _00939_ net195 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10838_ genblk2\[6\].wave_shpr.div.acc\[1\] genblk2\[6\].wave_shpr.div.b1\[1\] VGND
+ VGND VPWR VPWR _04982_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10769_ _04810_ _04765_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__or2b_1
X_13557_ clknet_leaf_97_clk net268 net169 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12508_ clknet_leaf_103_clk _00070_ net156 VGND VGND VPWR VPWR PWM.final_in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13488_ clknet_leaf_88_clk net330 net177 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10992__B2 _05052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12439_ genblk2\[11\].wave_shpr.div.acc\[24\] _03947_ _03944_ _06100_ VGND VGND VPWR
+ VPWR _01083_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07980_ _02685_ _02686_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__and2_1
Xfanout109 net127 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_2
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06931_ genblk1\[6\].osc.clkdiv_C.cnt\[9\] _01773_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__nor2_1
X_09650_ genblk2\[1\].wave_shpr.div.acc\[21\] _04007_ _04129_ VGND VGND VPWR VPWR
+ _04139_ sky130_fd_sc_hd__or3_1
X_06862_ net27 _01719_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__nor2_1
X_08601_ _03251_ _03252_ _03255_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__and3b_1
X_09581_ _03980_ _03966_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__nor2_1
X_06793_ genblk1\[5\].osc.clkdiv_C.cnt\[3\] _01592_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08532_ _02416_ _03238_ net2 _02364_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__o211a_1
XANTENNA__07921__B _01430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08463_ _03163_ _03164_ _03169_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__nand3_2
XFILLER_0_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07414_ genblk2\[1\].wave_shpr.div.busy _02157_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08394_ genblk1\[2\].osc.clkdiv_C.cnt\[11\] _01411_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07345_ genblk1\[11\].osc.clkdiv_C.cnt\[4\] _02101_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__nand2_1
XANTENNA__11224__A2 _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_16
X_07276_ genblk1\[10\].osc.clkdiv_C.cnt\[9\] _02046_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09015_ genblk2\[9\].wave_shpr.div.i\[0\] _02202_ genblk2\[9\].wave_shpr.div.i\[1\]
+ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__a21oi_1
X_06227_ _01174_ _01187_ _01188_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_131_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12185__B1 _03855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold130 genblk2\[9\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 smpl_rt_clkdiv.clkDiv_inst.cnt\[2\] VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__dlygate4sd3_1
X_06158_ net12 VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold152 genblk2\[7\].wave_shpr.div.quo\[11\] VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 genblk2\[7\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 genblk2\[5\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _01036_ VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 genblk2\[1\].wave_shpr.div.quo\[4\] VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09917_ net845 _04315_ _04322_ _04328_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_97_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_16
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ _03702_ _01416_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout66_A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09779_ _04239_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__clkbuf_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11810_ net886 _05652_ _05653_ _05659_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__a22o_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ clknet_leaf_57_clk _00123_ net182 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _02248_ _01145_ _05622_ net1073 VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__a22o_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ genblk2\[9\].wave_shpr.div.acc\[7\] genblk2\[9\].wave_shpr.div.b1\[7\] VGND
+ VGND VPWR VPWR _05564_ sky130_fd_sc_hd__or2b_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13411_ clknet_leaf_91_clk _00730_ net144 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10623_ _01747_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11215__A2 _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06890__A2 _01519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_16
X_13342_ clknet_leaf_7_clk _00663_ net49 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10554_ genblk2\[5\].wave_shpr.div.b1\[1\] genblk2\[5\].wave_shpr.div.acc\[1\] VGND
+ VGND VPWR VPWR _04782_ sky130_fd_sc_hd__xor2_1
XFILLER_0_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13273_ clknet_leaf_12_clk _00016_ net51 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
X_10485_ _04612_ _04567_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__or2b_1
XFILLER_0_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12224_ _05932_ _05960_ _05961_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12155_ _05783_ _05899_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__nor2_1
XANTENNA__10713__A _02183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11106_ genblk2\[7\].wave_shpr.div.acc\[15\] genblk2\[7\].wave_shpr.div.b1\[15\]
+ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__or2b_1
X_12086_ _05751_ _05851_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_88_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_16
X_11037_ _05003_ _05116_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12988_ clknet_leaf_124_clk net915 net71 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_148_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11939_ _05741_ _05759_ _05760_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10662__B1 _04857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10594__S _00015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13609_ clknet_leaf_58_clk _00922_ net194 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_12_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07130_ genblk1\[9\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07061_ genblk1\[8\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07916__B _01487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07963_ _01200_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01361_ _02668_ _02669_ VGND
+ VGND VPWR VPWR _02670_ sky130_fd_sc_hd__o311a_1
Xclkbuf_leaf_79_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08138__A2 _02309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09702_ _04169_ _04180_ _04181_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__a21o_1
X_06914_ genblk1\[6\].osc.clkdiv_C.cnt\[3\] _01763_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__and2_1
X_07894_ _02520_ net24 _02599_ _02600_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__o31a_1
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07932__A genblk2\[8\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09633_ _04003_ _04126_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__xnor2_1
X_06845_ genblk1\[5\].osc.clkdiv_C.cnt\[7\] _01705_ genblk1\[5\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__a21oi_1
X_09564_ _03970_ _03971_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__xor2_1
X_06776_ genblk1\[4\].osc.clkdiv_C.cnt\[15\] _01647_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__or2_1
X_08515_ _03127_ _03218_ _03204_ _03217_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09495_ net1271 net35 _04024_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08446_ _03024_ _03028_ VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__xor2_2
XFILLER_0_93_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08763__A net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08377_ _03073_ _03072_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12285__A _03702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07328_ _02091_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__buf_2
XANTENNA__09810__A2 _04253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07259_ genblk1\[10\].osc.clkdiv_C.cnt\[4\] _02034_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__or2_1
XANTENNA__07821__B2 _02527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10270_ genblk2\[4\].wave_shpr.div.acc\[2\] genblk2\[4\].wave_shpr.div.b1\[2\] VGND
+ VGND VPWR VPWR _04582_ sky130_fd_sc_hd__or2b_1
XANTENNA__10708__A1 _04855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12911_ clknet_leaf_34_clk _00242_ net107 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ clknet_leaf_65_clk _00175_ net197 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ clknet_leaf_47_clk _00106_ net119 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10644__B1 _04647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ genblk2\[9\].wave_shpr.div.fin_quo\[1\] net1328 _00023_ VGND VGND VPWR VPWR
+ _05615_ sky130_fd_sc_hd__mux2_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11655_ _05549_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout80 net83 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout91 net127 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_4
X_10606_ genblk2\[5\].wave_shpr.div.fin_quo\[6\] net1315 _00015_ VGND VGND VPWR VPWR
+ _04828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11586_ net922 _05447_ _05484_ _05500_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__a22o_1
XANTENNA__09262__B1 _03838_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09801__A2 _04248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10537_ genblk2\[5\].wave_shpr.div.acc\[15\] genblk2\[5\].wave_shpr.div.b1\[15\]
+ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__or2b_1
X_13325_ clknet_leaf_26_clk _00646_ net87 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10468_ _04604_ _04571_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__or2b_1
X_13256_ clknet_leaf_3_clk net773 net51 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12207_ _05940_ genblk2\[11\].wave_shpr.div.acc\[2\] _05944_ VGND VGND VPWR VPWR
+ _05945_ sky130_fd_sc_hd__o21a_1
XANTENNA__12134__S _05865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13187_ clknet_leaf_11_clk _00014_ net56 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
X_10399_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__and2_1
XANTENNA__11372__A1 _05248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07576__B1 _01234_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12138_ genblk2\[10\].wave_shpr.div.acc\[15\] _05891_ _05865_ VGND VGND VPWR VPWR
+ _05892_ sky130_fd_sc_hd__mux2_1
X_12069_ net247 _05812_ _05815_ net446 _05839_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_1_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11274__A _05245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06630_ genblk1\[3\].osc.clkdiv_C.cnt\[5\] genblk1\[3\].osc.clkdiv_C.cnt\[4\] _01530_
+ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06368__A _01309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06561_ genblk1\[2\].osc.clkdiv_C.cnt\[13\] genblk1\[2\].osc.clkdiv_C.cnt\[12\] _01470_
+ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08300_ _02927_ _03006_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__and2_1
X_09280_ genblk2\[0\].wave_shpr.div.acc\[2\] _03872_ _03804_ VGND VGND VPWR VPWR _03873_
+ sky130_fd_sc_hd__mux2_1
X_06492_ _01229_ _01182_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__nand2_2
XANTENNA__06303__A1 genblk1\[0\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08231_ _02937_ _02936_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06815__B _01355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08162_ _02866_ _02867_ _02868_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10938__A1 net792 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10938__B2 _05055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07113_ genblk1\[8\].osc.clkdiv_C.cnt\[15\] _01912_ _01915_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08093_ genblk1\[4\].osc.clkdiv_C.cnt\[14\] _01360_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09618__S _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07044_ _01854_ _01856_ _01857_ _01861_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__or4_1
XFILLER_0_100_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07567__B1 _01349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08995_ net428 _00024_ _03676_ _03677_ VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07946_ genblk1\[7\].osc.clkdiv_C.cnt\[6\] _01574_ _01802_ genblk1\[7\].osc.clkdiv_C.cnt\[5\]
+ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__a22o_1
X_07877_ _02571_ _02582_ _02583_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__a21o_1
XANTENNA__08531__A2 _02525_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09616_ _03996_ _03958_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__or2b_1
X_06828_ genblk1\[5\].osc.clkdiv_C.cnt\[2\] genblk1\[5\].osc.clkdiv_C.cnt\[1\] genblk1\[5\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__and3_1
XANTENNA__06278__A _01238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06759_ _01637_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__inv_2
X_09547_ net257 _04052_ _04053_ net417 _04064_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__a221o_1
X_09478_ _04027_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08429_ _03131_ _03132_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__xor2_1
XFILLER_0_81_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11440_ _05415_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__buf_2
XFILLER_0_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08598__A2 _02592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11371_ genblk2\[7\].wave_shpr.div.i\[1\] genblk2\[7\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _05351_ sky130_fd_sc_hd__nand2_1
X_10322_ genblk2\[4\].wave_shpr.div.fin_quo\[5\] genblk2\[4\].wave_shpr.div.quo\[4\]
+ _00013_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__mux2_1
X_13110_ clknet_leaf_114_clk _00435_ net133 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13041_ clknet_leaf_126_clk _00368_ net66 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10253_ genblk2\[4\].wave_shpr.div.acc\[17\] genblk2\[4\].wave_shpr.div.b1\[17\]
+ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__or2b_1
X_10184_ _04400_ _04515_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12303__B1 _06010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07572__A genblk1\[9\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12825_ clknet_leaf_62_clk _00158_ net190 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ clknet_leaf_50_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[15\] net110 VGND
+ VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11290__B1 _05283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11541__B genblk1\[8\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11707_ _05558_ _05597_ _05598_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12687_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[0\] net174 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11638_ _05412_ _05538_ _05471_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11569_ net898 _05447_ _05484_ _05487_ VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold707 genblk2\[5\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13308_ clknet_leaf_117_clk _00629_ net137 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold718 _00911_ VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 genblk2\[8\].wave_shpr.div.acc\[15\] VGND VGND VPWR VPWR net947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13239_ clknet_leaf_10_clk _00562_ net57 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06370__B _01313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09962__A _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07800_ _02475_ _02476_ _02478_ _02504_ _02506_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__o221a_1
X_08780_ _02583_ _03486_ _02582_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__or3b_1
X_07731_ genblk1\[1\].osc.clkdiv_C.cnt\[6\] _01360_ net37 _02437_ VGND VGND VPWR VPWR
+ _02438_ sky130_fd_sc_hd__a31o_1
XANTENNA__07482__A _02147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07662_ genblk1\[10\].osc.clkdiv_C.cnt\[5\] _01182_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__or2_1
X_06613_ _01485_ _01256_ _01511_ _01518_ _01520_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__o2111a_1
X_09401_ genblk2\[1\].wave_shpr.div.b1\[6\] VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07593_ _02270_ _02297_ _02299_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__or3b_1
X_09332_ genblk2\[0\].wave_shpr.div.acc\[14\] _03912_ _03889_ VGND VGND VPWR VPWR
+ _03913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06544_ genblk1\[2\].osc.clkdiv_C.cnt\[7\] _01461_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12073__A2 _05787_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09263_ _03853_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06475_ genblk1\[1\].osc.clkdiv_C.cnt\[14\] _01401_ _01404_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__o21a_1
X_08214_ _02747_ _02919_ _02920_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__nand3_1
XFILLER_0_8_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09194_ net1284 _01991_ _03822_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__mux2_1
XANTENNA__09226__B1 _03840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08145_ _01201_ genblk1\[3\].osc.clkdiv_C.cnt\[15\] genblk1\[3\].osc.clkdiv_C.cnt\[14\]
+ _01362_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_16_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07657__A net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08076_ genblk1\[5\].osc.clkdiv_C.cnt\[8\] _01678_ _02782_ VGND VGND VPWR VPWR _02783_
+ sky130_fd_sc_hd__a21bo_1
X_07027_ _01822_ _01847_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10083__A _02170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10139__A2 _04420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold12 _00818_ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 genblk2\[6\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _03661_ _03663_ _02248_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__mux2_1
Xhold34 _00468_ VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 genblk2\[8\].wave_shpr.div.quo\[17\] VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 genblk2\[8\].wave_shpr.div.acc_next\[0\] VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__buf_1
Xhold67 genblk2\[1\].wave_shpr.div.i\[4\] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _02221_ net30 VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__nor2_2
Xhold78 genblk2\[3\].wave_shpr.div.quo\[19\] VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 _00890_ VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10940_ net756 _05052_ _05056_ net792 VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10871_ _04851_ genblk2\[6\].wave_shpr.div.acc\[16\] _05014_ VGND VGND VPWR VPWR
+ _05015_ sky130_fd_sc_hd__a21o_1
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12610_ clknet_leaf_22_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[13\] net93 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13590_ clknet_leaf_73_clk _00905_ net215 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10075__A1 _01365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12541_ clknet_leaf_64_clk _00093_ net189 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12472_ clknet_leaf_32_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[6\] net99 VGND VGND
+ VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.cnt\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09768__A1 _01262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11423_ _05363_ _05397_ _05398_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09766__B _03727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11354_ net706 _05311_ _05315_ _05339_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__a22o_1
XANTENNA__07243__A2 _01235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10305_ _04565_ _04615_ _04616_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__a21o_1
X_11285_ net877 _05287_ _05222_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10236_ net1021 _04457_ _04454_ _04554_ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__a22o_1
X_13024_ clknet_leaf_114_clk _00351_ net132 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09782__A _03702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10167_ _04392_ _04502_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07951__B1 _01732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10098_ net538 _04457_ _04454_ genblk2\[3\].wave_shpr.div.quo\[8\] _04458_ VGND VGND
+ VPWR VPWR _00384_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12808_ clknet_leaf_60_clk net411 net187 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10066__A1 _04229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09022__A _03693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11263__B1 _05249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12739_ clknet_leaf_48_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[16\] net114 VGND
+ VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_155_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06260_ freq_div.state\[0\] freq_div.state\[1\] freq_div.state\[2\] VGND VGND VPWR
+ VPWR _01222_ sky130_fd_sc_hd__and3b_1
XFILLER_0_115_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06690__B1 _01578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06191_ PWM.counter\[1\] PWM.counter\[0\] PWM.counter\[2\] VGND VGND VPWR VPWR _01159_
+ sky130_fd_sc_hd__and3_1
Xhold504 genblk2\[8\].wave_shpr.div.b1\[14\] VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 _00463_ VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold526 _00796_ VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold537 genblk2\[1\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 _00028_ VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 genblk2\[4\].wave_shpr.div.acc\[25\] VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ net962 _04253_ _04251_ _04351_ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08901_ _03582_ _03577_ _03581_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_4_9_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _04213_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _03531_ _03537_ _03536_ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__a21oi_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07942__B1 _01925_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ net9 _02744_ _03469_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout183_A net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07714_ _02367_ _02420_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__xor2_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _03397_ _03400_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07940__A net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07645_ genblk2\[11\].wave_shpr.div.fin_quo\[0\] genblk2\[11\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07576_ genblk1\[9\].osc.clkdiv_C.cnt\[6\] _01512_ _01234_ genblk1\[9\].osc.clkdiv_C.cnt\[7\]
+ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10057__A1 _01329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09315_ net1004 _03870_ _03877_ _03899_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__a22o_1
X_06527_ net1051 _01452_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06458_ _01373_ _01392_ _01393_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_118_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09246_ net522 _03845_ _03847_ net543 _03851_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06681__B1 _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09177_ _03815_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__clkbuf_1
X_06389_ _01179_ _01332_ _01225_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__or3_1
X_08128_ _02826_ _02828_ _02832_ _02833_ _02834_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__o311a_1
XFILLER_0_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08059_ genblk1\[5\].osc.clkdiv_C.cnt\[5\] _01238_ net36 genblk1\[5\].osc.clkdiv_C.cnt\[4\]
+ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout96_A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11070_ _05019_ net21 VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10021_ genblk2\[3\].wave_shpr.div.acc\[22\] _04416_ VGND VGND VPWR VPWR _04417_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_101_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11972_ genblk2\[10\].wave_shpr.div.fin_quo\[3\] genblk2\[10\].wave_shpr.div.quo\[2\]
+ _00003_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13711_ clknet_leaf_31_clk _01022_ net100 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10923_ _05046_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07161__A1 genblk1\[9\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13642_ clknet_leaf_95_clk _00955_ net161 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_10854_ genblk2\[6\].wave_shpr.div.b1\[8\] genblk2\[6\].wave_shpr.div.acc\[8\] VGND
+ VGND VPWR VPWR _04998_ sky130_fd_sc_hd__and2b_1
XANTENNA__10048__A1 _01223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13573_ clknet_leaf_86_clk net227 net183 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10785_ genblk2\[5\].wave_shpr.div.acc\[19\] _04938_ VGND VGND VPWR VPWR _04941_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_27_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06185__B _01097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11796__A1 _03694_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09777__A _03701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12524_ clknet_leaf_59_clk _00076_ net193 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06672__B1 _01498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12480__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12455_ clknet_leaf_33_clk net4 net101 VGND VGND VPWR VPWR modein.delay_octave_down_in\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_151_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11406_ genblk2\[8\].wave_shpr.div.b1\[4\] genblk2\[8\].wave_shpr.div.acc\[4\] VGND
+ VGND VPWR VPWR _05382_ sky130_fd_sc_hd__and2b_1
XFILLER_0_34_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12386_ genblk2\[11\].wave_shpr.div.acc\[9\] _06061_ _06055_ VGND VGND VPWR VPWR
+ _06062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11337_ net924 _05311_ _05315_ _05327_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11268_ genblk2\[7\].wave_shpr.div.b1\[0\] _05222_ genblk2\[7\].wave_shpr.div.acc\[0\]
+ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13007_ clknet_leaf_138_clk net606 net40 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11547__A _05444_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12142__S _05865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10219_ net1055 _04518_ _04522_ _04542_ VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__a22o_1
X_11199_ _05240_ VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09017__A _03689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07760__A _02362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11484__B1 _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07430_ _02169_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__inv_2
XANTENNA__12028__A2 _05813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07361_ _02091_ _02116_ _02117_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09100_ genblk2\[0\].wave_shpr.div.acc\[15\] genblk2\[0\].wave_shpr.div.b1\[15\]
+ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__or2b_1
X_06312_ _01270_ _01271_ _01272_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07292_ _02026_ _02058_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09031_ _02155_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__buf_8
XFILLER_0_14_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06243_ genblk1\[0\].osc.clkdiv_C.cnt\[17\] _01197_ _01198_ VGND VGND VPWR VPWR _01205_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06174_ _01134_ _01136_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08404__A1 _01201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold301 genblk2\[1\].wave_shpr.div.quo\[13\] VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 genblk2\[9\].wave_shpr.div.quo\[17\] VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 genblk2\[9\].wave_shpr.div.quo\[13\] VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold334 genblk2\[1\].wave_shpr.div.quo\[17\] VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold345 genblk2\[7\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 genblk2\[2\].wave_shpr.div.quo\[9\] VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 genblk2\[7\].wave_shpr.div.quo\[17\] VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09626__S _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold378 genblk2\[4\].wave_shpr.div.quo\[14\] VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ net648 _04315_ _04322_ _04340_ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__a22o_1
Xhold389 genblk2\[3\].wave_shpr.div.quo\[21\] VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08707__A2 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ genblk2\[2\].wave_shpr.div.acc\[3\] _04287_ _04214_ VGND VGND VPWR VPWR _04288_
+ sky130_fd_sc_hd__mux2_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10514__A2 _04657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1001 _03812_ VGND VGND VPWR VPWR net1219 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07915__B1 _01487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1012 genblk2\[9\].wave_shpr.div.b1\[3\] VGND VGND VPWR VPWR net1230 sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ _03516_ _03520_ _03445_ _03450_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__a211o_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 genblk2\[10\].wave_shpr.div.acc\[6\] VGND VGND VPWR VPWR net1241 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _02152_ genblk2\[2\].wave_shpr.div.busy _02162_ VGND VGND VPWR VPWR _04249_
+ sky130_fd_sc_hd__and3_1
Xhold1034 genblk1\[7\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR net1252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 genblk2\[4\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net1263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1056 genblk2\[1\].wave_shpr.div.b1\[7\] VGND VGND VPWR VPWR net1274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 genblk2\[3\].wave_shpr.div.b1\[12\] VGND VGND VPWR VPWR net1285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08746_ _02217_ _02553_ genblk2\[6\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR
+ _03453_ sky130_fd_sc_hd__and3_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1078 genblk1\[9\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR net1296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 PWM.counter\[4\] VGND VGND VPWR VPWR net1307 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _03298_ _03333_ _03381_ _03382_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__a211oi_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07628_ genblk1\[11\].osc.clkdiv_C.cnt\[12\] _01256_ _02333_ _02334_ VGND VGND VPWR
+ VPWR _02335_ sky130_fd_sc_hd__a211o_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07559_ _01200_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01361_ genblk1\[9\].osc.clkdiv_C.cnt\[15\]
+ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__a211o_1
X_10570_ genblk2\[5\].wave_shpr.div.b1\[9\] genblk2\[5\].wave_shpr.div.acc\[9\] VGND
+ VGND VPWR VPWR _04798_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09229_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12240_ genblk2\[11\].wave_shpr.div.acc\[19\] _05977_ VGND VGND VPWR VPWR _05978_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_121_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06406__B1 genblk1\[1\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12171_ genblk2\[10\].wave_shpr.div.acc\[25\] _05785_ _05914_ VGND VGND VPWR VPWR
+ _05915_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07845__A net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11122_ genblk2\[7\].wave_shpr.div.acc\[0\] VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__inv_2
XANTENNA__10047__A2_N _04432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold890 genblk2\[4\].wave_shpr.div.i\[1\] VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__dlygate4sd3_1
X_11053_ net818 _05119_ _05126_ _05129_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__a22o_1
XANTENNA_hold944_A genblk1\[8\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10505__A2 _04715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10004_ _04368_ _04398_ _04399_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11955_ _05733_ _05775_ _05776_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08331__B1 _02526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10906_ _01805_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__inv_2
X_11886_ genblk2\[9\].wave_shpr.div.acc\[23\] _05610_ VGND VGND VPWR VPWR _05716_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11218__B1 _05250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13625_ clknet_leaf_68_clk _00938_ net194 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10837_ genblk2\[6\].wave_shpr.div.b1\[2\] VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__inv_2
XANTENNA__12661__RESET_B net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13556_ clknet_leaf_101_clk _00871_ net164 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08634__A1 genblk2\[8\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10768_ net835 _04918_ _04922_ _04928_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12507_ clknet_leaf_103_clk _00069_ net156 VGND VGND VPWR VPWR PWM.final_in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13487_ clknet_leaf_89_clk _00804_ net177 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10699_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12438_ genblk2\[11\].wave_shpr.div.acc\[23\] _05979_ _06099_ VGND VGND VPWR VPWR
+ _06100_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12369_ genblk2\[11\].wave_shpr.div.acc\[5\] _06048_ _05982_ VGND VGND VPWR VPWR
+ _06049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06930_ genblk1\[6\].osc.clkdiv_C.cnt\[9\] _01773_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__and2_1
X_06861_ genblk1\[5\].osc.clkdiv_C.cnt\[14\] _01717_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__and2_1
X_08600_ _03304_ _03306_ _03302_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__a21o_1
X_09580_ net825 _04076_ _04080_ _04086_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__a22o_1
X_06792_ _01659_ _01661_ _01662_ _01663_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__or4_1
X_08531_ genblk2\[10\].wave_shpr.div.fin_quo\[0\] _02525_ _02307_ genblk2\[10\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08462_ _02742_ _03167_ _03168_ _02745_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__o31a_1
XANTENNA__07676__A2 _01190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07413_ genblk2\[1\].wave_shpr.div.i\[1\] _02156_ genblk2\[1\].wave_shpr.div.i\[4\]
+ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__or3b_1
XFILLER_0_148_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08393_ genblk1\[2\].osc.clkdiv_C.cnt\[10\] _01420_ _01431_ genblk1\[2\].osc.clkdiv_C.cnt\[9\]
+ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout146_A net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07344_ _02104_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09210__A _02170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07275_ genblk1\[10\].osc.clkdiv_C.cnt\[9\] _02046_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06226_ _01178_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__buf_4
X_09014_ genblk2\[9\].wave_shpr.div.busy genblk2\[9\].wave_shpr.div.i\[0\] _03686_
+ _03687_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold120 smpl_rt_clkdiv.clkDiv_inst.cnt\[0\] VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__dlymetal6s2s_1
X_06157_ _01113_ _01117_ _01128_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__a21oi_1
Xhold131 genblk2\[9\].wave_shpr.div.quo\[16\] VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 _01090_ VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold153 _00723_ VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _00763_ VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 genblk2\[2\].wave_shpr.div.quo\[17\] VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 genblk2\[8\].wave_shpr.div.quo\[7\] VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _00212_ VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__dlygate4sd3_1
X_09916_ genblk2\[2\].wave_shpr.div.acc\[15\] _04327_ _04301_ VGND VGND VPWR VPWR
+ _04328_ sky130_fd_sc_hd__mux2_1
X_09847_ _04250_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__inv_2
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ net1297 _01487_ _04238_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout59_A net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11448__A0 genblk2\[8\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _03434_ _03435_ genblk2\[2\].wave_shpr.div.fin_quo\[5\] _02468_ VGND VGND
+ VPWR VPWR _03436_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08313__B1 _02525_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11999__A1 _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _01099_ _01149_ _05622_ net497 VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_68_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ genblk2\[9\].wave_shpr.div.acc\[8\] genblk2\[9\].wave_shpr.div.b1\[8\] VGND
+ VGND VPWR VPWR _05563_ sky130_fd_sc_hd__or2b_1
XFILLER_0_95_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13410_ clknet_leaf_90_clk _00729_ net144 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10622_ _04837_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13341_ clknet_leaf_7_clk _00662_ net49 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10553_ genblk2\[5\].wave_shpr.div.acc\[0\] VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13272_ clknet_leaf_136_clk _00595_ net41 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10484_ net784 _04715_ _04722_ _04728_ VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12223_ genblk2\[11\].wave_shpr.div.b1\[10\] genblk2\[11\].wave_shpr.div.acc\[10\]
+ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09041__A1 _03706_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12154_ net705 _05876_ _05883_ _05903_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__a22o_1
X_11105_ _05049_ genblk2\[7\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR _05165_
+ sky130_fd_sc_hd__nor2_1
X_12085_ _05752_ _05744_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__or2b_1
X_11036_ _05004_ _04972_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__or2b_1
XANTENNA__08552__B1 genblk2\[6\].wave_shpr.div.fin_quo\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12987_ clknet_leaf_125_clk net260 net69 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11938_ genblk2\[10\].wave_shpr.div.b1\[7\] genblk2\[10\].wave_shpr.div.acc\[7\]
+ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11869_ _05608_ _05646_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13608_ clknet_leaf_58_clk _00921_ net194 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09804__B1 _04252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13539_ clknet_leaf_100_clk _00854_ net165 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_42_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06373__B _01240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07060_ genblk1\[8\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07485__A _02209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07043__B1 _01858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09176__S _03722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07962_ genblk1\[7\].osc.clkdiv_C.cnt\[14\] _01361_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__nand2_1
X_09701_ genblk2\[2\].wave_shpr.div.b1\[4\] genblk2\[2\].wave_shpr.div.acc\[4\] VGND
+ VGND VPWR VPWR _04181_ sky130_fd_sc_hd__and2b_1
X_06913_ _01761_ _01763_ _01764_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07893_ _02529_ _02594_ _02518_ _02598_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__a22o_1
X_09632_ _04004_ _03954_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__or2b_1
XANTENNA__07932__B genblk2\[8\].wave_shpr.div.fin_quo\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06844_ genblk1\[5\].osc.clkdiv_C.cnt\[8\] genblk1\[5\].osc.clkdiv_C.cnt\[7\] _01705_
+ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09563_ _04045_ _04072_ _04073_ _04048_ genblk2\[1\].wave_shpr.div.acc\[1\] VGND
+ VGND VPWR VPWR _00234_ sky130_fd_sc_hd__a32o_1
X_06775_ genblk1\[4\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__inv_2
X_08514_ _03208_ _03215_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__or2b_1
X_09494_ _04037_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10102__B1 _04454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08445_ _03140_ _03150_ _03151_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_77_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08376_ _03081_ _03082_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06609__B1 _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07327_ _02069_ _02072_ _02073_ _02090_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__or4_4
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07258_ genblk1\[10\].osc.clkdiv_C.cnt\[4\] _02034_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07821__A2 _02521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06209_ _01170_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__buf_4
X_07189_ genblk1\[9\].osc.clkdiv_C.cnt\[11\] genblk1\[9\].osc.clkdiv_C.cnt\[10\] _01974_
+ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07585__A1 genblk1\[9\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08534__B1 _02308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12910_ clknet_leaf_33_clk _00241_ net100 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12841_ clknet_leaf_64_clk _00174_ net196 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ clknet_leaf_47_clk _00105_ net121 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _05614_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10644__A1 _03704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11654_ genblk2\[8\].wave_shpr.div.i\[1\] genblk2\[8\].wave_shpr.div.i\[0\] genblk2\[8\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout70 net75 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout81 net83 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10605_ _04827_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__clkbuf_1
Xfanout92 net94 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11585_ genblk2\[8\].wave_shpr.div.acc\[8\] _05499_ _05493_ VGND VGND VPWR VPWR _05500_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10947__A2 _05052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13324_ clknet_leaf_26_clk _00645_ net87 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10536_ _04649_ genblk2\[5\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR _04764_
+ sky130_fd_sc_hd__nor2_1
X_13255_ clknet_leaf_2_clk _00578_ net51 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10467_ _04651_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__clkbuf_4
X_12206_ _05941_ _05942_ _05943_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13186_ clknet_leaf_112_clk _00511_ net129 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10398_ net680 _04661_ _04663_ genblk2\[4\].wave_shpr.div.quo\[15\] _04667_ VGND
+ VGND VPWR VPWR _00475_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12137_ _05775_ _05890_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12068_ _05835_ genblk1\[10\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR _05839_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11555__A _05417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11019_ _04996_ _04976_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__or2b_1
XFILLER_0_149_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06368__B _01221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06560_ net1256 _01470_ _01473_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06491_ genblk1\[2\].osc.clkdiv_C.cnt\[16\] _01363_ _01416_ VGND VGND VPWR VPWR _01417_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06303__A2 _01256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08230_ _02798_ _02931_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08161_ genblk1\[3\].osc.clkdiv_C.cnt\[13\] _01498_ VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10938__A2 _05052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07112_ _01886_ _01914_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__nor2_1
X_08092_ _02791_ _02796_ _02798_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_70_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07043_ genblk1\[8\].osc.clkdiv_C.cnt\[5\] _01487_ _01858_ genblk1\[8\].osc.clkdiv_C.cnt\[6\]
+ _01860_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout109_A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11899__B1 _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07567__A1 genblk1\[9\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08994_ sig_norm.quo\[10\] _01099_ _01157_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__a21o_1
X_07945_ genblk1\[7\].osc.clkdiv_C.cnt\[5\] _01802_ _01805_ genblk1\[7\].osc.clkdiv_C.cnt\[4\]
+ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__o22a_1
XANTENNA__07662__B _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07876_ _02517_ _02570_ _02566_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__and3_1
X_09615_ _04046_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__buf_2
X_06827_ _01697_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[1\] sky130_fd_sc_hd__clkbuf_1
X_09546_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__and2_1
X_06758_ genblk1\[4\].osc.clkdiv_C.cnt\[11\] genblk1\[4\].osc.clkdiv_C.cnt\[10\] _01631_
+ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__and3_1
XANTENNA__10626__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09477_ genblk2\[2\].wave_shpr.div.b1\[6\] _01437_ _04024_ VGND VGND VPWR VPWR _04027_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06689_ genblk1\[4\].osc.clkdiv_C.cnt\[12\] _01574_ _01578_ genblk1\[4\].osc.clkdiv_C.cnt\[16\]
+ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__a2bb2o_1
X_08428_ _03129_ _03133_ _03010_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06294__A _01255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08359_ _03060_ _03065_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__xor2_1
XANTENNA__08047__A2 _01666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11370_ genblk2\[7\].wave_shpr.div.i\[1\] genblk2\[7\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _05350_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07053__A1_N genblk1\[8\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10321_ _04628_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13040_ clknet_leaf_126_clk _00367_ net61 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10252_ net333 _04563_ _04564_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__a21oi_1
X_10183_ _04401_ _04367_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__or2b_1
X_12824_ clknet_leaf_62_clk _00157_ net189 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12067__B1 _05815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ clknet_leaf_52_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[14\] net110 VGND
+ VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10093__A2 _04452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ genblk2\[9\].wave_shpr.div.b1\[13\] genblk2\[9\].wave_shpr.div.acc\[13\]
+ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__and2b_1
XFILLER_0_126_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ clknet_leaf_119_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[17\] net141 VGND
+ VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_1
X_11637_ genblk2\[8\].wave_shpr.div.acc\[22\] _05411_ VGND VGND VPWR VPWR _05538_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11568_ genblk2\[8\].wave_shpr.div.acc\[4\] _05486_ _05417_ VGND VGND VPWR VPWR _05487_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08994__B1 _01157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold708 genblk2\[4\].wave_shpr.div.acc\[17\] VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13307_ clknet_leaf_122_clk _00628_ net137 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold719 genblk2\[4\].wave_shpr.div.acc\[2\] VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__dlygate4sd3_1
X_10519_ genblk2\[4\].wave_shpr.div.acc\[25\] _04751_ VGND VGND VPWR VPWR _04753_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07747__B _01172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11499_ net709 _05442_ _05446_ net871 VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13238_ clknet_leaf_11_clk net236 net57 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13169_ clknet_leaf_127_clk _00494_ net66 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09454__S _00007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07730_ _01188_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07661_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _01190_ _01235_ genblk1\[10\].osc.clkdiv_C.cnt\[6\]
+ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__o22ai_1
XANTENNA__06524__A2 _01231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07721__A1 genblk1\[1\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09400_ genblk2\[1\].wave_shpr.div.acc\[7\] genblk2\[1\].wave_shpr.div.b1\[7\] VGND
+ VGND VPWR VPWR _03964_ sky130_fd_sc_hd__or2b_1
X_06612_ genblk1\[3\].osc.clkdiv_C.cnt\[1\] _01519_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__xor2_1
XANTENNA__08594__A net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07592_ _02298_ _02269_ _02272_ _02267_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_88_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09331_ _03790_ _03911_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__xnor2_1
X_06543_ _01452_ _01461_ _01462_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_5_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09262_ net454 _03835_ _03838_ net476 _03860_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__a221o_1
X_06474_ net29 _01403_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08213_ _02917_ _02916_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__xnor2_1
X_09193_ _03824_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_889 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09226__B2 net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08144_ genblk1\[3\].osc.clkdiv_C.cnt\[15\] _01576_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08075_ genblk1\[5\].osc.clkdiv_C.cnt\[8\] _01678_ _01726_ genblk1\[5\].osc.clkdiv_C.cnt\[9\]
+ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07026_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01846_ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold13 genblk2\[7\].wave_shpr.div.quo\[19\] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _03519_ _03662_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__xnor2_1
Xhold24 _00634_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 genblk2\[5\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 _00813_ VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 genblk2\[2\].wave_shpr.div.quo\[7\] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _02632_ _02633_ _02634_ genblk1\[8\].osc.clkdiv_C.cnt\[17\] genblk1\[8\].osc.clkdiv_C.cnt\[16\]
+ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__a311oi_2
Xhold68 PWM.final_sample_in\[7\] VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 _00395_ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06289__A _01246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07859_ _02563_ _02564_ _02565_ _02509_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10870_ _04967_ _05013_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09529_ net537 _04052_ _04053_ net645 _04054_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12540_ clknet_leaf_62_clk _00092_ net189 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12471_ clknet_leaf_31_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[5\] net100 VGND VGND
+ VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.cnt\[5\] sky130_fd_sc_hd__dfrtp_1
X_11422_ genblk2\[8\].wave_shpr.div.b1\[12\] genblk2\[8\].wave_shpr.div.acc\[12\]
+ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__and2b_1
XANTENNA__07228__B1 _01227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07779__A1 _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11353_ _05218_ _05273_ _05336_ genblk2\[7\].wave_shpr.div.acc\[21\] VGND VGND VPWR
+ VPWR _05339_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_104_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10304_ genblk2\[4\].wave_shpr.div.b1\[17\] genblk2\[4\].wave_shpr.div.acc\[17\]
+ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__and2b_1
X_11284_ _05179_ _05189_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__xor2_1
XANTENNA__08728__B1 _02224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13023_ clknet_leaf_113_clk _00350_ net128 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_10235_ _04552_ _04549_ _04553_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09782__B _01490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10166_ _04393_ _04371_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__or2b_1
XANTENNA__08398__B _01349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10097_ _04269_ genblk1\[3\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12807_ clknet_leaf_59_clk _00140_ net187 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10999_ _04985_ _05087_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12738_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[15\] net114 VGND
+ VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_2
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12669_ clknet_leaf_90_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[0\] net173 VGND VGND
+ VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06190_ net642 net361 VGND VGND VPWR VPWR PWM.next_counter\[1\] sky130_fd_sc_hd__xor2_1
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold505 genblk2\[10\].wave_shpr.div.quo\[4\] VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07477__B _02153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08431__A2 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold516 genblk2\[4\].wave_shpr.div.i\[2\] VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 genblk2\[5\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 genblk2\[6\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 genblk2\[11\].wave_shpr.div.quo\[4\] VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__buf_1
XFILLER_0_110_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08900_ sig_norm.acc\[2\] _03596_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _04186_ _04299_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__xnor2_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07493__A modein.delay_in\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _03531_ _03536_ _03537_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__and3_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12279__A0 _01308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ genblk2\[3\].wave_shpr.div.fin_quo\[0\] _02539_ _02939_ VGND VGND VPWR VPWR
+ _03469_ sky130_fd_sc_hd__a21o_1
X_07713_ _02414_ _02417_ _02419_ VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__a21bo_1
X_08693_ _03398_ _03399_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout176_A net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11743__A _02203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07940__B _02364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07644_ _02350_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__buf_2
XFILLER_0_76_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07575_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01925_ _02280_ _02281_ VGND VGND VPWR
+ VPWR _02282_ sky130_fd_sc_hd__a211o_1
X_09314_ genblk2\[0\].wave_shpr.div.acc\[10\] _03898_ _03889_ VGND VGND VPWR VPWR
+ _03899_ sky130_fd_sc_hd__mux2_1
X_06526_ _01451_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09245_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__and2_1
X_06457_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] _01387_ genblk1\[1\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09176_ genblk2\[10\].wave_shpr.div.b1\[1\] _01368_ _03722_ VGND VGND VPWR VPWR _03815_
+ sky130_fd_sc_hd__mux2_1
X_06388_ _01194_ _01176_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08127_ _02830_ _02827_ _02831_ _02829_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_133_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08058_ genblk1\[5\].osc.clkdiv_C.cnt\[6\] _01172_ _01180_ _02764_ VGND VGND VPWR
+ VPWR _02765_ sky130_fd_sc_hd__a31o_1
XFILLER_0_141_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07009_ _01823_ _01835_ _01836_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
X_10020_ genblk2\[3\].wave_shpr.div.acc\[21\] genblk2\[3\].wave_shpr.div.acc\[20\]
+ genblk2\[3\].wave_shpr.div.acc\[19\] _04415_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__or4_1
X_11971_ _05790_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__clkbuf_1
X_13710_ clknet_leaf_31_clk _01021_ net103 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10922_ net1301 _01811_ _05042_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__mux2_1
XANTENNA__07161__A2 genblk1\[9\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13641_ clknet_leaf_94_clk _00954_ net160 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10853_ _04976_ _04995_ _04996_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__a21o_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13572_ clknet_leaf_85_clk _00887_ net184 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10784_ net896 _04918_ _04922_ _04940_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__a22o_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11799__S _05613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12523_ clknet_leaf_103_clk PWM.next_counter\[7\] net157 VGND VGND VPWR VPWR PWM.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08661__A2 _02789_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12454_ clknet_leaf_39_clk net228 net115 VGND VGND VPWR VPWR modein.delay_octave_up_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11405_ _05372_ _05379_ _05380_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12385_ _05958_ _06060_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09071__C1 _03728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11336_ genblk2\[7\].wave_shpr.div.acc\[16\] _05326_ _05300_ VGND VGND VPWR VPWR
+ _05327_ sky130_fd_sc_hd__mux2_1
X_11267_ _05273_ _05182_ genblk2\[7\].wave_shpr.div.b1\[0\] VGND VGND VPWR VPWR _05274_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_120_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09374__A0 _03941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13006_ clknet_leaf_133_clk net581 net40 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10218_ net904 _04415_ _04541_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__a21bo_1
X_11198_ genblk2\[8\].wave_shpr.div.b1\[10\] _05239_ _05237_ VGND VGND VPWR VPWR _05240_
+ sky130_fd_sc_hd__mux2_1
X_10149_ net1057 _04486_ _04456_ _04489_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07688__B1 _02011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07360_ genblk1\[11\].osc.clkdiv_C.cnt\[7\] _02112_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06311_ genblk1\[0\].osc.clkdiv_C.cnt\[1\] genblk1\[0\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07291_ genblk1\[10\].osc.clkdiv_C.cnt\[15\] _02057_ VGND VGND VPWR VPWR _02058_
+ sky130_fd_sc_hd__and2_1
X_09030_ genblk2\[9\].wave_shpr.div.busy _03698_ net817 VGND VGND VPWR VPWR _03700_
+ sky130_fd_sc_hd__a21oi_1
X_06242_ genblk1\[0\].osc.clkdiv_C.cnt\[9\] _01193_ _01199_ _01202_ _01203_ VGND VGND
+ VPWR VPWR _01204_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06392__A _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06173_ _01141_ _01143_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__xor2_1
XFILLER_0_142_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold302 genblk2\[2\].wave_shpr.div.quo\[23\] VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold313 genblk2\[4\].wave_shpr.div.quo\[17\] VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 genblk2\[7\].wave_shpr.div.quo\[21\] VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 genblk2\[2\].wave_shpr.div.quo\[12\] VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 _00713_ VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 genblk2\[8\].wave_shpr.div.quo\[21\] VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ net605 _04336_ _04339_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__a21o_1
XANTENNA__11738__A _02248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold368 genblk2\[9\].wave_shpr.div.quo\[4\] VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 _00474_ VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _04178_ _04286_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__xnor2_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07915__A1 genblk1\[8\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _03445_ _03450_ _03516_ _03520_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__o211ai_2
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07915__B2 genblk1\[8\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1002 genblk1\[11\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR net1220 sky130_fd_sc_hd__clkbuf_2
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 genblk2\[9\].wave_shpr.div.b1\[10\] VGND VGND VPWR VPWR net1231 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _04247_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1024 genblk2\[11\].wave_shpr.div.b1\[6\] VGND VGND VPWR VPWR net1242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 genblk2\[7\].wave_shpr.div.b1\[10\] VGND VGND VPWR VPWR net1253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 _04631_ VGND VGND VPWR VPWR net1264 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ _03256_ _03257_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__nand2_1
Xhold1057 genblk2\[11\].wave_shpr.div.b1\[7\] VGND VGND VPWR VPWR net1275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 genblk2\[7\].wave_shpr.div.b1\[9\] VGND VGND VPWR VPWR net1286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 genblk2\[3\].wave_shpr.div.b1\[11\] VGND VGND VPWR VPWR net1297 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11475__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08676_ _03298_ _03333_ _03381_ _03382_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ genblk1\[11\].osc.clkdiv_C.cnt\[13\] _01209_ _01256_ genblk1\[11\].osc.clkdiv_C.cnt\[12\]
+ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__o22ai_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07558_ genblk2\[9\].wave_shpr.div.fin_quo\[4\] _02264_ VGND VGND VPWR VPWR _02265_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_36_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06509_ _01416_ _01365_ _01326_ genblk1\[2\].osc.clkdiv_C.cnt\[11\] genblk1\[2\].osc.clkdiv_C.cnt\[16\]
+ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07489_ _02147_ _02212_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__nor2_1
XANTENNA__10986__B1 _05054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09228_ _03835_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__clkbuf_4
X_09159_ genblk2\[0\].wave_shpr.div.fin_quo\[1\] genblk2\[0\].wave_shpr.div.quo\[0\]
+ _00001_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06406__A1 _01201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12170_ _05785_ genblk2\[10\].wave_shpr.div.acc\[25\] genblk2\[10\].wave_shpr.div.acc\[26\]
+ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__or3b_1
XFILLER_0_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06957__A2 _01227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11121_ genblk2\[7\].wave_shpr.div.acc\[2\] genblk2\[7\].wave_shpr.div.b1\[2\] VGND
+ VGND VPWR VPWR _05181_ sky130_fd_sc_hd__or2b_1
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold880 genblk2\[8\].wave_shpr.div.i\[1\] VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 genblk2\[1\].wave_shpr.div.acc\[21\] VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__dlygate4sd3_1
X_11052_ genblk2\[6\].wave_shpr.div.acc\[14\] _05128_ _05105_ VGND VGND VPWR VPWR
+ _05129_ sky130_fd_sc_hd__mux2_1
XANTENNA__11163__A0 genblk2\[7\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10003_ genblk2\[3\].wave_shpr.div.b1\[10\] genblk2\[3\].wave_shpr.div.acc\[10\]
+ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_13_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11466__A1 _02433_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11954_ genblk2\[10\].wave_shpr.div.b1\[15\] genblk2\[10\].wave_shpr.div.acc\[15\]
+ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10905_ _05036_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11885_ genblk2\[9\].wave_shpr.div.acc\[23\] _05610_ VGND VGND VPWR VPWR _05715_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13624_ clknet_leaf_68_clk _00937_ net194 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10836_ genblk2\[6\].wave_shpr.div.acc\[3\] genblk2\[6\].wave_shpr.div.b1\[3\] VGND
+ VGND VPWR VPWR _04980_ sky130_fd_sc_hd__or2b_1
XFILLER_0_39_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13555_ clknet_leaf_101_clk net587 net164 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10767_ genblk2\[5\].wave_shpr.div.acc\[14\] _04927_ _04907_ VGND VGND VPWR VPWR
+ _04928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08634__A2 genblk2\[8\].wave_shpr.div.fin_quo\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12506_ clknet_leaf_104_clk _00068_ net154 VGND VGND VPWR VPWR PWM.final_in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13486_ clknet_leaf_79_clk net405 net206 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10698_ net459 _02183_ _04856_ net471 _04876_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12437_ _05980_ _06088_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12368_ _06047_ _05950_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11319_ genblk2\[7\].wave_shpr.div.acc\[12\] _05313_ _05300_ VGND VGND VPWR VPWR
+ _05314_ sky130_fd_sc_hd__mux2_1
X_12299_ net430 _06009_ _06010_ _05982_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__a22o_1
X_06860_ net1229 _01715_ _01718_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09462__S _00007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06791_ genblk1\[5\].osc.clkdiv_C.cnt\[16\] _01578_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08530_ _03141_ _03236_ net3 net163 VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08461_ _02217_ _02553_ genblk2\[6\].wave_shpr.div.fin_quo\[4\] VGND VGND VPWR VPWR
+ _03168_ sky130_fd_sc_hd__and3_1
XFILLER_0_148_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07412_ genblk2\[1\].wave_shpr.div.i\[2\] genblk2\[1\].wave_shpr.div.i\[3\] genblk2\[1\].wave_shpr.div.i\[0\]
+ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08392_ genblk1\[2\].osc.clkdiv_C.cnt\[9\] _01431_ _03096_ _03097_ _03098_ VGND VGND
+ VPWR VPWR _03099_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07343_ _02092_ _02102_ _02103_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07274_ _02027_ _02046_ _02047_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_61_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09013_ _02171_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__buf_6
XFILLER_0_14_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06225_ _01176_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold110 genblk2\[7\].wave_shpr.div.i\[4\] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08389__B2 _02011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06156_ _01126_ _01127_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__or2_1
Xhold121 genblk2\[2\].wave_shpr.div.quo\[18\] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold132 _00882_ VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold143 PWM.counter\[0\] VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__buf_1
Xhold154 sig_norm.quo\[8\] VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 genblk2\[10\].wave_shpr.div.quo\[20\] VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 genblk2\[0\].wave_shpr.div.b1\[6\] VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 _00803_ VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold198 genblk2\[9\].wave_shpr.div.quo\[21\] VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _04202_ _04326_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10499__A2 _04715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09846_ genblk2\[2\].wave_shpr.div.acc_next\[0\] _04247_ _04250_ net259 _04274_ VGND
+ VGND VPWR VPWR _00316_ sky130_fd_sc_hd__a221o_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _03701_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__buf_4
X_06989_ genblk1\[7\].osc.clkdiv_C.cnt\[1\] genblk1\[7\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01824_ sky130_fd_sc_hd__xnor2_1
X_08728_ genblk2\[2\].wave_shpr.div.fin_quo\[4\] _03113_ _03117_ _02224_ VGND VGND
+ VPWR VPWR _03435_ sky130_fd_sc_hd__a31o_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _02939_ _03365_ _02943_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__o21ai_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11670_ genblk2\[9\].wave_shpr.div.acc\[9\] genblk2\[9\].wave_shpr.div.b1\[9\] VGND
+ VGND VPWR VPWR _05562_ sky130_fd_sc_hd__or2b_1
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10621_ genblk2\[6\].wave_shpr.div.b1\[4\] _04836_ _04834_ VGND VGND VPWR VPWR _04837_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13340_ clknet_leaf_7_clk _00661_ net49 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10552_ genblk2\[5\].wave_shpr.div.acc\[2\] genblk2\[5\].wave_shpr.div.b1\[2\] VGND
+ VGND VPWR VPWR _04780_ sky130_fd_sc_hd__or2b_1
XFILLER_0_91_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13271_ clknet_leaf_137_clk _00594_ net41 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10483_ genblk2\[4\].wave_shpr.div.acc\[14\] _04727_ _04704_ VGND VGND VPWR VPWR
+ _04728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12222_ _05933_ _05958_ _05959_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12153_ genblk2\[10\].wave_shpr.div.acc\[19\] _05900_ VGND VGND VPWR VPWR _05903_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11104_ genblk2\[7\].wave_shpr.div.acc\[17\] genblk2\[7\].wave_shpr.div.b1\[17\]
+ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__or2b_1
X_12084_ _05815_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__clkbuf_4
X_11035_ net900 _05086_ _05093_ _05115_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__a22o_1
XANTENNA__08001__B1 _01675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08552__A1 genblk2\[6\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12986_ clknet_leaf_13_clk _00315_ net69 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12100__A2 _05844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11937_ _03821_ genblk2\[10\].wave_shpr.div.acc\[6\] _05758_ VGND VGND VPWR VPWR
+ _05759_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10662__A2 _04853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11868_ net669 _05684_ _05685_ _05703_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10819_ genblk2\[5\].wave_shpr.div.busy _04962_ net855 VGND VGND VPWR VPWR _04964_
+ sky130_fd_sc_hd__a21oi_1
X_13607_ clknet_leaf_68_clk _00920_ net194 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11799_ genblk2\[9\].wave_shpr.div.acc\[1\] _05650_ _05613_ VGND VGND VPWR VPWR _05651_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13538_ clknet_leaf_100_clk _00853_ net165 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_40_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13469_ clknet_leaf_85_clk _00786_ net204 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07043__A1 genblk1\[8\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10192__A _04455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07043__B2 genblk1\[8\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07961_ genblk1\[7\].osc.clkdiv_C.cnt\[14\] _01360_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__or2_1
X_09700_ _04170_ _04178_ _04179_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__a21o_1
X_06912_ genblk1\[6\].osc.clkdiv_C.cnt\[1\] net837 genblk1\[6\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__a21oi_1
X_07892_ _02529_ _02594_ _02518_ _02598_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__and4_1
XANTENNA__09192__S _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08543__A1 _02225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09631_ net973 _04109_ _04113_ _04125_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06843_ net1072 _01705_ _01707_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__07932__C genblk2\[8\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09562_ genblk2\[1\].wave_shpr.div.b1\[0\] _04011_ net752 VGND VGND VPWR VPWR _04073_
+ sky130_fd_sc_hd__a21o_1
X_06774_ _01649_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[14\] sky130_fd_sc_hd__clkbuf_1
X_08513_ _03210_ _03214_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__or2b_1
XFILLER_0_77_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09493_ net1277 _04036_ _04024_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08444_ _03145_ _03149_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08059__B1 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08375_ _02600_ _03080_ net24 _02520_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__a211o_1
XANTENNA__10367__A _02152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07326_ _02074_ _02084_ _02088_ _02089_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__nand4_1
XFILLER_0_34_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07257_ _02027_ _02034_ _02035_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_116_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06208_ freq_div.state\[1\] freq_div.state\[2\] freq_div.state\[0\] VGND VGND VPWR
+ VPWR _01170_ sky130_fd_sc_hd__or3b_1
XFILLER_0_131_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07188_ genblk1\[9\].osc.clkdiv_C.cnt\[10\] _01974_ genblk1\[9\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06139_ _01107_ _01110_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__xor2_1
XFILLER_0_112_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07585__A2 _01311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09829_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__and2_1
X_12840_ clknet_leaf_65_clk net1306 net197 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ clknet_leaf_93_clk _00104_ net148 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ genblk2\[9\].wave_shpr.div.fin_quo\[0\] _05613_ _00023_ VGND VGND VPWR VPWR
+ _05614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ genblk2\[8\].wave_shpr.div.i\[1\] genblk2\[8\].wave_shpr.div.i\[0\] genblk2\[8\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout60 net63 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout71 net72 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10604_ genblk2\[5\].wave_shpr.div.fin_quo\[5\] net1330 _00015_ VGND VGND VPWR VPWR
+ _04827_ sky130_fd_sc_hd__mux2_1
XANTENNA__09798__B1 _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout82 net83 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
X_11584_ _05389_ _05498_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__xnor2_1
Xfanout93 net94 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13323_ clknet_leaf_26_clk _00644_ net87 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10535_ genblk2\[5\].wave_shpr.div.acc\[17\] genblk2\[5\].wave_shpr.div.b1\[17\]
+ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__or2b_1
XFILLER_0_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13254_ clknet_leaf_2_clk _00577_ net43 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10466_ net1008 _04683_ _04690_ _04714_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12205_ genblk2\[11\].wave_shpr.div.b1\[1\] genblk2\[11\].wave_shpr.div.acc\[1\]
+ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__or2b_1
X_13185_ clknet_leaf_112_clk _00510_ net128 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10397_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12136_ _05776_ _05733_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__or2b_1
XANTENNA__13081__RESET_B net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12067_ net446 _05812_ _05815_ genblk2\[10\].wave_shpr.div.quo\[23\] _05838_ VGND
+ VGND VPWR VPWR _00973_ sky130_fd_sc_hd__a221o_1
X_11018_ net826 _05086_ _05093_ _05102_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_138_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_138_clk sky130_fd_sc_hd__clkbuf_16
X_12969_ clknet_leaf_111_clk _00298_ net128 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06490_ genblk1\[2\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__inv_2
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10187__A _04451_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06384__B _01327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08160_ _01489_ genblk1\[3\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07111_ genblk1\[8\].osc.clkdiv_C.cnt\[15\] genblk1\[8\].osc.clkdiv_C.cnt\[14\] _01910_
+ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08091_ _02797_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__buf_2
XFILLER_0_141_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10915__A _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07042_ genblk1\[8\].osc.clkdiv_C.cnt\[1\] _01436_ _01855_ _01859_ genblk1\[8\].osc.clkdiv_C.cnt\[10\]
+ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__a32o_1
XFILLER_0_141_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11899__A1 _03839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08993_ _03572_ _03675_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07944_ genblk1\[7\].osc.clkdiv_C.cnt\[8\] _01920_ _01514_ genblk1\[7\].osc.clkdiv_C.cnt\[9\]
+ VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__o22a_1
XANTENNA__07319__A2 _01242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07875_ _02575_ _02580_ _02581_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__a21o_1
XANTENNA__11520__B1 _05449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09614_ net865 _04109_ _04080_ _04112_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__a22o_1
X_06826_ _01694_ _01695_ _01696_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__and3_1
X_09545_ net417 _04052_ _04053_ net426 _04063_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_129_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_129_clk sky130_fd_sc_hd__clkbuf_16
X_06757_ genblk1\[4\].osc.clkdiv_C.cnt\[10\] genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01627_
+ genblk1\[4\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09476_ _04026_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06575__A _01196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06688_ _01577_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__buf_4
XFILLER_0_136_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08427_ _03010_ _03129_ _03133_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__nor3_1
XFILLER_0_136_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10097__A _04269_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08358_ _02846_ _03064_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07309_ genblk1\[11\].osc.clkdiv_C.cnt\[7\] _01430_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08289_ _02993_ _02994_ _02995_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10320_ genblk2\[4\].wave_shpr.div.fin_quo\[4\] net1333 _00013_ VGND VGND VPWR VPWR
+ _04628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12000__A1 _03706_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10251_ net333 _04563_ _03855_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08014__B _01367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10182_ net791 _04486_ _04490_ _04514_ VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__a22o_1
XANTENNA__12303__A2 _06009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06518__B1 _01439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07572__C _01437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11511__B1 _05449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11484__A1_N _03727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09180__A1 _01356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12823_ clknet_leaf_62_clk _00156_ net189 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12474__RESET_B net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10078__B1 _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06485__A _01241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12754_ clknet_leaf_51_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[13\] net110 VGND
+ VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_2
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _05559_ _05595_ _05596_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__a21o_1
X_12685_ clknet_leaf_119_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[16\] net141 VGND
+ VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_2
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11290__A2 _05279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11636_ _05449_ _05536_ _05537_ _05448_ net456 VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__a32o_1
XFILLER_0_142_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11567_ _05485_ _05381_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10518_ net777 _04657_ _04655_ _04752_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__a22o_1
X_13306_ clknet_leaf_3_clk _00627_ net51 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold709 genblk2\[5\].wave_shpr.div.acc\[8\] VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__dlygate4sd3_1
X_11498_ genblk2\[8\].wave_shpr.div.quo\[1\] _05442_ _05446_ net743 VGND VGND VPWR
+ VPWR _00796_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13237_ clknet_leaf_10_clk _00560_ net57 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13262__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10449_ net971 _04683_ _04690_ _04701_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09735__S _00009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13168_ clknet_leaf_127_clk _00493_ net66 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11750__B1 _05624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06889__A2_N _01519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12119_ _05768_ _05737_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__or2b_1
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13099_ clknet_leaf_137_clk _00426_ net42 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09036__A _03702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06509__B1 _01326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11502__B1 _05446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07660_ _02359_ _02360_ _02363_ _02366_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06611_ _01186_ _01354_ _01171_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__o21a_2
XANTENNA__07721__A2 _02425_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07591_ _01928_ _01801_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__nor2_1
XANTENNA__08594__B _02364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09330_ _03791_ _03749_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__or2b_1
X_06542_ genblk1\[2\].osc.clkdiv_C.cnt\[6\] _01459_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09261_ _03853_ genblk1\[0\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__and2_1
X_06473_ genblk1\[1\].osc.clkdiv_C.cnt\[14\] _01401_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__and2_1
XANTENNA__08682__B1 _02224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08212_ _02697_ _02698_ _02746_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09192_ net1244 _02002_ _03822_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09226__A2 _03836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08143_ genblk2\[3\].wave_shpr.div.fin_quo\[6\] VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07237__A1 _01242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08434__B1 _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07237__B2 _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08074_ _02763_ _02765_ _02769_ _02778_ _02780_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__o41a_1
XFILLER_0_113_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07025_ _01822_ _01845_ _01846_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_12_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_129_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10380__A _04651_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold14 _00731_ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _03656_ _03523_ _03521_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__o21a_1
Xhold25 genblk2\[9\].wave_shpr.div.quo\[12\] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 _00549_ VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__A2 _01514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold47 genblk2\[0\].wave_shpr.div.quo\[21\] VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 _00299_ VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _01200_ genblk1\[8\].osc.clkdiv_C.cnt\[14\] _01362_ genblk1\[8\].osc.clkdiv_C.cnt\[15\]
+ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__a211o_1
Xhold69 PWM.next_pwm_out VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06289__B _01250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07858_ _02216_ _02552_ genblk2\[0\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR
+ _02565_ sky130_fd_sc_hd__and3_1
X_06809_ _01676_ _01677_ _01679_ _01680_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__or4b_1
X_07789_ genblk1\[0\].osc.clkdiv_C.cnt\[11\] _01263_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09528_ _03853_ genblk1\[1\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__and2_1
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09459_ _04017_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12470_ clknet_leaf_33_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[4\] net100 VGND VGND
+ VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.cnt\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__13773__RESET_B net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11421_ _05364_ _05395_ _05396_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__a21o_1
XANTENNA__10232__B1 _04457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11352_ net679 _05311_ _05315_ _05338_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10303_ _04566_ _04613_ _04614_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_120_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11283_ net877 _05279_ _05283_ _05286_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold967_A genblk1\[8\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13022_ clknet_leaf_128_clk _00349_ net67 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_10234_ genblk2\[3\].wave_shpr.div.acc\[24\] _04480_ _04549_ VGND VGND VPWR VPWR
+ _04553_ sky130_fd_sc_hd__or3b_1
X_10165_ net890 _04486_ _04490_ _04501_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07951__A2 _01556_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10096_ _04451_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12806_ clknet_leaf_59_clk _00139_ net187 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10998_ genblk2\[6\].wave_shpr.div.b1\[2\] genblk2\[6\].wave_shpr.div.acc\[2\] VGND
+ VGND VPWR VPWR _05087_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11263__A2 _05245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12737_ clknet_leaf_37_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[14\] net114 VGND
+ VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_2
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12668_ clknet_leaf_24_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[17\] net92 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11619_ net991 _05507_ _05445_ _05525_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12599_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[2\] net97 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_106_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold506 genblk2\[10\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold517 _00514_ VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11995__S _05802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold528 genblk2\[9\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold539 genblk2\[1\].wave_shpr.div.i\[2\] VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07927__C1 genblk1\[8\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _03482_ _03530_ _03529_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07942__A2 _01311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ net10 _02744_ _03467_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__and3_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07712_ _02418_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__buf_2
X_08692_ _03187_ _03194_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__xnor2_1
X_07643_ genblk1\[11\].osc.clkdiv_C.cnt\[16\] genblk1\[11\].osc.clkdiv_C.cnt\[17\]
+ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout169_A net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07574_ _01336_ _01437_ _01226_ genblk1\[9\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR
+ VPWR _02281_ sky130_fd_sc_hd__o31a_1
X_09313_ _03782_ _03897_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__xnor2_1
X_06525_ _01450_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__buf_2
XFILLER_0_8_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_60_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_118_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09244_ net543 _03845_ _03847_ genblk2\[0\].wave_shpr.div.quo\[14\] _03850_ VGND
+ VGND VPWR VPWR _00138_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06456_ genblk1\[1\].osc.clkdiv_C.cnt\[8\] genblk1\[1\].osc.clkdiv_C.cnt\[7\] _01387_
+ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__and3_1
XANTENNA__07949__A _01172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09175_ _03814_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06681__A2 _01362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06387_ genblk1\[1\].osc.clkdiv_C.cnt\[3\] _01323_ _01329_ _01330_ VGND VGND VPWR
+ VPWR _01331_ sky130_fd_sc_hd__a22o_1
X_08126_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] _01340_ _02829_ VGND VGND VPWR VPWR _02833_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09080__B1 _03733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08057_ genblk1\[5\].osc.clkdiv_C.cnt\[7\] _01223_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07008_ genblk1\[7\].osc.clkdiv_C.cnt\[7\] _01832_ genblk1\[7\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11190__A1 _03831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08959_ sig_norm.quo\[4\] _03647_ _02248_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__mux2_1
X_11970_ genblk2\[10\].wave_shpr.div.fin_quo\[2\] net220 _00003_ VGND VGND VPWR VPWR
+ _05790_ sky130_fd_sc_hd__mux2_1
X_10921_ _05045_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13640_ clknet_leaf_94_clk net683 net160 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10852_ genblk2\[6\].wave_shpr.div.b1\[7\] genblk2\[6\].wave_shpr.div.acc\[7\] VGND
+ VGND VPWR VPWR _04996_ sky130_fd_sc_hd__and2b_1
XFILLER_0_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10783_ _04938_ _04939_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__nand2_1
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ clknet_leaf_56_clk _00886_ net182 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_51_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08110__A2 _01313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12522_ clknet_leaf_103_clk PWM.next_counter\[6\] net156 VGND VGND VPWR VPWR PWM.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12453_ clknet_leaf_42_clk net5 net123 VGND VGND VPWR VPWR modein.delay_octave_up_in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07578__B _01234_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11404_ genblk2\[8\].wave_shpr.div.b1\[3\] genblk2\[8\].wave_shpr.div.acc\[3\] VGND
+ VGND VPWR VPWR _05380_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12384_ _05959_ _05933_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__or2b_1
XFILLER_0_62_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09071__B1 _01302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11335_ _05325_ _05212_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11266_ _05219_ _05220_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__nor2_2
XFILLER_0_120_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09374__A1 _03942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10217_ genblk2\[3\].wave_shpr.div.acc\[19\] _04538_ VGND VGND VPWR VPWR _04541_
+ sky130_fd_sc_hd__or2_1
X_13005_ clknet_leaf_138_clk _00334_ net40 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11197_ _01859_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__inv_2
XANTENNA__11181__A1 _03819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10148_ net976 _04488_ _04420_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__mux2_1
XANTENNA__11844__A _03693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10079_ _03833_ net1227 VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13769_ clknet_leaf_71_clk _01080_ net217 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_42_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_16
X_06310_ genblk1\[0\].osc.clkdiv_C.cnt\[1\] genblk1\[0\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01271_ sky130_fd_sc_hd__or2_1
X_07290_ _02027_ _02056_ _02057_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_57_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06241_ _01201_ genblk1\[0\].osc.clkdiv_C.cnt\[7\] genblk1\[0\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06172_ _01141_ _01143_ _01119_ _01126_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_53_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08404__A3 _01362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold303 genblk2\[10\].wave_shpr.div.quo\[13\] VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold314 _00476_ VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold325 genblk2\[0\].wave_shpr.div.quo\[15\] VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold336 _00303_ VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold347 genblk2\[9\].wave_shpr.div.quo\[23\] VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 genblk2\[11\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09931_ _04210_ net22 VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__nor2_1
Xhold369 _00870_ VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _04179_ _04170_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__or2b_1
XANTENNA__06690__A2_N _01209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08813_ _03511_ _03515_ _03513_ _03514_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__o211ai_2
Xhold1003 _01059_ VGND VGND VPWR VPWR net1221 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09969__B_N genblk2\[3\].wave_shpr.div.b1\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 genblk2\[4\].wave_shpr.div.b1\[10\] VGND VGND VPWR VPWR net1232 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _02164_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 genblk2\[0\].wave_shpr.div.b1\[1\] VGND VGND VPWR VPWR net1243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 genblk2\[10\].wave_shpr.div.b1\[7\] VGND VGND VPWR VPWR net1254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 genblk2\[11\].wave_shpr.div.b1\[3\] VGND VGND VPWR VPWR net1265 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _03422_ _03427_ _03449_ _03450_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__a211oi_2
Xhold1058 genblk2\[0\].wave_shpr.div.b1\[9\] VGND VGND VPWR VPWR net1276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1069 genblk2\[5\].wave_shpr.div.b1\[4\] VGND VGND VPWR VPWR net1287 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _03359_ _03380_ _03379_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__o21a_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07626_ _02081_ _01241_ _02331_ _02332_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__a211o_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06351__A1 genblk1\[0\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07557_ genblk2\[9\].wave_shpr.div.fin_quo\[3\] _02263_ VGND VGND VPWR VPWR _02264_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_33_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_16
X_06508_ _01201_ _01410_ _01432_ _01412_ genblk1\[2\].osc.clkdiv_C.cnt\[7\] VGND VGND
+ VPWR VPWR _01434_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07679__A _01489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07488_ genblk2\[11\].wave_shpr.div.busy _02211_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09840__A2 _04247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06439_ genblk1\[1\].osc.clkdiv_C.cnt\[3\] _01378_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__and2_1
X_09227_ net277 _03836_ _03840_ net379 VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09158_ _03805_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08109_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01323_ _02811_ _02815_ VGND VGND VPWR
+ VPWR _02816_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06406__A2 genblk1\[1\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09089_ _03737_ modein.delay_octave_down_in\[1\] _01197_ _03738_ VGND VGND VPWR VPWR
+ _03740_ sky130_fd_sc_hd__or4_1
X_11120_ genblk2\[7\].wave_shpr.div.acc\[3\] genblk2\[7\].wave_shpr.div.b1\[3\] VGND
+ VGND VPWR VPWR _05180_ sky130_fd_sc_hd__or2b_1
Xhold870 sig_norm.b1\[3\] VGND VGND VPWR VPWR net1088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 genblk2\[3\].wave_shpr.div.b1\[5\] VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 genblk2\[2\].wave_shpr.div.i\[1\] VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ _05009_ _05127_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11163__A1 _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10002_ _04369_ _04396_ _04397_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11953_ _05734_ _05773_ _05774_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10904_ net1200 _01799_ _04848_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11884_ net892 _03696_ _03694_ _05714_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13623_ clknet_leaf_85_clk _00936_ net204 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11218__A2 _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10835_ genblk2\[6\].wave_shpr.div.acc\[4\] genblk2\[6\].wave_shpr.div.b1\[4\] VGND
+ VGND VPWR VPWR _04979_ sky130_fd_sc_hd__or2b_1
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_109_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13554_ clknet_leaf_100_clk _00869_ net164 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12451__CLK clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10766_ _04807_ _04926_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12505_ clknet_leaf_104_clk _00067_ net154 VGND VGND VPWR VPWR PWM.final_in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13485_ clknet_leaf_97_clk _00802_ net167 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10697_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12436_ net619 _06072_ _06073_ _06098_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12367_ _05951_ _05937_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__or2b_1
XFILLER_0_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11318_ _05204_ _05312_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__xnor2_1
X_12298_ _03941_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__buf_4
X_11249_ net400 _05255_ _05256_ net585 _05264_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09743__S _00009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06790_ genblk1\[5\].osc.clkdiv_C.cnt\[5\] net36 VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08460_ _03165_ _03166_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07411_ genblk2\[0\].wave_shpr.div.start VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__buf_8
XFILLER_0_148_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08391_ _01412_ _01302_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_15_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_18_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07499__A net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07342_ genblk1\[11\].osc.clkdiv_C.cnt\[3\] _02097_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11090__A0 _05054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07273_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _02041_ net1183 VGND VGND VPWR VPWR _02047_
+ sky130_fd_sc_hd__a21oi_1
X_09012_ genblk2\[9\].wave_shpr.div.i\[0\] _02202_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__nand2_1
X_06224_ _01179_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold100 _00718_ VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__dlygate4sd3_1
X_06155_ _01124_ _01125_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold111 genblk2\[8\].wave_shpr.div.quo\[9\] VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout201_A net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold122 genblk2\[1\].wave_shpr.div.quo\[22\] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 genblk2\[11\].wave_shpr.div.quo\[15\] VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 genblk2\[9\].wave_shpr.div.quo\[19\] VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09219__A _03838_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold155 genblk2\[10\].wave_shpr.div.quo\[14\] VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 genblk2\[11\].wave_shpr.div.b1\[14\] VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold177 smpl_rt_clkdiv.clkDiv_inst.cnt\[7\] VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 genblk2\[1\].wave_shpr.div.b1\[15\] VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _04203_ _04158_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__or2b_1
Xhold199 genblk2\[1\].wave_shpr.div.quo\[19\] VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09845_ _04269_ genblk1\[2\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__and2_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _04237_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__clkbuf_1
X_06988_ net1058 _01823_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07311__A2_N _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08727_ _03113_ _03117_ genblk2\[2\].wave_shpr.div.fin_quo\[4\] VGND VGND VPWR VPWR
+ _03434_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13546__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ genblk2\[3\].wave_shpr.div.fin_quo\[3\] _02467_ _03364_ _02592_ VGND VGND
+ VPWR VPWR _03365_ sky130_fd_sc_hd__a22o_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _02222_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__clkbuf_4
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _03275_ _03276_ _03295_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10620_ _01730_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10551_ genblk2\[5\].wave_shpr.div.acc\[3\] genblk2\[5\].wave_shpr.div.b1\[3\] VGND
+ VGND VPWR VPWR _04779_ sky130_fd_sc_hd__or2b_1
XFILLER_0_52_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13270_ clknet_leaf_1_clk _00593_ net43 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10482_ _04609_ _04726_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12221_ genblk2\[11\].wave_shpr.div.b1\[9\] genblk2\[11\].wave_shpr.div.acc\[9\]
+ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__and2b_1
XANTENNA__11659__A _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12152_ net1135 _05876_ _05883_ _05902_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__a22o_1
X_11103_ net280 _05162_ _05163_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12083_ net969 _05844_ _05817_ _05849_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11034_ genblk2\[6\].wave_shpr.div.acc\[10\] _05114_ _05105_ VGND VGND VPWR VPWR
+ _05115_ sky130_fd_sc_hd__mux2_1
XANTENNA__07591__B _01801_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12985_ clknet_leaf_13_clk _00314_ net69 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09501__A1 _03831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09799__A _04250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11936_ _03821_ genblk2\[10\].wave_shpr.div.acc\[6\] _05757_ VGND VGND VPWR VPWR
+ _05758_ sky130_fd_sc_hd__o21a_1
XANTENNA__08907__S _01157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11867_ genblk2\[9\].wave_shpr.div.acc\[17\] _05702_ _05673_ VGND VGND VPWR VPWR
+ _05703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08068__A1 _01196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13606_ clknet_leaf_67_clk _00919_ net194 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10818_ _04855_ _04961_ _04963_ _04858_ net783 VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__a32o_1
XANTENNA__09804__A2 _04248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11798_ _05575_ _05649_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13537_ clknet_leaf_81_clk _00852_ net200 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10749_ genblk2\[5\].wave_shpr.div.acc\[10\] _04913_ _04907_ VGND VGND VPWR VPWR
+ _04914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13468_ clknet_leaf_75_clk _00785_ net203 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07766__B _01255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12419_ genblk2\[11\].wave_shpr.div.acc\[17\] _06086_ _05981_ VGND VGND VPWR VPWR
+ _06087_ sky130_fd_sc_hd__mux2_1
X_13399_ clknet_leaf_119_clk net318 net139 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07043__A2 _01487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09039__A _02147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07960_ genblk1\[7\].osc.clkdiv_C.cnt\[9\] _01514_ _02651_ _02665_ _02666_ VGND VGND
+ VPWR VPWR _02667_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_4_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_16
X_06911_ genblk1\[6\].osc.clkdiv_C.cnt\[2\] genblk1\[6\].osc.clkdiv_C.cnt\[1\] genblk1\[6\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__and3_1
X_07891_ _02509_ _02597_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__or2_1
X_09630_ genblk2\[1\].wave_shpr.div.acc\[16\] _04124_ _04095_ VGND VGND VPWR VPWR
+ _04125_ sky130_fd_sc_hd__mux2_1
X_06842_ genblk1\[5\].osc.clkdiv_C.cnt\[7\] _01705_ _01694_ VGND VGND VPWR VPWR _01707_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__06398__A _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06773_ _01599_ _01646_ _01648_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__and3_1
X_09561_ genblk2\[1\].wave_shpr.div.b1\[0\] net752 _04011_ VGND VGND VPWR VPWR _04072_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08512_ _03204_ _03217_ _03127_ _03218_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__o211a_1
X_09492_ _01411_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10102__A2 _04457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08443_ _03145_ _03149_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__xor2_2
XANTENNA_fanout151_A net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08374_ _02520_ net1354 _03080_ _02600_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12939__RESET_B net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07325_ genblk1\[11\].osc.clkdiv_C.cnt\[1\] _01321_ _01925_ genblk1\[11\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_129_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09271__A3 _03804_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07256_ genblk1\[10\].osc.clkdiv_C.cnt\[3\] _02032_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06207_ genblk1\[0\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10383__A _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07187_ genblk1\[9\].osc.clkdiv_C.cnt\[10\] _01974_ _01976_ _01954_ VGND VGND VPWR
+ VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o211a_1
XFILLER_0_103_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06138_ _01108_ _01109_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08534__A2 _02526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09828_ net393 _04257_ _04259_ net573 _04264_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__a221o_1
X_09759_ _04228_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ clknet_leaf_93_clk _00103_ net148 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _05612_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__buf_4
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _05449_ _05546_ _05547_ _05448_ net1098 VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__a32o_1
XANTENNA__08028__A genblk2\[6\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout50 net85 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
Xfanout61 net62 VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10603_ _04826_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__clkbuf_1
Xfanout72 net75 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09798__B2 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout83 net84 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_153_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11583_ _05390_ _05367_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__or2b_1
Xfanout94 net98 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13322_ clknet_leaf_26_clk _00643_ net87 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10534_ net281 _04761_ _04762_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13253_ clknet_leaf_1_clk _00576_ net41 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10465_ genblk2\[4\].wave_shpr.div.acc\[10\] _04713_ _04704_ VGND VGND VPWR VPWR
+ _04714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12204_ genblk2\[11\].wave_shpr.div.acc\[0\] genblk2\[11\].wave_shpr.div.b1\[0\]
+ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__and2b_1
XANTENNA__08222__A1 _02789_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13184_ clknet_leaf_112_clk _00509_ net129 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10396_ genblk2\[4\].wave_shpr.div.quo\[15\] _04661_ _04663_ net596 _04666_ VGND
+ VGND VPWR VPWR _00474_ sky130_fd_sc_hd__a221o_1
X_12135_ net944 _05876_ _05883_ _05889_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__a22o_1
XANTENNA__06784__A1 _01436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09293__S _03804_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12306__B1 _06010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12066_ _05835_ genblk1\[10\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR _05838_
+ sky130_fd_sc_hd__and2_1
X_11017_ genblk2\[6\].wave_shpr.div.acc\[6\] _05101_ _05023_ VGND VGND VPWR VPWR _05102_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12968_ clknet_leaf_111_clk _00297_ net130 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11919_ genblk2\[10\].wave_shpr.div.acc\[7\] genblk2\[10\].wave_shpr.div.b1\[7\]
+ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__or2b_1
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12899_ clknet_leaf_30_clk net341 net102 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07110_ genblk1\[8\].osc.clkdiv_C.cnt\[14\] _01910_ _01913_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08090_ net11 _02364_ _02365_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__and3_1
XANTENNA__07777__A genblk1\[0\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07041_ _01439_ _01576_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__nand2_2
XFILLER_0_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08992_ _03134_ _03571_ _03009_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__o21a_1
XANTENNA__10931__A _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07943_ genblk1\[7\].osc.clkdiv_C.cnt\[11\] _01925_ _02649_ VGND VGND VPWR VPWR _02650_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout199_A net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07874_ _02517_ _02579_ _02577_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__and3_1
XANTENNA__07724__B1 _01313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09613_ genblk2\[1\].wave_shpr.div.acc\[12\] _04111_ _04095_ VGND VGND VPWR VPWR
+ _04112_ sky130_fd_sc_hd__mux2_1
X_06825_ genblk1\[5\].osc.clkdiv_C.cnt\[1\] genblk1\[5\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01696_ sky130_fd_sc_hd__nand2_1
X_09544_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__and2_1
X_06756_ genblk1\[4\].osc.clkdiv_C.cnt\[10\] _01631_ _01635_ _01600_ VGND VGND VPWR
+ VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o211a_1
XFILLER_0_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09475_ genblk2\[2\].wave_shpr.div.b1\[5\] _01248_ _04024_ VGND VGND VPWR VPWR _04026_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06687_ _01576_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06575__B _01327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08426_ _03131_ _03132_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08357_ genblk2\[4\].wave_shpr.div.fin_quo\[5\] _02521_ _02838_ _03063_ VGND VGND
+ VPWR VPWR _03064_ sky130_fd_sc_hd__a211o_1
XFILLER_0_117_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_863 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07308_ genblk1\[11\].osc.clkdiv_C.cnt\[4\] _01513_ _02070_ _02071_ VGND VGND VPWR
+ VPWR _02072_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08288_ _02972_ _02991_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_833 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07239_ genblk1\[10\].osc.clkdiv_C.cnt\[10\] _01215_ VGND VGND VPWR VPWR _02021_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10250_ _03690_ _04562_ _04563_ VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__nor3_1
X_10181_ genblk2\[3\].wave_shpr.div.acc\[10\] _04513_ _04507_ VGND VGND VPWR VPWR
+ _04514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10052__S _04238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12822_ clknet_leaf_62_clk _00155_ net189 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09468__B1 _03733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10078__A1 _03714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12753_ clknet_leaf_51_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[12\] net110 VGND
+ VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06485__B _01337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ genblk2\[9\].wave_shpr.div.b1\[12\] genblk2\[9\].wave_shpr.div.acc\[12\]
+ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__and2b_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[15\] net141 VGND
+ VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_4
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11635_ genblk2\[8\].wave_shpr.div.acc\[21\] _05534_ VGND VGND VPWR VPWR _05537_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11566_ _05382_ _05371_ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__or2b_1
X_13305_ clknet_leaf_96_clk _00626_ net161 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08994__A2 _01099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10517_ _04750_ _04621_ _04751_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11497_ _05444_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__clkbuf_4
X_13236_ clknet_leaf_15_clk _00559_ net74 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10448_ genblk2\[4\].wave_shpr.div.acc\[6\] _04700_ _04623_ VGND VGND VPWR VPWR _04701_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13649__RESET_B net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13167_ clknet_leaf_123_clk net972 net76 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10379_ net251 _04652_ _04656_ net408 VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12118_ _05812_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__clkbuf_4
X_13098_ clknet_leaf_137_clk _00425_ net39 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12049_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__and2_1
XANTENNA__09036__B _01432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06610_ genblk1\[3\].osc.clkdiv_C.cnt\[10\] _01231_ _01515_ _01516_ _01517_ VGND
+ VGND VPWR VPWR _01518_ sky130_fd_sc_hd__o2111a_1
X_07590_ genblk1\[9\].osc.clkdiv_C.cnt\[9\] _01991_ _01923_ genblk1\[9\].osc.clkdiv_C.cnt\[10\]
+ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10069__A1 _04444_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06541_ genblk1\[2\].osc.clkdiv_C.cnt\[6\] _01459_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__and2_1
XANTENNA__09052__A _03689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06472_ genblk1\[1\].osc.clkdiv_C.cnt\[13\] _01399_ _01402_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__o21a_1
X_09260_ genblk2\[0\].wave_shpr.div.quo\[22\] _03835_ _03847_ net265 _03859_ VGND
+ VGND VPWR VPWR _00145_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08211_ _02916_ _02917_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__or2b_1
XFILLER_0_118_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09191_ _03823_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06693__B1 _01340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08142_ _02848_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07300__A _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08073_ _02761_ _02762_ _02779_ _02764_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout114_A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07024_ genblk1\[7\].osc.clkdiv_C.cnt\[14\] genblk1\[7\].osc.clkdiv_C.cnt\[13\] _01842_
+ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07954__B _01805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11741__A1 _02248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07945__B1 _01805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08131__A _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08975_ sig_norm.quo\[7\] VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__inv_2
Xhold15 genblk2\[5\].wave_shpr.div.quo\[19\] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 _00878_ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 genblk2\[4\].wave_shpr.div.quo\[18\] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _02607_ _02608_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__or2b_1
Xhold48 _00145_ VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 genblk2\[0\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dlygate4sd3_1
X_07857_ genblk2\[0\].wave_shpr.div.fin_quo\[0\] genblk2\[0\].wave_shpr.div.fin_quo\[1\]
+ _02510_ _02316_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__a31oi_1
XANTENNA__11492__A _05441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10600__S _00015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06808_ genblk1\[5\].osc.clkdiv_C.cnt\[15\] _01359_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__or2_1
XANTENNA__06586__A _01342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07788_ _02493_ _02494_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__or2_1
XANTENNA__11257__B1 _05249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09527_ _04046_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__buf_2
XFILLER_0_149_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06739_ _01600_ _01621_ _01622_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08122__B1 _01304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09458_ genblk2\[1\].wave_shpr.div.fin_quo\[5\] net414 _00007_ VGND VGND VPWR VPWR
+ _04017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08409_ genblk2\[2\].wave_shpr.div.fin_quo\[2\] _03115_ VGND VGND VPWR VPWR _03116_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_19_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09389_ net288 _03952_ _03953_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11420_ genblk2\[8\].wave_shpr.div.b1\[11\] genblk2\[8\].wave_shpr.div.acc\[11\]
+ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11351_ _05336_ _05337_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11980__A1 genblk2\[10\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10302_ _04449_ genblk2\[4\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR _04614_
+ sky130_fd_sc_hd__and2_1
X_11282_ genblk2\[7\].wave_shpr.div.acc\[3\] _05285_ _05222_ VGND VGND VPWR VPWR _05286_
+ sky130_fd_sc_hd__mux2_1
X_13021_ clknet_leaf_122_clk _00348_ net76 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10233_ genblk2\[3\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10164_ genblk2\[3\].wave_shpr.div.acc\[6\] _04500_ _04420_ VGND VGND VPWR VPWR _04501_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07951__A3 _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10095_ genblk2\[3\].wave_shpr.div.quo\[8\] _04452_ _04456_ net401 VGND VGND VPWR
+ VPWR _00383_ sky130_fd_sc_hd__a22o_1
XANTENNA__11496__B1 _05417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12805_ clknet_leaf_59_clk net544 net187 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_812 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10997_ _05051_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08113__B1 _01592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12624__RESET_B net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ clknet_leaf_37_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[13\] net114 VGND
+ VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09861__B1 _04252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12667_ clknet_leaf_24_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[16\] net88 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_25_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11618_ genblk2\[8\].wave_shpr.div.acc\[16\] _05524_ _05416_ VGND VGND VPWR VPWR
+ _05525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12598_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[1\] net97 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07120__A _01432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11549_ genblk2\[8\].wave_shpr.div.acc\[0\] _00020_ _05471_ net274 _05472_ VGND VGND
+ VPWR VPWR _00821_ sky130_fd_sc_hd__o221a_1
XFILLER_0_123_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold507 genblk2\[3\].wave_shpr.div.i\[2\] VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 genblk2\[7\].wave_shpr.div.quo\[10\] VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 genblk2\[6\].wave_shpr.div.b1\[14\] VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13219_ clknet_leaf_3_clk _00542_ net47 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07774__B _01215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07927__B1 _01362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09047__A _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ genblk2\[4\].wave_shpr.div.fin_quo\[0\] _02521_ _02838_ VGND VGND VPWR VPWR
+ _03467_ sky130_fd_sc_hd__a21o_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07711_ net2 net163 _02312_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__and3_1
X_08691_ _03340_ _03350_ _03349_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_79_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07642_ net33 VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__clkbuf_4
X_07573_ _02278_ _02279_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__nand2_1
XANTENNA__08104__B1 _01592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09312_ _03783_ _03753_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__or2b_1
X_06524_ _01410_ _01231_ _01413_ _01429_ _01449_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_146_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09510__A _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06666__B1 _01223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09243_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06455_ _01391_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[7\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__07949__B _02011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10656__A _04856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06386_ genblk1\[1\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__inv_2
X_09174_ genblk2\[10\].wave_shpr.div.b1\[0\] _03813_ _03722_ VGND VGND VPWR VPWR _03814_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08125_ _01570_ _01870_ _02829_ _02830_ _02831_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09080__A1 _03732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08056_ _02761_ _02762_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07007_ genblk1\[7\].osc.clkdiv_C.cnt\[8\] genblk1\[7\].osc.clkdiv_C.cnt\[7\] _01832_
+ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__and3_1
XANTENNA__12082__S _05787_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10391__A _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08958_ _03565_ _03646_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07501__A_N net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07909_ genblk1\[8\].osc.clkdiv_C.cnt\[11\] _01869_ _02613_ _02614_ _02615_ VGND
+ VGND VPWR VPWR _02616_ sky130_fd_sc_hd__o221a_1
X_08889_ sig_norm.acc\[11\] sig_norm.acc\[12\] _03591_ _03594_ VGND VGND VPWR VPWR
+ _03595_ sky130_fd_sc_hd__or4_1
X_10920_ genblk2\[7\].wave_shpr.div.b1\[11\] _02433_ _05042_ VGND VGND VPWR VPWR _05045_
+ sky130_fd_sc_hd__mux2_1
X_10851_ _04977_ _04993_ _04994_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13570_ clknet_leaf_56_clk net363 net182 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10782_ _04815_ _04880_ net630 VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ clknet_leaf_103_clk PWM.next_counter\[5\] net156 VGND VGND VPWR VPWR PWM.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12452_ clknet_leaf_116_clk net222 net150 VGND VGND VPWR VPWR modein.delay_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11403_ _05373_ _05377_ _05378_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12383_ net762 _06039_ _06040_ _06059_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__a22o_1
XANTENNA__09071__A1 _03726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09071__B2 _03727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11334_ _05213_ _05165_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07621__A2 _01430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11265_ _03819_ net1255 _00018_ genblk2\[7\].wave_shpr.div.acc\[0\] _05272_ VGND
+ VGND VPWR VPWR _00737_ sky130_fd_sc_hd__o221a_1
X_13004_ clknet_leaf_138_clk _00333_ net39 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10216_ net904 _04518_ _04522_ _04540_ VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__a22o_1
X_11196_ _05238_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11181__A2 _01242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10147_ _04383_ _04487_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10078_ _03714_ _04449_ _03736_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07688__A2 _01215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07115__A genblk1\[8\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_128_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13768_ clknet_leaf_71_clk _01079_ net217 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08637__A1 _02592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12719_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[14\] net181 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_127_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__10476__A _04654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13699_ clknet_leaf_94_clk _01010_ net160 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06240_ _01201_ genblk1\[0\].osc.clkdiv_C.cnt\[7\] genblk1\[0\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06171_ _01121_ _01123_ _01142_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold304 genblk2\[0\].wave_shpr.div.quo\[16\] VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 genblk2\[9\].wave_shpr.div.quo\[20\] VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold326 _00138_ VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 genblk2\[10\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 genblk2\[5\].wave_shpr.div.acc\[21\] VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ net605 _04315_ _04322_ _04338_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__a22o_1
Xhold359 genblk2\[0\].wave_shpr.div.b1\[15\] VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ net918 _04282_ _04252_ _04285_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__a22o_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ _03517_ _03518_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__or2b_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _04246_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__clkbuf_1
Xhold1004 genblk2\[8\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR net1222 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 genblk2\[6\].wave_shpr.div.b1\[11\] VGND VGND VPWR VPWR net1233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 genblk2\[10\].wave_shpr.div.b1\[8\] VGND VGND VPWR VPWR net1244 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _03447_ _03448_ _03445_ _03446_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__a211oi_4
Xhold1037 genblk1\[7\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR net1255 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__B genblk1\[9\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09505__A _04042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1048 genblk2\[5\].wave_shpr.div.b1\[11\] VGND VGND VPWR VPWR net1266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 genblk2\[2\].wave_shpr.div.b1\[12\] VGND VGND VPWR VPWR net1277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout181_A net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08325__B1 _02223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _03359_ _03379_ _03380_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__nor3_2
XFILLER_0_95_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ genblk1\[11\].osc.clkdiv_C.cnt\[13\] _01208_ _01576_ genblk1\[11\].osc.clkdiv_C.cnt\[15\]
+ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07556_ genblk2\[9\].wave_shpr.div.fin_quo\[2\] _02262_ VGND VGND VPWR VPWR _02263_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_76_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06507_ _01200_ _01432_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__nand2_2
XFILLER_0_118_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07487_ genblk2\[11\].wave_shpr.div.i\[1\] _02210_ genblk2\[11\].wave_shpr.div.i\[4\]
+ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__or3b_1
XANTENNA__06583__B _01250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10986__A2 _05051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09226_ genblk2\[0\].wave_shpr.div.quo\[7\] _03836_ _03840_ net269 VGND VGND VPWR
+ VPWR _00130_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06438_ _01373_ _01378_ _01379_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_106_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09157_ genblk2\[0\].wave_shpr.div.fin_quo\[0\] _03804_ _00001_ VGND VGND VPWR VPWR
+ _03805_ sky130_fd_sc_hd__mux2_1
X_06369_ _01192_ _01208_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__nand2_4
X_08108_ _02812_ _02809_ _02813_ _02814_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__or4_1
XFILLER_0_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09088_ _03737_ modein.delay_octave_down_in\[1\] _01591_ _03738_ VGND VGND VPWR VPWR
+ _03739_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08039_ _02741_ _02743_ _02745_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__o21a_1
Xhold860 genblk2\[11\].wave_shpr.div.acc\[25\] VGND VGND VPWR VPWR net1078 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout94_A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold871 genblk1\[0\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR net1089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 genblk2\[4\].wave_shpr.div.b1\[1\] VGND VGND VPWR VPWR net1100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 PWM.final_sample_in\[0\] VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ _05010_ _04969_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__or2b_1
XFILLER_0_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10001_ genblk2\[3\].wave_shpr.div.b1\[9\] genblk2\[3\].wave_shpr.div.acc\[9\] VGND
+ VGND VPWR VPWR _04397_ sky130_fd_sc_hd__and2b_1
XANTENNA__07772__D1 _02336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11952_ genblk2\[10\].wave_shpr.div.b1\[14\] genblk2\[10\].wave_shpr.div.acc\[14\]
+ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10903_ _05035_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11883_ net646 _05609_ _05713_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13622_ clknet_leaf_75_clk _00935_ net204 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10834_ genblk2\[6\].wave_shpr.div.acc\[5\] genblk2\[6\].wave_shpr.div.b1\[5\] VGND
+ VGND VPWR VPWR _04978_ sky130_fd_sc_hd__or2b_1
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13553_ clknet_leaf_100_clk net687 net164 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10765_ _04808_ _04766_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12504_ clknet_leaf_106_clk _00066_ net154 VGND VGND VPWR VPWR PWM.final_in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13484_ clknet_leaf_99_clk _00801_ net168 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10696_ genblk2\[5\].wave_shpr.div.quo\[22\] _02183_ _04856_ net245 _04875_ VGND
+ VGND VPWR VPWR _00565_ sky130_fd_sc_hd__a221o_1
XFILLER_0_152_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12435_ genblk2\[11\].wave_shpr.div.acc\[22\] _06096_ VGND VGND VPWR VPWR _06098_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12366_ net958 _06039_ _06040_ _06046_ VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11317_ _05205_ _05169_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__or2b_1
XFILLER_0_50_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12297_ _03942_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11248_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10362__B1 _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11179_ _03831_ net864 _03705_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_89_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07410_ _02154_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08390_ genblk1\[2\].osc.clkdiv_C.cnt\[8\] _01442_ _02011_ genblk1\[2\].osc.clkdiv_C.cnt\[7\]
+ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__a22o_1
XANTENNA__09807__B1 _04252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07341_ _02101_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__inv_2
XANTENNA__11090__A1 _05051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07272_ genblk1\[10\].osc.clkdiv_C.cnt\[8\] genblk1\[10\].osc.clkdiv_C.cnt\[7\] _02041_
+ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07833__A2 _02539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09011_ _03685_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06223_ _01184_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10934__A _05051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06154_ _01124_ _01125_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold101 genblk2\[8\].wave_shpr.div.i\[4\] VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold112 _00805_ VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _00230_ VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold134 _01049_ VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _00885_ VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 genblk2\[9\].wave_shpr.div.b1\[14\] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 genblk2\[6\].wave_shpr.div.quo\[23\] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 genblk2\[0\].wave_shpr.div.b1\[16\] VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ net1036 _04315_ _04322_ _04325_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__a22o_1
Xhold189 smpl_rt_clkdiv.clkDiv_inst.cnt\[5\] VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ net259 _04247_ _04250_ net520 _04273_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__a221o_1
XANTENNA__07962__B _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08010__A2 _01365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ genblk2\[3\].wave_shpr.div.b1\[10\] _02336_ _04039_ VGND VGND VPWR VPWR _04237_
+ sky130_fd_sc_hd__mux2_1
X_06987_ _01822_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__clkbuf_4
X_08726_ _03397_ _03400_ _03432_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__a21oi_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ genblk2\[3\].wave_shpr.div.fin_quo\[2\] _03363_ VGND VGND VPWR VPWR _03364_
+ sky130_fd_sc_hd__xnor2_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07608_ _02306_ _02311_ _02314_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__o21a_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _03293_ _03294_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07539_ PWM.final_sample_in\[1\] net1103 PWM.start VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10550_ _04776_ _04777_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09209_ _03714_ _03832_ _03736_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__o21ai_1
X_10481_ _04610_ _04568_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__or2b_1
XFILLER_0_17_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12220_ _05934_ _05956_ _05957_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12030__B1 _05817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08314__A _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12151_ _05900_ _05901_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10055__S _04238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11102_ net280 _05162_ _03855_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__o21ai_1
X_12082_ genblk2\[10\].wave_shpr.div.acc\[2\] _05848_ _05787_ VGND VGND VPWR VPWR
+ _05849_ sky130_fd_sc_hd__mux2_1
Xhold690 genblk2\[8\].wave_shpr.div.acc\[10\] VGND VGND VPWR VPWR net908 sky130_fd_sc_hd__dlygate4sd3_1
X_11033_ _05001_ _05113_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08001__A2 _01577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12984_ clknet_leaf_13_clk net262 net69 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11935_ _05742_ _05755_ _05756_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_115_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11866_ _05605_ _05701_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12344__B_N _03941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13605_ clknet_leaf_59_clk _00918_ net193 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_145_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10817_ _04962_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11797_ genblk2\[9\].wave_shpr.div.b1\[0\] _05573_ _05574_ VGND VGND VPWR VPWR _05649_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_131_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13536_ clknet_leaf_81_clk _00851_ net199 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10748_ _04799_ _04912_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13467_ clknet_leaf_75_clk _00784_ net203 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10679_ net249 _04861_ _04862_ net294 _04866_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12021__B1 _05787_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12418_ _05974_ _06085_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__xnor2_1
X_13398_ clknet_leaf_117_clk _00717_ net140 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12349_ genblk2\[11\].wave_shpr.div.acc\[1\] _05981_ VGND VGND VPWR VPWR _06033_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12891__RESET_B net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06910_ _01761_ _01762_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[1\]
+ sky130_fd_sc_hd__nor2_1
X_07890_ genblk2\[0\].wave_shpr.div.fin_quo\[7\] _02539_ _02596_ _02592_ VGND VGND
+ VPWR VPWR _02597_ sky130_fd_sc_hd__a22o_1
X_06841_ _01693_ _01705_ _01706_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
X_09560_ _03819_ genblk1\[1\].osc.clkdiv_C.cnt\[17\] _00006_ net752 _04071_ VGND VGND
+ VPWR VPWR _00233_ sky130_fd_sc_hd__o221a_1
X_06772_ _01647_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__inv_2
X_08511_ _03079_ _03126_ _03125_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__o21ai_1
X_09491_ _04035_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08442_ _02416_ _03148_ _02419_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__o21a_1
XFILLER_0_81_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08373_ _02599_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__inv_2
XANTENNA__08059__A2 _01238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout144_A net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07324_ genblk1\[11\].osc.clkdiv_C.cnt\[3\] _01334_ _02086_ _01197_ _02087_ VGND
+ VGND VPWR VPWR _02088_ sky130_fd_sc_hd__o221a_1
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07255_ genblk1\[10\].osc.clkdiv_C.cnt\[3\] _02032_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12355__S _05982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06206_ net399 _01166_ VGND VGND VPWR VPWR PWM.next_counter\[7\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07186_ genblk1\[9\].osc.clkdiv_C.cnt\[10\] _01974_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__nand2_1
X_06137_ net1 net7 VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__or2_1
XANTENNA__11495__A _05444_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07692__B _02011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09827_ _04058_ _01412_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__nor2_1
XANTENNA__12079__B1 _05817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09758_ genblk2\[3\].wave_shpr.div.b1\[2\] _04227_ _04039_ VGND VGND VPWR VPWR _04228_
+ sky130_fd_sc_hd__mux2_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout57_A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08709_ _03114_ _03415_ _03122_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__o21a_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09495__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09689_ genblk2\[2\].wave_shpr.div.acc\[4\] genblk2\[2\].wave_shpr.div.b1\[4\] VGND
+ VGND VPWR VPWR _04169_ sky130_fd_sc_hd__or2b_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _05610_ _05611_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ genblk2\[8\].wave_shpr.div.i\[1\] genblk2\[8\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _05547_ sky130_fd_sc_hd__nand2_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout40 net44 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_49_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08028__B genblk2\[6\].wave_shpr.div.fin_quo\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout51 net53 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_4
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout62 net63 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_4
X_10602_ genblk2\[5\].wave_shpr.div.fin_quo\[4\] net1326 _00015_ VGND VGND VPWR VPWR
+ _04826_ sky130_fd_sc_hd__mux2_1
XANTENNA__09798__A2 _04248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout73 net74 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_4
X_11582_ net978 _05447_ _05484_ _05497_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__a22o_1
Xfanout84 net85 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_2
Xfanout95 net98 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13321_ clknet_leaf_26_clk _00642_ net87 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10533_ net281 _04761_ _03855_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12265__S _05802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13252_ clknet_leaf_1_clk _00575_ net41 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10464_ _04601_ _04712_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12203_ genblk2\[11\].wave_shpr.div.acc\[1\] genblk2\[11\].wave_shpr.div.b1\[1\]
+ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13183_ clknet_leaf_112_clk _00508_ net129 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10395_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__and2_1
X_12134_ genblk2\[10\].wave_shpr.div.acc\[14\] _05888_ _05865_ VGND VGND VPWR VPWR
+ _05889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06784__A2 _01304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12306__B2 net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12065_ genblk2\[10\].wave_shpr.div.quo\[23\] _05812_ _05815_ net474 _05837_ VGND
+ VGND VPWR VPWR _00972_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11016_ _04993_ _05100_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12967_ clknet_leaf_111_clk net697 net130 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11918_ genblk2\[10\].wave_shpr.div.acc\[8\] genblk2\[10\].wave_shpr.div.b1\[8\]
+ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__or2b_1
XFILLER_0_59_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12898_ clknet_leaf_31_clk _00229_ net102 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07123__A _01432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11849_ _05598_ _05558_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__or2b_1
XFILLER_0_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09749__S _00009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13519_ clknet_leaf_79_clk _00836_ net206 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07040_ _01489_ _01344_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__nand2_4
XANTENNA__06472__A1 genblk1\[1\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11114__B_N genblk2\[7\].wave_shpr.div.b1\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08991_ _03674_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__clkbuf_1
X_07942_ genblk1\[7\].osc.clkdiv_C.cnt\[10\] _01311_ _01925_ genblk1\[7\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__o22a_1
XANTENNA__11264__B_N _05249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07873_ _02517_ _02577_ _02579_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__a21o_1
X_09612_ _03993_ _04110_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__xnor2_1
X_06824_ genblk1\[5\].osc.clkdiv_C.cnt\[1\] genblk1\[5\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01695_ sky130_fd_sc_hd__or2_1
XANTENNA__11762__B genblk1\[9\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09543_ net426 _04052_ _04053_ genblk2\[1\].wave_shpr.div.quo\[17\] _04062_ VGND
+ VGND VPWR VPWR _00225_ sky130_fd_sc_hd__a221o_1
X_06755_ genblk1\[4\].osc.clkdiv_C.cnt\[10\] _01631_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09477__A1 _01437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09474_ _04025_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06686_ _01575_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__buf_4
XFILLER_0_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08425_ _03011_ _03128_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08356_ _03061_ _03062_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__nor2_1
XANTENNA__06872__A _01441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07307_ genblk1\[11\].osc.clkdiv_C.cnt\[0\] _01223_ _01678_ VGND VGND VPWR VPWR _02071_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_144_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08287_ _02964_ _02958_ _02963_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06463__A1 genblk1\[1\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07238_ genblk1\[10\].osc.clkdiv_C.cnt\[12\] _02011_ _02012_ _02014_ _02019_ VGND
+ VGND VPWR VPWR _02020_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07169_ _01964_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10180_ _04398_ _04512_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07963__A1 _01200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11511__A2 _05448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12821_ clknet_leaf_67_clk net824 net196 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09468__A1 _03732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ clknet_leaf_50_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[11\] net111 VGND
+ VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11703_ _05560_ _05593_ _05594_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__a21o_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[14\] net81 VGND VGND
+ VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_84_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ genblk2\[8\].wave_shpr.div.acc\[21\] _05534_ VGND VGND VPWR VPWR _05536_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11565_ _05444_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13304_ clknet_leaf_96_clk _00625_ net161 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10516_ _04750_ _04748_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__nand2_1
X_11496_ net743 _05442_ _05417_ _05445_ VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__a22o_1
X_13235_ clknet_leaf_15_clk net250 net73 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10447_ _04593_ _04699_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13166_ clknet_leaf_127_clk _00491_ net79 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10378_ net408 _04652_ _04656_ net508 VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__a22o_1
X_12117_ net844 _05844_ _05850_ _05875_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__a22o_1
XANTENNA__11750__A2 _05623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13097_ clknet_leaf_137_clk _00424_ net41 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08221__B _02789_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12048_ net357 _05823_ _05825_ net373 _05828_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__a221o_1
XANTENNA__06509__A2 _01365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08903__B1 _01157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06676__B _01565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06540_ _01452_ _01459_ _01460_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__09052__B _01242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06471_ _01373_ _01401_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__nor2_1
X_08210_ _02315_ _02421_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__xor2_1
X_09190_ net1254 _03706_ _03822_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__mux2_1
XANTENNA_hold82_A genblk2\[2\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08141_ _02799_ _02847_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__xor2_2
XFILLER_0_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12844__D _00007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08072_ genblk1\[5\].osc.clkdiv_C.cnt\[6\] _01309_ _01180_ _02767_ _02766_ VGND VGND
+ VPWR VPWR _02779_ sky130_fd_sc_hd__a311o_1
XANTENNA__07300__B _01226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07023_ genblk1\[7\].osc.clkdiv_C.cnt\[13\] _01842_ genblk1\[7\].osc.clkdiv_C.cnt\[14\]
+ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10529__B1 _04657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout107_A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10153__S _04420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08974_ _03660_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08131__B _02837_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold16 _00563_ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 genblk2\[5\].wave_shpr.div.quo\[21\] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ _02609_ _02616_ _02629_ _02631_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__o22a_1
Xhold38 _00478_ VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 genblk2\[9\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__buf_1
XANTENNA__11773__A _04676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1124_A genblk2\[5\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07856_ genblk2\[0\].wave_shpr.div.fin_quo\[0\] net31 genblk2\[0\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__a21o_1
X_06807_ genblk1\[5\].osc.clkdiv_C.cnt\[9\] _01678_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__nor2_1
X_07787_ genblk1\[0\].osc.clkdiv_C.cnt\[8\] _01193_ _01184_ genblk1\[0\].osc.clkdiv_C.cnt\[9\]
+ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__a22o_1
XANTENNA__06586__B _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09526_ _04042_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__buf_2
X_06738_ genblk1\[4\].osc.clkdiv_C.cnt\[6\] _01616_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__or2_1
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09457_ _04016_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__clkbuf_1
X_06669_ _01349_ _01180_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__nand2_2
XFILLER_0_109_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08408_ genblk2\[2\].wave_shpr.div.fin_quo\[0\] genblk2\[2\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10480__A2 _04715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09388_ net288 _03952_ _03819_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_124_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08339_ genblk2\[6\].wave_shpr.div.fin_quo\[5\] _02467_ _02742_ VGND VGND VPWR VPWR
+ _03046_ sky130_fd_sc_hd__a21o_1
XANTENNA__10328__S _04440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10232__A2 _04454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11350_ genblk2\[7\].wave_shpr.div.acc\[20\] _05334_ VGND VGND VPWR VPWR _05337_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07633__B1 _01494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10301_ _04567_ _04611_ _04612_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11281_ _05187_ _05284_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__xnor2_1
X_13020_ clknet_leaf_123_clk _00347_ net77 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10232_ _04418_ _04454_ _04551_ _04457_ net1064 VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__a32o_1
XFILLER_0_30_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10163_ _04390_ _04499_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10940__B1 _05056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08041__B _01576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10094_ net401 _04452_ _04456_ net820 VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11999__B1_N _03705_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12804_ clknet_leaf_59_clk net496 net188 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12445__B1 _03944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10996_ _05055_ _05083_ _05085_ _05057_ net1165 VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__a32o_1
XFILLER_0_85_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12735_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[12\] net114 VGND
+ VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_2
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10471__A2 _04715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ clknet_leaf_25_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[15\] net88 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_154_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12664__RESET_B net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11617_ _05523_ _05405_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12597_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[0\] net97 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_154_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07120__B _01221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11548_ _03719_ genblk1\[8\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__or2_1
XANTENNA__07624__B1 _01172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold508 genblk2\[8\].wave_shpr.div.i\[2\] VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold519 genblk2\[3\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11479_ _05436_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13218_ clknet_leaf_5_clk _00541_ net46 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08232__A _02225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07927__A1 _01200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ clknet_leaf_121_clk net597 net80 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09047__B _02374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09762__S _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ genblk2\[10\].wave_shpr.div.fin_quo\[7\] _02362_ _02416_ VGND VGND VPWR VPWR
+ _02417_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07790__B _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08690_ _02798_ _03370_ _03375_ _03396_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__a31o_1
XANTENNA__06687__A _01576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07641_ _02330_ _02335_ _02343_ _02347_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_79_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07572_ genblk1\[9\].osc.clkdiv_C.cnt\[5\] _01186_ _01437_ _01225_ VGND VGND VPWR
+ VPWR _02279_ sky130_fd_sc_hd__or4_1
XFILLER_0_87_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09311_ net934 _03870_ _03877_ _03896_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__a22o_1
X_06523_ genblk1\[2\].osc.clkdiv_C.cnt\[10\] _01431_ _01448_ VGND VGND VPWR VPWR _01449_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10937__A _05054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09852__B2 _04248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09242_ genblk2\[0\].wave_shpr.div.quo\[14\] _03845_ _03847_ net495 _03849_ VGND
+ VGND VPWR VPWR _00137_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06454_ _01374_ _01389_ _01390_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08407__A _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09173_ _01342_ _01441_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__nor2_2
XANTENNA__10148__S _04420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06385_ _01326_ _01328_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__and2_2
XFILLER_0_44_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08124_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] _01340_ _01304_ genblk1\[4\].osc.clkdiv_C.cnt\[6\]
+ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__a22oi_1
XANTENNA__10214__A2 _04480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08055_ _01309_ _01180_ genblk1\[5\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _02762_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__07091__A1 genblk1\[8\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10672__A _04672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput17 net17 VGND VGND VPWR VPWR mode_out[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07006_ _01823_ _01834_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09238__A _03838_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08957_ _03506_ _03566_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__nor2_1
X_07908_ genblk1\[8\].osc.clkdiv_C.cnt\[10\] _01870_ _02610_ VGND VGND VPWR VPWR _02615_
+ sky130_fd_sc_hd__or3_1
XANTENNA__11478__A1 _01227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08888_ _03582_ _03581_ _03593_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__nor3_1
X_07839_ _02541_ _02545_ _02529_ _02518_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__and4b_1
X_10850_ genblk2\[6\].wave_shpr.div.b1\[6\] genblk2\[6\].wave_shpr.div.acc\[6\] VGND
+ VGND VPWR VPWR _04994_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09509_ _04044_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10781_ _04816_ _04880_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__or2_1
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12520_ clknet_leaf_104_clk PWM.next_counter\[4\] net157 VGND VGND VPWR VPWR PWM.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ clknet_4_0_0_clk net6 net38 VGND VGND VPWR VPWR modein.delay_in\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11402_ genblk2\[8\].wave_shpr.div.b1\[2\] genblk2\[8\].wave_shpr.div.acc\[2\] VGND
+ VGND VPWR VPWR _05378_ sky130_fd_sc_hd__and2b_1
XFILLER_0_90_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12382_ genblk2\[11\].wave_shpr.div.acc\[8\] _06058_ _06055_ VGND VGND VPWR VPWR
+ _06059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11333_ net1010 _05311_ _05315_ _05324_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11264_ net540 _05249_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__or2b_1
XANTENNA__07909__A1 genblk1\[8\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13003_ clknet_leaf_133_clk _00332_ net59 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10215_ _04538_ _04539_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__nand2_1
X_11195_ net1246 _05236_ _05237_ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__mux2_1
XANTENNA__11181__A3 _02064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10146_ _04384_ _04378_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__or2b_1
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06593__B1 _01500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10077_ net667 VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13767_ clknet_leaf_71_clk _01078_ net214 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10979_ _05074_ genblk1\[6\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12718_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[13\] net181 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
X_13698_ clknet_leaf_94_clk _01009_ net160 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12649_ clknet_leaf_10_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[16\] net55 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_111_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06170_ _01119_ _01126_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold305 genblk2\[6\].wave_shpr.div.quo\[7\] VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_810 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold316 genblk2\[7\].wave_shpr.div.quo\[24\] VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold327 genblk2\[3\].wave_shpr.div.quo\[20\] VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold338 genblk2\[9\].wave_shpr.div.acc\[21\] VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 genblk2\[6\].wave_shpr.div.quo\[20\] VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09058__A _02170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__13633__RESET_B net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09860_ genblk2\[2\].wave_shpr.div.acc\[2\] _04284_ _04214_ VGND VGND VPWR VPWR _04285_
+ sky130_fd_sc_hd__mux2_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _03512_ _03516_ _03223_ _03509_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__a211o_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _03833_ net1190 VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__and2_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 genblk2\[5\].wave_shpr.div.b1\[17\] VGND VGND VPWR VPWR net1223 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1016 genblk2\[7\].wave_shpr.div.b1\[17\] VGND VGND VPWR VPWR net1234 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ _03445_ _03446_ _03447_ _03448_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__o211a_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1027 genblk2\[3\].wave_shpr.div.b1\[4\] VGND VGND VPWR VPWR net1245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 genblk1\[2\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR net1256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 genblk2\[1\].wave_shpr.div.b1\[4\] VGND VGND VPWR VPWR net1267 sky130_fd_sc_hd__dlygate4sd3_1
X_08673_ _03357_ _03358_ _03334_ _03335_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06210__A _01171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout174_A net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07624_ genblk1\[11\].osc.clkdiv_C.cnt\[14\] _02085_ _01172_ VGND VGND VPWR VPWR
+ _02331_ sky130_fd_sc_hd__o21a_1
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12586__RESET_B net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07555_ genblk2\[9\].wave_shpr.div.fin_quo\[0\] genblk2\[9\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__or2_1
X_06506_ _01230_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__buf_8
XFILLER_0_118_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07836__B1 _02261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07486_ genblk2\[11\].wave_shpr.div.i\[2\] genblk2\[11\].wave_shpr.div.i\[3\] genblk2\[11\].wave_shpr.div.i\[0\]
+ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_76_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09225_ net269 _03836_ _03840_ net652 VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07041__A _01439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06437_ genblk1\[1\].osc.clkdiv_C.cnt\[1\] genblk1\[1\].osc.clkdiv_C.cnt\[0\] genblk1\[1\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09156_ _03803_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__buf_4
X_06368_ _01309_ _01221_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__and2_2
X_08107_ _01192_ _01208_ _01588_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__a21oi_1
X_09087_ modein.delay_octave_up_in\[1\] modein.delay_octave_up_in\[0\] VGND VGND VPWR
+ VPWR _03738_ sky130_fd_sc_hd__and2b_1
XANTENNA__10606__S _00015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_110_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_110_clk sky130_fd_sc_hd__clkbuf_16
X_06299_ _01176_ _01178_ _01194_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08038_ net12 _02744_ _02365_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__and3_2
Xhold850 genblk2\[4\].wave_shpr.div.acc\[3\] VGND VGND VPWR VPWR net1068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 genblk2\[3\].wave_shpr.div.i\[1\] VGND VGND VPWR VPWR net1079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 genblk2\[10\].wave_shpr.div.i\[1\] VGND VGND VPWR VPWR net1090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 genblk1\[3\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 _02252_ VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ _04370_ _04394_ _04395_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout87_A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09989_ _04378_ _04383_ _04384_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__a21o_1
XANTENNA__09513__B1 _04047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11951_ _05735_ _05771_ _05772_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__a21o_1
XANTENNA__11320__B1 _05283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10902_ net1250 _01923_ _04848_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__mux2_1
X_11882_ _05610_ _05611_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__and2b_1
X_10833_ genblk2\[6\].wave_shpr.div.acc\[6\] genblk2\[6\].wave_shpr.div.b1\[6\] VGND
+ VGND VPWR VPWR _04977_ sky130_fd_sc_hd__or2b_1
X_13621_ clknet_leaf_74_clk _00934_ net212 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10764_ net902 _04918_ _04922_ _04925_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__a22o_1
X_13552_ clknet_leaf_100_clk net650 net165 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12503_ clknet_leaf_106_clk _00065_ net154 VGND VGND VPWR VPWR PWM.final_in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13483_ clknet_leaf_99_clk _00800_ net168 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10695_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__and2_1
X_12434_ net955 _06072_ _06073_ _06097_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12365_ genblk2\[11\].wave_shpr.div.acc\[4\] _06045_ _05982_ VGND VGND VPWR VPWR
+ _06046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_101_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_101_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_105_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11316_ _05245_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12296_ _03687_ net409 _03735_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_10_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11247_ genblk2\[7\].wave_shpr.div.quo\[17\] _05255_ _05256_ net548 _05263_ VGND
+ VGND VPWR VPWR _00728_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11178_ net1216 VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10362__A1 _03726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10129_ net490 _04451_ _04455_ net529 _04475_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__a221o_1
XANTENNA__12032__A _02155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07678__A2_N _01215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11311__B1 _05283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06965__A _01213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09807__A1 genblk2\[2\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07340_ genblk1\[11\].osc.clkdiv_C.cnt\[3\] _02097_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07271_ _02045_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09010_ net1128 sig_norm.quo\[6\] _01154_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__mux2_1
X_06222_ _01172_ _01180_ _01183_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06153_ net3 _01100_ _01101_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold102 genblk2\[10\].wave_shpr.div.quo\[7\] VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold113 genblk2\[7\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 genblk2\[11\].wave_shpr.div.quo\[13\] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 genblk2\[10\].wave_shpr.div.quo\[16\] VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 smpl_rt_clkdiv.clkDiv_inst.cnt\[1\] VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 genblk2\[3\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold168 _00651_ VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09912_ genblk2\[2\].wave_shpr.div.acc\[14\] _04324_ _04301_ VGND VGND VPWR VPWR
+ _04325_ sky130_fd_sc_hd__mux2_1
Xhold179 genblk2\[11\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ _04269_ genblk1\[2\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__and2_1
XANTENNA__11765__B genblk1\[9\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _03831_ net614 _03733_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__a21bo_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ genblk1\[7\].osc.clkdiv_C.cnt\[2\] _01227_ _01793_ _01821_ VGND VGND VPWR
+ VPWR _01822_ sky130_fd_sc_hd__o211a_2
X_08725_ _03399_ _03398_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__and2b_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _03188_ _03189_ _02885_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__a21o_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_54_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07607_ _02313_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__buf_2
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _03237_ _03239_ _03243_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10397__A _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07538_ net1112 VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07469_ _02198_ VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09208_ net959 VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10480_ net850 _04715_ _04722_ _04725_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09139_ genblk2\[0\].wave_shpr.div.b1\[12\] genblk2\[0\].wave_shpr.div.acc\[12\]
+ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10336__S _04440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12030__A1 genblk2\[10\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12150_ _05781_ _05899_ genblk2\[10\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR
+ _05901_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11101_ _03690_ _05161_ _05162_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__nor3_1
XFILLER_0_130_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12081_ _05749_ _05847_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_127_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold680 genblk2\[8\].wave_shpr.div.acc\[5\] VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold691 genblk2\[8\].wave_shpr.div.acc\[12\] VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ _05002_ _04973_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__or2b_1
XANTENNA__10071__S _04440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09860__S _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12983_ clknet_leaf_125_clk _00312_ net69 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11934_ genblk2\[10\].wave_shpr.div.b1\[5\] genblk2\[10\].wave_shpr.div.acc\[5\]
+ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__and2b_1
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11865_ _05606_ _05554_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__or2b_1
X_13604_ clknet_leaf_97_clk _00003_ net166 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
X_10816_ genblk2\[5\].wave_shpr.div.i\[1\] genblk2\[5\].wave_shpr.div.i\[0\] genblk2\[5\].wave_shpr.div.i\[2\]
+ genblk2\[5\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__and4_1
XFILLER_0_95_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11796_ _03694_ _05647_ _05648_ _03696_ net1059 VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__a32o_1
XFILLER_0_54_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13535_ clknet_leaf_81_clk _00850_ net199 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10747_ _04800_ _04770_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__or2b_1
XFILLER_0_54_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10678_ _04672_ genblk1\[5\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__and2_1
X_13466_ clknet_leaf_75_clk _00783_ net203 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12021__A1 genblk2\[10\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12417_ _05975_ _05925_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__or2b_1
XANTENNA__12021__B2 _05816_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13397_ clknet_leaf_117_clk net662 net140 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12348_ _03944_ _06031_ _06032_ _03947_ net1044 VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__a32o_1
XFILLER_0_121_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12279_ _01308_ genblk2\[1\].wave_shpr.div.b1\[8\] _03719_ VGND VGND VPWR VPWR _06001_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06840_ genblk1\[5\].osc.clkdiv_C.cnt\[6\] _01703_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__nor2_1
XANTENNA__09770__S _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06771_ genblk1\[4\].osc.clkdiv_C.cnt\[14\] genblk1\[4\].osc.clkdiv_C.cnt\[13\] _01641_
+ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__and3_1
X_08510_ _03204_ _03205_ _03216_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__nor3b_2
XANTENNA__11805__S _05613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09490_ genblk2\[2\].wave_shpr.div.b1\[11\] _04034_ _04024_ VGND VGND VPWR VPWR _04035_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08441_ _02525_ _03146_ _03147_ _02361_ genblk2\[10\].wave_shpr.div.fin_quo\[3\]
+ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__a32o_1
XFILLER_0_93_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08372_ _03055_ _03077_ _03001_ _03078_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_46_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07323_ genblk1\[11\].osc.clkdiv_C.cnt\[3\] _01334_ _01321_ genblk1\[11\].osc.clkdiv_C.cnt\[1\]
+ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_73_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout137_A net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07254_ _02027_ _02032_ _02033_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_155_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08415__A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06205_ _01168_ VGND VGND VPWR VPWR PWM.next_counter\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10156__S _04420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07185_ _01953_ _01974_ _01975_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_143_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06136_ net1 net7 VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10680__A _04676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09192__A1 _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09826_ genblk2\[2\].wave_shpr.div.quo\[16\] _04257_ _04259_ net315 _04263_ VGND
+ VGND VPWR VPWR _00307_ sky130_fd_sc_hd__a221o_1
X_09757_ _01496_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__inv_2
X_06969_ _01179_ _01233_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__or2_2
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _03413_ _03414_ genblk2\[2\].wave_shpr.div.fin_quo\[4\] _02468_ VGND VGND
+ VPWR VPWR _03415_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12400__A _03942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09688_ genblk2\[2\].wave_shpr.div.acc\[5\] genblk2\[2\].wave_shpr.div.b1\[5\] VGND
+ VGND VPWR VPWR _04168_ sky130_fd_sc_hd__or2b_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _02685_ _02681_ _02686_ _02526_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__o31a_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08309__B _02361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ genblk2\[8\].wave_shpr.div.i\[1\] genblk2\[8\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _05546_ sky130_fd_sc_hd__or2_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout41 net43 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10601_ _04825_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__clkbuf_1
Xfanout52 net53 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_4
Xfanout63 net85 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
X_11581_ genblk2\[8\].wave_shpr.div.acc\[7\] _05496_ _05493_ VGND VGND VPWR VPWR _05497_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout74 net75 VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout85 net16 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10532_ _03690_ _04760_ _04761_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__nor3_1
XFILLER_0_52_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13320_ clknet_leaf_26_clk net499 net87 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout96 net98 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13251_ clknet_leaf_2_clk _00574_ net41 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10463_ _04602_ _04572_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__or2b_1
XANTENNA__10066__S _04440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09955__B1 _04253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12202_ genblk2\[11\].wave_shpr.div.b1\[2\] VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__inv_2
X_13182_ clknet_leaf_130_clk net473 net129 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10394_ net596 _04661_ _04663_ net637 _04665_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__a221o_1
X_12133_ _05773_ _05887_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08979__B _01157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12306__A2 _06009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12064_ _03833_ _01995_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__nor2_1
X_11015_ _04994_ _04977_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__or2b_1
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12966_ clknet_leaf_111_clk net337 net130 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11917_ genblk2\[10\].wave_shpr.div.acc\[9\] genblk2\[10\].wave_shpr.div.b1\[9\]
+ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__or2b_1
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ clknet_leaf_31_clk net258 net99 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07123__B _01344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11848_ net967 _05684_ _05685_ _05688_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__a22o_1
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11779_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06962__B _01797_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13518_ clknet_leaf_78_clk _00835_ net206 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13449_ clknet_leaf_91_clk _00766_ net144 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08749__A1 genblk2\[8\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09946__B1 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11753__B1 _05624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08990_ net1261 _03673_ _01158_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07941_ _02646_ _02647_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__nor2_2
XFILLER_0_76_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09174__A1 _03813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07872_ _02469_ _02578_ _02529_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__o21a_1
XANTENNA__07724__A2 _01323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09611_ _03994_ _03959_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__or2b_1
X_06823_ net1355 VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__inv_2
X_06754_ _01634_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[9\] sky130_fd_sc_hd__clkbuf_1
X_09542_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__and2_1
X_09473_ genblk2\[2\].wave_shpr.div.b1\[4\] _04023_ _04024_ VGND VGND VPWR VPWR _04025_
+ sky130_fd_sc_hd__mux2_1
X_06685_ _01194_ _01175_ _01191_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_90_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08424_ _03083_ _03124_ _03130_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08355_ genblk2\[4\].wave_shpr.div.fin_quo\[4\] _02932_ _02841_ _02222_ VGND VGND
+ VPWR VPWR _03062_ sky130_fd_sc_hd__a31o_1
XFILLER_0_129_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08437__B1 _02361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07306_ _01223_ _01678_ genblk1\[11\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR _02070_
+ sky130_fd_sc_hd__o21ai_1
X_08286_ _02964_ _02958_ _02963_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__nand3_1
XFILLER_0_61_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07237_ _01242_ _02015_ _02017_ _01197_ _02018_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__o221a_1
XFILLER_0_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07168_ _01954_ _01962_ _01963_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06119_ net365 _01088_ VGND VGND VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.next_cnt\[6\]
+ sky130_fd_sc_hd__xor2_1
X_07099_ genblk1\[8\].osc.clkdiv_C.cnt\[11\] _01904_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09809_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12820_ clknet_leaf_66_clk _00153_ net196 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ clknet_leaf_50_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[10\] net111 VGND
+ VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_2
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ genblk2\[9\].wave_shpr.div.b1\[11\] genblk2\[9\].wave_shpr.div.acc\[11\]
+ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__and2b_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[13\] net81 VGND VGND
+ VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ net1018 _05507_ _05445_ _05535_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11564_ net980 _05447_ _05446_ _05483_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11983__B1 _05796_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13303_ clknet_leaf_87_clk _00624_ net201 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10515_ genblk2\[4\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11495_ _05444_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_150_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10446_ _04594_ _04576_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__or2b_1
X_13234_ clknet_leaf_16_clk net295 net73 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13165_ clknet_leaf_127_clk _00490_ net68 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10377_ net508 _04652_ _04656_ net781 VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__a22o_1
XANTENNA__11204__A1_N _03727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12116_ genblk2\[10\].wave_shpr.div.acc\[10\] _05874_ _05865_ VGND VGND VPWR VPWR
+ _05875_ sky130_fd_sc_hd__mux2_1
X_13096_ clknet_leaf_137_clk _00423_ net41 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12452__RESET_B net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12047_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12949_ clknet_leaf_121_clk _00278_ net77 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06470_ genblk1\[1\].osc.clkdiv_C.cnt\[13\] genblk1\[1\].osc.clkdiv_C.cnt\[12\] _01398_
+ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07890__B2 _02592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08140_ _02838_ _02845_ _02846_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_43_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08071_ _02772_ _02774_ _02776_ _02777_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__o31a_1
XFILLER_0_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07022_ genblk1\[7\].osc.clkdiv_C.cnt\[13\] _01842_ _01844_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__06609__A2_N _01514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10529__A1 _04655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08973_ net1300 _03659_ _01158_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold17 genblk2\[5\].wave_shpr.div.quo\[17\] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 _00565_ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ _02609_ _02613_ _02630_ _02614_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__or4b_1
Xhold39 genblk2\[1\].wave_shpr.div.quo\[20\] VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09524__A _03853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07855_ _02509_ _02551_ _02554_ _02560_ _02518_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__o311a_1
X_06806_ _01336_ _01564_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__nor2_4
X_07786_ genblk1\[0\].osc.clkdiv_C.cnt\[8\] _01193_ _01184_ genblk1\[0\].osc.clkdiv_C.cnt\[9\]
+ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_79_866 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09525_ net645 _04048_ _04045_ net610 _04051_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11257__A2 _05245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06737_ _01620_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_63_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08122__A2 _01340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07979__A genblk2\[7\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09456_ genblk2\[1\].wave_shpr.div.fin_quo\[4\] net1316 _00007_ VGND VGND VPWR VPWR
+ _04016_ sky130_fd_sc_hd__mux2_1
X_06668_ genblk1\[4\].osc.clkdiv_C.cnt\[6\] _01557_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08407_ _02221_ _03113_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__nor2_2
X_06599_ _01441_ _01249_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__nor2_2
X_09387_ _03726_ _03951_ _03952_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__nor3_1
XFILLER_0_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08338_ _03043_ _03044_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_871 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08269_ _02973_ _02974_ _02975_ _02360_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10300_ genblk2\[4\].wave_shpr.div.b1\[15\] genblk2\[4\].wave_shpr.div.acc\[15\]
+ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__and2b_1
XFILLER_0_62_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_868 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11280_ _05188_ _05180_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__or2b_1
X_10231_ _04549_ _04550_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10162_ _04391_ _04372_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__or2b_1
XANTENNA__10940__B2 net792 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10093_ genblk2\[3\].wave_shpr.div.quo\[6\] _04452_ _04456_ net814 VGND VGND VPWR
+ VPWR _00381_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06496__C _01327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12803_ clknet_leaf_59_clk _00136_ net188 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10995_ _05023_ _05084_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_54_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08113__A2 _01323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12734_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[11\] net113 VGND
+ VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ clknet_leaf_25_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[14\] net86 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ _05406_ _05359_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__or2b_1
XFILLER_0_65_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12596_ clknet_leaf_15_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[17\] net73 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_80_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11547_ _05444_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__inv_2
Xhold509 genblk2\[0\].wave_shpr.div.b1\[5\] VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__dlygate4sd3_1
X_11478_ net1231 _01227_ _05433_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12633__RESET_B net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13217_ clknet_leaf_6_clk _00540_ net48 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10429_ net937 _04683_ _04656_ _04686_ VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08232__B _02885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07927__A2 genblk1\[8\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ clknet_leaf_121_clk _00473_ net81 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ clknet_leaf_125_clk _00406_ net61 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07790__C _01801_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08352__A2 _02521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07640_ _02335_ _02344_ _02345_ _02346_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07560__B1 _01328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07571_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01186_ _01355_ VGND VGND VPWR VPWR _02278_
+ sky130_fd_sc_hd__or3_1
XANTENNA__08104__A2 _01323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_16
X_09310_ genblk2\[0\].wave_shpr.div.acc\[9\] _03895_ _03889_ VGND VGND VPWR VPWR _03896_
+ sky130_fd_sc_hd__mux2_1
X_06522_ genblk1\[2\].osc.clkdiv_C.cnt\[10\] _01431_ _01447_ VGND VGND VPWR VPWR _01448_
+ sky130_fd_sc_hd__o21bai_1
XANTENNA__07312__B1 _01578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06453_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] _01387_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__or2_1
X_09241_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06666__A2 _01221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09172_ net1219 VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06384_ _01186_ _01327_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__nor2_4
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08123_ genblk1\[4\].osc.clkdiv_C.cnt\[5\] _01224_ _01249_ _01565_ genblk1\[4\].osc.clkdiv_C.cnt\[4\]
+ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__o32a_1
XFILLER_0_32_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout217_A net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08054_ genblk1\[5\].osc.clkdiv_C.cnt\[7\] _01223_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__or2_1
XANTENNA__09519__A _04042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07005_ genblk1\[7\].osc.clkdiv_C.cnt\[7\] _01832_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput18 net18 VGND VGND VPWR VPWR mode_out[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10164__S _04420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07039__A genblk1\[8\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_wire32_A _02302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10922__A1 _01811_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08956_ _03645_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__clkbuf_1
X_07907_ genblk1\[8\].osc.clkdiv_C.cnt\[8\] _01865_ _01859_ genblk1\[8\].osc.clkdiv_C.cnt\[9\]
+ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__o22a_1
X_08887_ sig_norm.b1\[0\] _03578_ _03592_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06597__B _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07838_ genblk2\[0\].wave_shpr.div.fin_quo\[5\] _02539_ _02509_ _02544_ VGND VGND
+ VPWR VPWR _02545_ sky130_fd_sc_hd__a211o_1
X_07769_ genblk1\[0\].osc.clkdiv_C.cnt\[13\] _01256_ _01240_ genblk1\[0\].osc.clkdiv_C.cnt\[12\]
+ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_36_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09508_ genblk2\[1\].wave_shpr.div.quo\[0\] _04043_ _04011_ _04045_ VGND VGND VPWR
+ VPWR _00207_ sky130_fd_sc_hd__a22o_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10780_ net630 _04918_ _04922_ _04937_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__a22o_1
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07303__B1 _01595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07502__A _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09439_ _03955_ _04001_ _04002_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__o21bai_1
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12450_ clknet_leaf_107_clk _00029_ net153 VGND VGND VPWR VPWR sig_norm.i\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11401_ _05374_ _05375_ _05376_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12381_ _05956_ _06057_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11332_ genblk2\[7\].wave_shpr.div.acc\[15\] _05323_ _05300_ VGND VGND VPWR VPWR
+ _05324_ sky130_fd_sc_hd__mux2_1
X_11263_ net540 _05245_ _05249_ net534 _05271_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13002_ clknet_leaf_133_clk _00331_ net59 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07909__A2 _01869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10214_ _04414_ _04480_ genblk2\[3\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR
+ _04539_ sky130_fd_sc_hd__o21ai_1
X_11194_ _03707_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10913__A1 _01819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10145_ _04451_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__06788__A _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10076_ _04448_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10103__A _04451_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13766_ clknet_leaf_69_clk _01077_ net213 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10978_ _04268_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12717_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[12\] net181 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13697_ clknet_leaf_96_clk _01008_ net160 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07131__B _01250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12648_ clknet_leaf_9_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[15\] net54 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12579_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[0\] net70 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_80_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold306 genblk2\[3\].wave_shpr.div.acc\[21\] VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08243__A _02225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold317 _00735_ VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold328 _00396_ VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 genblk2\[9\].wave_shpr.div.quo\[10\] VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10904__A1 _01799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08810_ _03223_ _03509_ _03512_ _03516_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__o211a_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09770__A1 _02077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _03714_ _04245_ _03736_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__o21ai_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 genblk2\[10\].wave_shpr.div.b1\[10\] VGND VGND VPWR VPWR net1224 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06584__B2 _01490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1017 genblk2\[1\].wave_shpr.div.b1\[3\] VGND VGND VPWR VPWR net1235 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ _03410_ _03417_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__or2_2
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1028 genblk2\[8\].wave_shpr.div.b1\[9\] VGND VGND VPWR VPWR net1246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 genblk2\[10\].wave_shpr.div.acc\[22\] VGND VGND VPWR VPWR net1257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08672_ _03361_ _03378_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07623_ _02317_ _02328_ _02329_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__a21oi_2
XANTENNA__06887__A2 _01738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10948__A _05051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_18_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout167_A net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07554_ _02223_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__buf_4
XANTENNA__08089__B2 _02527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06505_ _01362_ _01430_ _01196_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_146_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07485_ _02209_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09224_ genblk2\[0\].wave_shpr.div.quo\[5\] _03836_ _03840_ net600 VGND VGND VPWR
+ VPWR _00128_ sky130_fd_sc_hd__a22o_1
XANTENNA__07041__B _01576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06487__A2_N _01411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06436_ genblk1\[1\].osc.clkdiv_C.cnt\[2\] genblk1\[1\].osc.clkdiv_C.cnt\[1\] genblk1\[1\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09155_ genblk2\[0\].wave_shpr.div.acc\[25\] genblk2\[0\].wave_shpr.div.acc\[24\]
+ genblk2\[0\].wave_shpr.div.acc\[26\] _03802_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__or4_2
X_06367_ _01310_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__buf_4
XFILLER_0_17_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08106_ genblk1\[4\].osc.clkdiv_C.cnt\[11\] _01574_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09249__A _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09086_ modein.delay_octave_down_in\[0\] VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__inv_2
X_06298_ genblk1\[0\].osc.clkdiv_C.cnt\[14\] _01256_ _01240_ genblk1\[0\].osc.clkdiv_C.cnt\[13\]
+ _01259_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_142_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08037_ _02364_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__buf_2
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold840 genblk1\[7\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR net1058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 sig_norm.acc\[2\] VGND VGND VPWR VPWR net1069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 genblk1\[10\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR net1080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 genblk2\[1\].wave_shpr.div.i\[1\] VGND VGND VPWR VPWR net1091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 PWM.final_in\[2\] VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold895 genblk2\[7\].wave_shpr.div.i\[1\] VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06425__A2_N _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09988_ genblk2\[3\].wave_shpr.div.b1\[2\] genblk2\[3\].wave_shpr.div.acc\[2\] VGND
+ VGND VPWR VPWR _04384_ sky130_fd_sc_hd__and2b_1
XANTENNA__07772__B1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08939_ sig_norm.quo\[1\] _03631_ _00024_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10659__B1 _04857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11950_ genblk2\[10\].wave_shpr.div.b1\[13\] genblk2\[10\].wave_shpr.div.acc\[13\]
+ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__and2b_1
XANTENNA__07216__B _01442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold546_A genblk2\[1\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10901_ _05034_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11881_ net646 _05684_ _05685_ _05712_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13620_ clknet_leaf_75_clk _00933_ net204 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10832_ genblk2\[6\].wave_shpr.div.acc\[7\] genblk2\[6\].wave_shpr.div.b1\[7\] VGND
+ VGND VPWR VPWR _04976_ sky130_fd_sc_hd__or2b_1
X_13551_ clknet_leaf_100_clk _00866_ net165 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10069__S _04440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10763_ genblk2\[5\].wave_shpr.div.acc\[13\] _04924_ _04907_ VGND VGND VPWR VPWR
+ _04925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12502_ clknet_leaf_106_clk _00064_ net154 VGND VGND VPWR VPWR PWM.final_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09029__B1 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13482_ clknet_leaf_99_clk net347 net168 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10694_ net245 _02183_ _04856_ net503 _04874_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12433_ genblk2\[11\].wave_shpr.div.acc\[21\] _06095_ _06096_ VGND VGND VPWR VPWR
+ _06097_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_63_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06790__B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12364_ _06044_ _05948_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11315_ net852 _05279_ _05283_ _05310_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12295_ _03687_ net425 _03716_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__a21bo_1
X_11246_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09752__A1 _04223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11177_ net1215 genblk2\[7\].wave_shpr.div.quo\[6\] _00019_ VGND VGND VPWR VPWR _05230_
+ sky130_fd_sc_hd__mux2_1
X_10128_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10059_ net1206 _01263_ _04238_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__mux2_1
XANTENNA__06965__B _01344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09807__A2 _04248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07142__A genblk1\[9\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13749_ clknet_leaf_75_clk _01060_ net211 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07270_ _02028_ _02043_ _02044_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__and3_1
XANTENNA__09768__S _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06221_ _01181_ _01182_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__nor2_8
XFILLER_0_155_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06152_ _01121_ _01123_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09069__A _03701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold103 _00957_ VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10050__A1 _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold114 _00715_ VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold125 _01047_ VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _00966_ VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold147 smpl_rt_clkdiv.clkDiv_inst.cnt\[6\] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold158 genblk2\[3\].wave_shpr.div.quo\[16\] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _04200_ _04323_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__xnor2_1
Xhold169 genblk2\[3\].wave_shpr.div.quo\[12\] VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ net520 _04247_ _04250_ net639 _04272_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _04236_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__clkbuf_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06221__A _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ _01795_ _01796_ _01798_ _01818_ _01820_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__o2111a_1
X_08724_ _03429_ _03430_ VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__xnor2_2
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _03263_ _03274_ _03273_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__a21boi_1
XANTENNA__10678__A _04672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12369__S _05982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07606_ net15 net163 _02312_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ _03280_ _03292_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07052__A _01441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07537_ net1111 PWM.final_in\[0\] PWM.start VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07809__B2 _02468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07987__A _02225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07468_ _02147_ _02197_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09207_ _03831_ net674 _03717_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__a21bo_1
XANTENNA__06493__B1 _01418_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06419_ _01362_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__buf_4
X_07399_ _02146_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09138_ _03752_ _03784_ _03785_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__a21o_1
XANTENNA__08234__A1 _02885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12030__A2 _05813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09069_ _03701_ _01221_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__nand2_8
X_11100_ genblk2\[6\].wave_shpr.div.i\[3\] _02187_ _05159_ VGND VGND VPWR VPWR _05162_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07993__B1 _01519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12080_ _05750_ _05745_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__or2b_1
Xhold670 genblk2\[5\].wave_shpr.div.acc\[4\] VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold681 genblk2\[6\].wave_shpr.div.acc\[17\] VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 genblk2\[5\].wave_shpr.div.acc\[2\] VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ net1003 _05086_ _05093_ _05112_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__a22o_1
XANTENNA__10352__S _04637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07745__B1 _01337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06131__A net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12982_ clknet_leaf_125_clk net323 net70 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11933_ _05743_ _05753_ _05754_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__o21ba_1
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12279__S _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11183__S _05042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06785__B _01483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08170__B1 _01507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11864_ net987 _05684_ _05685_ _05700_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12477__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13603_ clknet_leaf_45_clk _00002_ net121 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
X_10815_ genblk2\[5\].wave_shpr.div.i\[1\] genblk2\[5\].wave_shpr.div.i\[0\] genblk2\[5\].wave_shpr.div.i\[2\]
+ genblk2\[5\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__a31o_1
X_11795_ genblk2\[9\].wave_shpr.div.b1\[0\] _05613_ genblk2\[9\].wave_shpr.div.acc\[0\]
+ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__a21o_1
XANTENNA__10804__B1 _04855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13534_ clknet_leaf_81_clk _00849_ net199 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10746_ genblk2\[5\].wave_shpr.div.acc\[10\] _04886_ _04890_ _04911_ VGND VGND VPWR
+ VPWR _00579_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09670__B1 _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13465_ clknet_leaf_75_clk _00782_ net203 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10677_ net294 _04861_ _04862_ net453 _04865_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__a221o_1
XFILLER_0_153_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11212__A _05245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12416_ net878 _06072_ _06073_ _06084_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12021__A2 _05813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13396_ clknet_leaf_117_clk net332 net140 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12347_ genblk2\[11\].wave_shpr.div.b1\[0\] _05982_ genblk2\[11\].wave_shpr.div.acc\[0\]
+ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12309__B1 _03944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08521__A _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12278_ _06000_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13265__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11229_ _05074_ genblk1\[7\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12043__A _04676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07137__A genblk1\[9\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12088__A2 _05844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06770_ genblk1\[4\].osc.clkdiv_C.cnt\[13\] genblk1\[4\].osc.clkdiv_C.cnt\[12\] _01637_
+ genblk1\[4\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06695__B _01323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08440_ _02407_ _02403_ genblk2\[10\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR
+ _03147_ sky130_fd_sc_hd__or3b_1
XFILLER_0_148_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08371_ _02998_ _03000_ _02999_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__o21a_1
XFILLER_0_147_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09498__S _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07322_ genblk1\[11\].osc.clkdiv_C.cnt\[16\] _02085_ VGND VGND VPWR VPWR _02086_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09661__B1 _04045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07600__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07253_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] genblk1\[10\].osc.clkdiv_C.cnt\[0\] genblk1\[10\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06204_ _01166_ _01167_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__and2_1
X_07184_ genblk1\[9\].osc.clkdiv_C.cnt\[9\] _01972_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06135_ net11 _01106_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__xor2_1
XANTENNA__11220__B1 _05250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09527__A _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09825_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__and2_1
XANTENNA__07047__A _01336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09756_ _04226_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10900__S _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06968_ genblk1\[7\].osc.clkdiv_C.cnt\[1\] _01801_ _01803_ VGND VGND VPWR VPWR _01804_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__12079__A2 _05844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08707_ genblk2\[2\].wave_shpr.div.fin_quo\[3\] net25 _03116_ _02224_ VGND VGND VPWR
+ VPWR _03414_ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12099__S _05787_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09687_ genblk2\[2\].wave_shpr.div.acc\[6\] genblk2\[2\].wave_shpr.div.b1\[6\] VGND
+ VGND VPWR VPWR _04167_ sky130_fd_sc_hd__or2b_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06899_ genblk1\[6\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__inv_2
XANTENNA__08152__B1 _01250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _02682_ _02686_ _02685_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__o21ai_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08569_ _03273_ _03274_ _03263_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10600_ genblk2\[5\].wave_shpr.div.fin_quo\[3\] genblk2\[5\].wave_shpr.div.quo\[2\]
+ _00015_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__mux2_1
Xfanout42 net43 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout53 net58 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_2
XFILLER_0_119_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11580_ _05387_ _05495_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout64 net65 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09201__S _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout75 net84 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout86 net88 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10531_ genblk2\[4\].wave_shpr.div.i\[3\] _02176_ _04758_ VGND VGND VPWR VPWR _04761_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout97 net98 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10347__S _04637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13250_ clknet_leaf_2_clk _00573_ net43 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10462_ net1024 _04683_ _04690_ _04711_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06126__A _01097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06218__B1 _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12201_ genblk2\[11\].wave_shpr.div.acc\[3\] genblk2\[11\].wave_shpr.div.b1\[3\]
+ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__or2b_1
XANTENNA__09955__A1 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13181_ clknet_leaf_112_clk _00506_ net68 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10393_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__and2_1
XANTENNA__07966__B1 _01675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12132_ _05774_ _05734_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12063_ genblk2\[10\].wave_shpr.div.quo\[22\] _05812_ _05825_ net334 _05836_ VGND
+ VGND VPWR VPWR _00971_ sky130_fd_sc_hd__a221o_1
XANTENNA__08060__B _01238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06499__C net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11014_ net819 _05086_ _05093_ _05099_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11278__B1 _05250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12965_ clknet_leaf_110_clk _00294_ net130 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11916_ genblk2\[10\].wave_shpr.div.acc\[10\] genblk2\[10\].wave_shpr.div.b1\[10\]
+ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__or2b_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ clknet_leaf_32_clk _00227_ net99 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09900__A _04247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11847_ genblk2\[9\].wave_shpr.div.acc\[12\] _05687_ _05673_ VGND VGND VPWR VPWR
+ _05688_ sky130_fd_sc_hd__mux2_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ net362 _05628_ _05629_ net513 _05638_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13517_ clknet_leaf_77_clk _00834_ net208 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06457__B1 genblk1\[1\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10729_ net863 _04886_ _04890_ _04898_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13448_ clknet_leaf_91_clk _00765_ net147 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08749__A2 _02309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13379_ clknet_leaf_81_clk _00698_ net199 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11753__A1 net526 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07940_ net13 _02364_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__nand2_1
X_07871_ genblk2\[1\].wave_shpr.div.fin_quo\[0\] _02524_ _02307_ genblk2\[1\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__a22o_1
XANTENNA__08382__B1 _01418_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09610_ _04042_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__buf_2
XANTENNA__11816__S _05613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06822_ net1120 _01693_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09541_ net552 _04052_ _04053_ net462 _04061_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__a221o_1
X_06753_ _01599_ _01632_ _01633_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__and3_1
X_09472_ _03701_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__clkbuf_4
X_06684_ _01173_ _01187_ _01188_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__mux2_4
XFILLER_0_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08423_ _03085_ _03123_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__or2_1
XANTENNA__06696__B1 _01574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10956__A _05051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_126_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08354_ _02932_ _02841_ genblk2\[4\].wave_shpr.div.fin_quo\[4\] VGND VGND VPWR VPWR
+ _03061_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08437__A1 _02525_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07305_ _02063_ _02066_ _02067_ _02068_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08285_ _02972_ _02991_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__and2b_1
XFILLER_0_132_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11992__A1 _01855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07236_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] _02001_ _02002_ _02003_ VGND VGND VPWR
+ VPWR _02018_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07167_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01960_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09257__A _03853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06118_ _01088_ _01092_ VGND VGND VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.next_cnt\[5\]
+ sky130_fd_sc_hd__nor2_1
X_07098_ genblk1\[8\].osc.clkdiv_C.cnt\[10\] _01902_ _01905_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[10\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07963__A3 _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout210 net218 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__buf_2
XANTENNA__11726__S _00023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09808_ _04247_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10630__S _04834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout62_A net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09739_ genblk2\[2\].wave_shpr.div.fin_quo\[2\] net1343 _00009_ VGND VGND VPWR VPWR
+ _04217_ sky130_fd_sc_hd__mux2_1
X_12750_ clknet_leaf_46_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[9\] net119 VGND VGND
+ VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_2
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _05561_ _05591_ _05592_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__a21o_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[12\] net82 VGND VGND
+ VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_139_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ genblk2\[8\].wave_shpr.div.acc\[20\] _05533_ _05534_ VGND VGND VPWR VPWR
+ _05535_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11563_ genblk2\[8\].wave_shpr.div.acc\[3\] _05482_ _05417_ VGND VGND VPWR VPWR _05483_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13302_ clknet_leaf_87_clk _00623_ net179 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11983__A1 _03732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10514_ net1144 _04657_ _04655_ _04749_ VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11494_ _05443_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__buf_2
XFILLER_0_107_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13233_ clknet_leaf_15_clk _00556_ net73 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10445_ net998 _04683_ _04690_ _04698_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13164_ clknet_leaf_127_clk net843 net67 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10376_ genblk2\[4\].wave_shpr.div.quo\[5\] _04652_ _04656_ net749 VGND VGND VPWR
+ VPWR _00464_ sky130_fd_sc_hd__a22o_1
X_12115_ _05765_ _05873_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06611__B1 _01171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13095_ clknet_leaf_1_clk _00422_ net41 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12046_ net373 _05823_ _05825_ net521 _05827_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__a221o_1
XANTENNA__11499__B1 _05446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07415__A _02155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12948_ clknet_leaf_125_clk _00277_ net71 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08667__B2 _02362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ clknet_leaf_119_clk _00210_ net139 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07890__A2 _02539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08070_ _02770_ _02771_ _02775_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07021_ genblk1\[7\].osc.clkdiv_C.cnt\[13\] _01842_ _01822_ VGND VGND VPWR VPWR _01844_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11400__A genblk2\[8\].wave_shpr.div.b1\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08972_ _03657_ _03658_ sig_norm.quo\[6\] _01098_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07309__B _01430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07923_ genblk1\[8\].osc.clkdiv_C.cnt\[8\] _01865_ VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__and2_1
Xhold18 _00561_ VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 genblk2\[10\].wave_shpr.div.acc_next\[0\] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08355__B1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout197_A net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07854_ _02518_ _02555_ _02560_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__a21oi_1
X_06805_ genblk1\[5\].osc.clkdiv_C.cnt\[9\] _01362_ _01226_ VGND VGND VPWR VPWR _01677_
+ sky130_fd_sc_hd__and3_1
X_07785_ _02482_ _02488_ _02491_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__o21ba_1
X_09524_ _03853_ genblk1\[1\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__and2_1
X_06736_ genblk1\[4\].osc.clkdiv_C.cnt\[6\] _01616_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__and2_1
XANTENNA__08658__B2 _02592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09540__A _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09455_ _04015_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06667_ _01556_ _01344_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08406_ net25 VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__buf_2
XFILLER_0_143_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09386_ genblk2\[11\].wave_shpr.div.i\[3\] _02212_ _03949_ VGND VGND VPWR VPWR _03952_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_81_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06598_ genblk1\[3\].osc.clkdiv_C.cnt\[16\] _01197_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07060__A genblk1\[8\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08337_ genblk2\[6\].wave_shpr.div.fin_quo\[4\] _02734_ _02737_ _02261_ VGND VGND
+ VPWR VPWR _03044_ sky130_fd_sc_hd__a31o_1
XANTENNA__09428__A_N genblk2\[1\].wave_shpr.div.b1\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08268_ genblk2\[11\].wave_shpr.div.fin_quo\[5\] _02361_ VGND VGND VPWR VPWR _02975_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07219_ _01358_ net37 VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__nand2_2
X_08199_ _02404_ _02410_ _02405_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10230_ genblk2\[3\].wave_shpr.div.acc\[23\] _04417_ VGND VGND VPWR VPWR _04550_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_30_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06404__A genblk1\[1\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10161_ net941 _04486_ _04490_ _04498_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__a22o_1
XANTENNA__07219__B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold576_A genblk2\[3\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10940__A2 _05052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10092_ net814 _04452_ _04456_ net849 VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__a22o_1
XANTENNA__07149__B2 genblk1\[9\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12802_ clknet_leaf_59_clk _00135_ net193 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09846__B1 _04250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10994_ _04982_ _04983_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12445__A2 _03947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12733_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[10\] net115 VGND
+ VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06793__B _01592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11191__S _05042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ clknet_leaf_26_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[13\] net88 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11615_ net802 _05507_ _05445_ _05522_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09074__A1 _01592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12595_ clknet_leaf_11_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[16\] net56 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09596__S _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11546_ net274 _05441_ _05444_ net445 _05470_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11477_ _03704_ net1042 _04233_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13216_ clknet_leaf_6_clk _00539_ net46 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10428_ genblk2\[4\].wave_shpr.div.acc\[1\] _04685_ _04623_ VGND VGND VPWR VPWR _04686_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_880 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13147_ clknet_leaf_121_clk net638 net80 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10359_ genblk2\[5\].wave_shpr.div.b1\[15\] _01365_ _04637_ VGND VGND VPWR VPWR _04648_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07129__B _01801_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13078_ clknet_leaf_125_clk _00405_ net61 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08337__B1 _02261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12029_ net320 _05813_ _05817_ genblk2\[10\].wave_shpr.div.quo\[6\] VGND VGND VPWR
+ VPWR _00956_ sky130_fd_sc_hd__a22o_1
XANTENNA__12051__A _03833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10144__B1 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11892__B1 _03694_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07560__A1 genblk1\[9\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07570_ _02267_ _02273_ _02276_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__a21o_1
X_06521_ _01433_ _01434_ _01435_ _01436_ _01446_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09240_ net495 _03845_ _03847_ net584 _03848_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__a221o_1
X_06452_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] _01387_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09171_ net1218 genblk2\[0\].wave_shpr.div.quo\[6\] _00001_ VGND VGND VPWR VPWR _03812_
+ sky130_fd_sc_hd__mux2_1
X_06383_ _01254_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__clkbuf_8
X_08122_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] _01340_ _01304_ genblk1\[4\].osc.clkdiv_C.cnt\[6\]
+ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08053_ _02756_ _02757_ _02758_ _02759_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout112_A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07004_ _01823_ _01832_ _01833_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_102_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput19 net19 VGND VGND VPWR VPWR sigout sky130_fd_sc_hd__buf_2
XFILLER_0_113_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06224__A _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08576__B1 _02361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07039__B _01487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09535__A _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08955_ net1339 _03644_ _00024_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__mux2_1
X_07906_ genblk1\[8\].osc.clkdiv_C.cnt\[9\] _01859_ _02610_ _02611_ _02612_ VGND VGND
+ VPWR VPWR _02613_ sky130_fd_sc_hd__a2111o_1
X_08886_ sig_norm.b1\[3\] sig_norm.acc\[3\] VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__xnor2_1
X_07837_ _02542_ _02543_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__nor2_1
X_07768_ _02472_ _02473_ _02474_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__or3b_1
XANTENNA__13549__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09507_ _04044_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__clkbuf_4
X_06719_ genblk1\[4\].osc.clkdiv_C.cnt\[1\] genblk1\[4\].osc.clkdiv_C.cnt\[0\] genblk1\[4\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07699_ genblk2\[10\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__inv_2
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09438_ genblk2\[1\].wave_shpr.div.b1\[16\] genblk2\[1\].wave_shpr.div.acc\[16\]
+ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__and2b_1
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09369_ _03937_ _03938_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09056__A1 _01201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11400_ genblk2\[8\].wave_shpr.div.b1\[1\] genblk2\[8\].wave_shpr.div.acc\[1\] VGND
+ VGND VPWR VPWR _05376_ sky130_fd_sc_hd__or2b_1
XFILLER_0_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12380_ _05957_ _05934_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__or2b_1
XFILLER_0_62_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10610__A1 _01189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11331_ _05210_ _05322_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10355__S _04637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11040__A _05051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11262_ _04676_ _01813_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13001_ clknet_leaf_133_clk _00330_ net59 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10213_ _04415_ _04480_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__or2_1
X_11193_ _01865_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__inv_2
X_10144_ net976 _04452_ _04456_ _04485_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08319__B1 _02316_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06788__B _01262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11186__S _05042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10075_ genblk2\[4\].wave_shpr.div.b1\[15\] _01365_ _04440_ VGND VGND VPWR VPWR _04448_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13765_ clknet_leaf_69_clk _01076_ net213 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10977_ genblk2\[6\].wave_shpr.div.quo\[21\] _05062_ _05064_ net567 _05073_ VGND
+ VGND VPWR VPWR _00648_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12716_ clknet_leaf_56_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[11\] net175 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
X_13696_ clknet_leaf_96_clk _01007_ net161 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_127_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12647_ clknet_leaf_9_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[14\] net54 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07058__B1 _01246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12578_ clknet_leaf_29_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[17\] net96 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08524__A _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11529_ net263 _05454_ _05458_ net502 _05461_ VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold307 genblk2\[3\].wave_shpr.div.quo\[11\] VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_40_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold318 genblk2\[10\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 genblk2\[10\].wave_shpr.div.quo\[17\] VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08558__B1 _02223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06584__A2 _01231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _03412_ _03416_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__nand2_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 genblk2\[4\].wave_shpr.div.b1\[7\] VGND VGND VPWR VPWR net1225 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1018 genblk2\[9\].wave_shpr.div.b1\[8\] VGND VGND VPWR VPWR net1236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 genblk2\[2\].wave_shpr.div.b1\[1\] VGND VGND VPWR VPWR net1247 sky130_fd_sc_hd__dlygate4sd3_1
X_08671_ _03362_ _03377_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11824__S _05613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07622_ genblk1\[11\].osc.clkdiv_C.cnt\[7\] _01211_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07603__A _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07553_ _01157_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08089__A2 _02309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06504_ _01224_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07484_ _02206_ _02153_ genblk2\[10\].wave_shpr.div.busy VGND VGND VPWR VPWR _02209_
+ sky130_fd_sc_hd__and3b_2
XANTENNA__06219__A _01174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09223_ net600 _03836_ _03840_ net728 VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__a22o_1
X_06435_ _01377_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09154_ genblk2\[0\].wave_shpr.div.acc\[23\] _03801_ VGND VGND VPWR VPWR _03802_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_146_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06366_ _01308_ _01309_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__nand2_1
X_08105_ _01588_ _01192_ _01208_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__and3_1
X_09085_ _03714_ _03734_ _03736_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06297_ genblk1\[0\].osc.clkdiv_C.cnt\[2\] _01190_ _01258_ genblk1\[0\].osc.clkdiv_C.cnt\[5\]
+ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_130_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06272__A1 _01229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08036_ genblk2\[6\].wave_shpr.div.fin_quo\[7\] _02539_ _02742_ VGND VGND VPWR VPWR
+ _02743_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold830 genblk2\[7\].wave_shpr.div.acc\[19\] VGND VGND VPWR VPWR net1048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold841 genblk2\[9\].wave_shpr.div.acc\[1\] VGND VGND VPWR VPWR net1059 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12345__A1 _03819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold852 genblk2\[7\].wave_shpr.div.acc\[1\] VGND VGND VPWR VPWR net1070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold863 genblk2\[10\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR net1081 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08013__A2 _01367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold874 genblk1\[8\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 PWM.final_in\[1\] VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 genblk2\[8\].wave_shpr.div.acc\[19\] VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09265__A _03853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09987_ _04379_ genblk2\[3\].wave_shpr.div.acc\[1\] _04382_ VGND VGND VPWR VPWR _04383_
+ sky130_fd_sc_hd__a21o_1
X_08938_ sig_norm.quo\[0\] _01098_ _03629_ _03630_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__a22o_1
XANTENNA__07323__A2_N _01334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09513__A2 _04043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08869_ sig_norm.b1\[3\] VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11734__S _00023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10900_ net1288 _01991_ _04848_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__mux2_1
X_11880_ _05609_ _05646_ _05709_ genblk2\[9\].wave_shpr.div.acc\[21\] VGND VGND VPWR
+ VPWR _05712_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_86_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10831_ genblk2\[6\].wave_shpr.div.acc\[8\] genblk2\[6\].wave_shpr.div.b1\[8\] VGND
+ VGND VPWR VPWR _04975_ sky130_fd_sc_hd__or2b_1
XFILLER_0_39_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13550_ clknet_leaf_100_clk _00865_ net170 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10762_ _04805_ _04923_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06129__A net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07827__A2 _02309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06594__A2_N _01500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12501_ clknet_leaf_106_clk _00063_ net153 VGND VGND VPWR VPWR PWM.final_in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13481_ clknet_leaf_100_clk _00798_ net168 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09029__A1 _03694_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10693_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12432_ genblk2\[11\].wave_shpr.div.acc\[21\] genblk2\[11\].wave_shpr.div.acc\[20\]
+ _05978_ net20 VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__or4_1
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12363_ _05949_ _05938_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__or2b_1
XANTENNA__08063__B _01238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11314_ genblk2\[7\].wave_shpr.div.acc\[11\] _05309_ _05300_ VGND VGND VPWR VPWR
+ _05310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12294_ _03732_ net406 _03733_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11245_ net548 _05255_ _05256_ net550 _05262_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__a221o_1
XANTENNA__09201__A1 _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08004__A2 _01519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07212__B1 _01214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11176_ _05229_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__clkbuf_1
X_10127_ net529 _04451_ _04455_ net607 _04474_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10058_ _04438_ VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11311__A2 _05279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08519__A _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07142__B _01514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13748_ clknet_leaf_85_clk net1221 net184 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13679_ clknet_leaf_43_clk net860 net190 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06220_ _01177_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_26_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12024__B1 _05817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06151_ _01107_ _01110_ _01122_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_81_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09069__B _01221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold104 genblk2\[2\].wave_shpr.div.quo\[19\] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold115 genblk2\[3\].wave_shpr.div.i\[4\] VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold126 genblk2\[6\].wave_shpr.div.quo\[10\] VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold137 genblk2\[11\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkbuf_2
Xhold148 genblk2\[1\].wave_shpr.div.acc\[11\] VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ _04201_ _04159_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__or2b_1
XFILLER_0_1_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold159 _00392_ VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09841_ _04269_ genblk1\[2\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__and2_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11550__A2 _05417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ net1298 _01256_ _04039_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06984_ genblk1\[7\].osc.clkdiv_C.cnt\[8\] _01819_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__xnor2_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06221__B _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _02536_ _02586_ VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__and2b_1
XANTENNA__09813__A _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10959__A _05054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08654_ _03320_ _03325_ _03360_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__o21bai_2
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07605_ net17 net18 VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__or2_2
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08585_ _03284_ _03291_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__xnor2_2
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07536_ net279 _02249_ _02251_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07052__B _01226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07467_ genblk2\[8\].wave_shpr.div.busy _02196_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09206_ _02171_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__buf_8
XFILLER_0_151_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06493__A1 _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06418_ _01361_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__buf_4
XANTENNA__08164__A _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07398_ _02091_ _02144_ _02145_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__and3_1
X_09137_ genblk2\[0\].wave_shpr.div.b1\[11\] genblk2\[0\].wave_shpr.div.acc\[11\]
+ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06349_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] _01295_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09068_ _03725_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__buf_8
X_08019_ genblk1\[6\].osc.clkdiv_C.cnt\[8\] _01732_ _02725_ _01753_ VGND VGND VPWR
+ VPWR _02726_ sky130_fd_sc_hd__o2bb2a_1
Xhold660 genblk2\[11\].wave_shpr.div.acc\[17\] VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 genblk2\[0\].wave_shpr.div.acc\[12\] VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08611__B _02223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold682 genblk2\[6\].wave_shpr.div.acc\[11\] VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ genblk2\[6\].wave_shpr.div.acc\[9\] _05111_ _05105_ VGND VGND VPWR VPWR _05112_
+ sky130_fd_sc_hd__mux2_1
Xhold693 _00571_ VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06412__A _01226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07745__A1 genblk1\[1\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07745__B2 genblk1\[1\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12981_ clknet_leaf_124_clk _00310_ net75 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09498__A1 _01327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11932_ genblk2\[10\].wave_shpr.div.b1\[4\] genblk2\[10\].wave_shpr.div.acc\[4\]
+ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__and2b_1
XFILLER_0_87_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ genblk2\[9\].wave_shpr.div.acc\[16\] _05699_ _05673_ VGND VGND VPWR VPWR
+ _05700_ sky130_fd_sc_hd__mux2_1
XANTENNA__09869__S _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10814_ _04855_ _04959_ _04960_ _04858_ net1154 VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__a32o_1
X_13602_ clknet_leaf_77_clk _00917_ net209 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11794_ _05646_ _05573_ genblk2\[9\].wave_shpr.div.b1\[0\] VGND VGND VPWR VPWR _05647_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10745_ net772 _04910_ _04907_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__mux2_1
X_13533_ clknet_leaf_81_clk _00848_ net199 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09670__A1 _04045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13464_ clknet_leaf_83_clk _00781_ net203 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10676_ _04672_ genblk1\[5\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12415_ genblk2\[11\].wave_shpr.div.acc\[16\] _06083_ _06055_ VGND VGND VPWR VPWR
+ _06084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13395_ clknet_leaf_116_clk _00714_ net140 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10109__A _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12346_ genblk2\[11\].wave_shpr.div.b1\[0\] genblk2\[11\].wave_shpr.div.acc\[0\]
+ _05982_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__nand3_1
XFILLER_0_23_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12309__B2 net355 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12277_ net1274 _02001_ _05994_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__mux2_1
XANTENNA__12324__A _03689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07418__A _02160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11228_ net302 _05251_ _05248_ net492 _05252_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11159_ genblk2\[7\].wave_shpr.div.acc\[22\] _05218_ VGND VGND VPWR VPWR _05219_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06976__B _01811_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08370_ _03054_ _03075_ _03076_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__or3_2
XFILLER_0_58_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07321_ genblk1\[11\].osc.clkdiv_C.cnt\[15\] _01359_ VGND VGND VPWR VPWR _02085_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06475__A1 genblk1\[1\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07600__B net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07252_ genblk1\[10\].osc.clkdiv_C.cnt\[2\] genblk1\[10\].osc.clkdiv_C.cnt\[1\] genblk1\[10\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06203_ PWM.counter\[6\] _01164_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__or2_1
XANTENNA__08415__C _02365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07183_ genblk1\[9\].osc.clkdiv_C.cnt\[9\] _01972_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06227__A1 _01174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06134_ _01104_ _01105_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__nand2_1
XANTENNA__09808__A _04247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10453__S _04704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09824_ net315 _04257_ _04259_ net480 _04262_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__a221o_1
XANTENNA__07047__B _01223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09755_ genblk2\[3\].wave_shpr.div.b1\[1\] _04225_ _04039_ VGND VGND VPWR VPWR _04226_
+ sky130_fd_sc_hd__mux2_1
X_06967_ genblk1\[7\].osc.clkdiv_C.cnt\[7\] _01574_ _01802_ genblk1\[7\].osc.clkdiv_C.cnt\[6\]
+ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__a22o_1
X_08706_ _03113_ _03116_ genblk2\[2\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR
+ _03413_ sky130_fd_sc_hd__a21oi_1
X_09686_ genblk2\[2\].wave_shpr.div.acc\[7\] genblk2\[2\].wave_shpr.div.b1\[7\] VGND
+ VGND VPWR VPWR _04166_ sky130_fd_sc_hd__or2b_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08159__A _01489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06898_ genblk1\[6\].osc.clkdiv_C.cnt\[6\] _01367_ _01750_ genblk1\[6\].osc.clkdiv_C.cnt\[7\]
+ _01751_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__a221o_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _02592_ _03342_ _03343_ _02636_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__a211o_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _03263_ _03273_ _03274_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__nand3_1
XFILLER_0_49_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07519_ _01163_ PWM.final_sample_in\[4\] _02233_ _02238_ VGND VGND VPWR VPWR _02239_
+ sky130_fd_sc_hd__a22o_1
Xfanout43 net44 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08499_ _02547_ _02586_ _02588_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout54 net58 VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10628__S _04834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout65 net68 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout76 net84 VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_4
X_10530_ _00012_ _04758_ net1160 VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__a21oi_1
Xfanout87 net88 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07663__B1 _01241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout98 net127 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_2
XFILLER_0_134_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10461_ genblk2\[4\].wave_shpr.div.acc\[9\] _04710_ _04704_ VGND VGND VPWR VPWR _04711_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06218__A1 _01174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12200_ genblk2\[11\].wave_shpr.div.acc\[4\] genblk2\[11\].wave_shpr.div.b1\[4\]
+ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__or2b_1
XFILLER_0_33_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13180_ clknet_leaf_130_clk _00505_ net68 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10392_ net637 _04661_ _04663_ genblk2\[4\].wave_shpr.div.quo\[12\] _04664_ VGND
+ VGND VPWR VPWR _00472_ sky130_fd_sc_hd__a221o_1
X_12131_ net945 _05876_ _05883_ _05886_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12062_ _05835_ genblk1\[10\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR _05836_
+ sky130_fd_sc_hd__and2_1
Xhold490 genblk2\[5\].wave_shpr.div.b1\[6\] VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06142__A net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11013_ genblk2\[6\].wave_shpr.div.acc\[5\] _05098_ _05023_ VGND VGND VPWR VPWR _05099_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12964_ clknet_leaf_111_clk _00293_ net130 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11915_ genblk2\[10\].wave_shpr.div.acc\[11\] genblk2\[10\].wave_shpr.div.b1\[11\]
+ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__or2b_1
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ clknet_leaf_32_clk _00226_ net99 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11846_ _05595_ _05686_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__xnor2_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _04676_ _02268_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06457__A1 genblk1\[1\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10728_ genblk2\[5\].wave_shpr.div.acc\[5\] _04897_ _04821_ VGND VGND VPWR VPWR _04898_
+ sky130_fd_sc_hd__mux2_1
X_13516_ clknet_leaf_78_clk _00833_ net208 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10659_ net745 _04853_ _04857_ net882 VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__a22o_1
X_13447_ clknet_leaf_90_clk _00764_ net144 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09946__A2 _04253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13378_ clknet_leaf_81_clk _00697_ net205 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10781__B _04880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11753__A2 _05623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12329_ net509 _06014_ _06015_ net510 _06022_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__a221o_1
XANTENNA__07148__A genblk1\[9\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07870_ _02221_ _02510_ _02576_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__o21bai_1
X_06821_ net27 VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11269__A1 _05248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09540_ _04058_ _02444_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__nor2_1
X_06752_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01627_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__or2_1
X_09471_ _01418_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06683_ _01566_ _01567_ _01569_ _01572_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__or4b_1
XFILLER_0_92_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08422_ _03011_ _03128_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__and2b_1
XFILLER_0_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10492__A2 _04715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08353_ _03058_ _03059_ _02798_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout142_A net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07304_ genblk1\[11\].osc.clkdiv_C.cnt\[5\] _02064_ _01925_ genblk1\[11\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_117_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08284_ _02984_ _02989_ _02990_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07235_ genblk1\[10\].osc.clkdiv_C.cnt\[16\] _02016_ VGND VGND VPWR VPWR _02017_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11787__B genblk1\[9\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07166_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01960_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06117_ net380 _01087_ net407 VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__a21oi_1
X_07097_ _01887_ _01904_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08161__B _01498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout200 net210 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_2
Xfanout211 net212 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10911__S _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09807_ genblk2\[2\].wave_shpr.div.quo\[8\] _04248_ _04252_ net275 VGND VGND VPWR
+ VPWR _00299_ sky130_fd_sc_hd__a22o_1
X_07999_ _01200_ genblk1\[6\].osc.clkdiv_C.cnt\[15\] _01361_ _02704_ _02705_ VGND
+ VGND VPWR VPWR _02706_ sky130_fd_sc_hd__o311a_1
XANTENNA__07581__C1 genblk1\[9\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09738_ _04216_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout55_A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _04151_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ genblk2\[9\].wave_shpr.div.b1\[10\] genblk2\[9\].wave_shpr.div.acc\[10\]
+ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__and2b_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[11\] net82 VGND VGND
+ VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _05410_ _05416_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__and2b_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11562_ _05379_ _05481_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06137__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10513_ genblk2\[4\].wave_shpr.div.acc\[23\] _04620_ _04748_ VGND VGND VPWR VPWR
+ _04749_ sky130_fd_sc_hd__a21o_1
X_13301_ clknet_leaf_84_clk _00622_ net202 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11493_ _02152_ genblk2\[8\].wave_shpr.div.busy _02196_ VGND VGND VPWR VPWR _05443_
+ sky130_fd_sc_hd__and3_1
X_13232_ clknet_leaf_15_clk net501 net73 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10444_ genblk2\[4\].wave_shpr.div.acc\[5\] _04697_ _04623_ VGND VGND VPWR VPWR _04698_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13163_ clknet_leaf_114_clk _00488_ net67 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10375_ genblk2\[4\].wave_shpr.div.quo\[4\] _04652_ _04656_ net732 VGND VGND VPWR
+ VPWR _00463_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10943__B1 _05056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12114_ _05766_ _05738_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__or2b_1
XFILLER_0_20_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13094_ clknet_leaf_1_clk _00421_ net38 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12045_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__and2_1
XANTENNA__12160__A2 _05818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06600__A _01241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10122__A _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12947_ clknet_leaf_125_clk _00276_ net69 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ clknet_leaf_119_clk net685 net143 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07431__A _02152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11829_ genblk2\[9\].wave_shpr.div.acc\[8\] _05672_ _05673_ VGND VGND VPWR VPWR _05674_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07627__B1 _01256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07020_ net1189 _01841_ _01843_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_141_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08971_ _03656_ _03523_ _01098_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__a21o_1
X_07922_ _02624_ _02626_ _02627_ _02628_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__o211a_1
Xhold19 genblk2\[8\].wave_shpr.div.quo\[14\] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07606__A net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07853_ _02558_ _02559_ _02424_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06510__A _01349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06804_ genblk1\[5\].osc.clkdiv_C.cnt\[15\] _01362_ genblk1\[5\].osc.clkdiv_C.cnt\[17\]
+ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__a21o_1
X_07784_ genblk1\[0\].osc.clkdiv_C.cnt\[5\] _02486_ _02489_ _02490_ VGND VGND VPWR
+ VPWR _02491_ sky130_fd_sc_hd__o31ai_1
XANTENNA__12439__B1 _03944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08107__A1 _01192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09821__A _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06735_ _01619_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[5\] sky130_fd_sc_hd__clkbuf_1
X_09523_ net610 _04048_ _04045_ net517 _04050_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__a221o_1
XANTENNA__08658__A2 _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09454_ genblk2\[1\].wave_shpr.div.fin_quo\[3\] genblk2\[1\].wave_shpr.div.quo\[2\]
+ _00007_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__mux2_1
X_06666_ _01230_ _01221_ _01223_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__a21o_4
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08405_ genblk1\[2\].osc.clkdiv_C.cnt\[16\] _01578_ _03111_ genblk1\[2\].osc.clkdiv_C.cnt\[17\]
+ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09385_ _00004_ _03949_ net1163 VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06597_ genblk1\[3\].osc.clkdiv_C.cnt\[16\] _01197_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08336_ _02734_ _02737_ genblk2\[6\].wave_shpr.div.fin_quo\[4\] VGND VGND VPWR VPWR
+ _03043_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08267_ genblk2\[11\].wave_shpr.div.fin_quo\[4\] net33 _02350_ _02354_ _02222_ VGND
+ VGND VPWR VPWR _02974_ sky130_fd_sc_hd__a41o_1
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07218_ genblk1\[10\].osc.clkdiv_C.cnt\[14\] _01246_ _01442_ genblk1\[10\].osc.clkdiv_C.cnt\[13\]
+ _01999_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__a221o_1
XANTENNA__09268__A _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08198_ _02902_ _02903_ _02904_ _02360_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07149_ genblk1\[9\].osc.clkdiv_C.cnt\[12\] _01799_ _01947_ genblk1\[9\].osc.clkdiv_C.cnt\[1\]
+ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_132_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06404__B _01327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10160_ genblk2\[3\].wave_shpr.div.acc\[5\] _04497_ _04420_ VGND VGND VPWR VPWR _04498_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10091_ genblk2\[3\].wave_shpr.div.quo\[4\] _04452_ _04456_ net779 VGND VGND VPWR
+ VPWR _00379_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12801_ clknet_leaf_59_clk net570 net193 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10993_ genblk2\[6\].wave_shpr.div.acc\[1\] _05022_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__or2_1
XANTENNA__11102__B1 _03855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[9\] net115 VGND VGND
+ VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07857__B1 _02316_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold903_A genblk2\[1\].wave_shpr.div.b1\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ clknet_leaf_26_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[12\] net88 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09877__S _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11614_ genblk2\[8\].wave_shpr.div.acc\[15\] _05521_ _05493_ VGND VGND VPWR VPWR
+ _05522_ sky130_fd_sc_hd__mux2_1
X_12594_ clknet_leaf_12_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[15\] net52 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_53_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11545_ _05464_ genblk1\[8\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_131_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_131_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_67_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13760__RESET_B net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11476_ _05435_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10427_ _04585_ _04684_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__nor2_1
X_13215_ clknet_leaf_6_clk _00538_ net48 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_892 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10358_ _03704_ net800 _04647_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__a21o_1
X_13146_ clknet_leaf_121_clk _00471_ net81 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13077_ clknet_leaf_125_clk _00404_ net62 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _04573_ _04599_ _04600_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_125_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12332__A _03833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12028_ genblk2\[10\].wave_shpr.div.quo\[6\] _05813_ _05817_ net555 VGND VGND VPWR
+ VPWR _00955_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06984__B _01819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06520_ _01438_ _01443_ _01444_ _01445_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__or4_1
XFILLER_0_87_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07312__A2 _01210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06451_ _01373_ _01387_ _01388_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__09787__S _04238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09170_ _03811_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06382_ _01229_ _01325_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__nand2_4
X_08121_ genblk1\[4\].osc.clkdiv_C.cnt\[3\] _01439_ _02827_ VGND VGND VPWR VPWR _02828_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_122_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_122_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_114_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08052_ _01489_ genblk1\[5\].osc.clkdiv_C.cnt\[9\] net37 _01667_ genblk1\[5\].osc.clkdiv_C.cnt\[10\]
+ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__a32o_1
XFILLER_0_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07003_ genblk1\[7\].osc.clkdiv_C.cnt\[6\] _01830_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__nor2_1
XANTENNA__08576__A1 _02525_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09816__A _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10461__S _04704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08954_ sig_norm.quo\[3\] _03643_ _02248_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__mux2_1
XANTENNA__09525__B1 _04045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07905_ genblk1\[8\].osc.clkdiv_C.cnt\[10\] _01870_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__xnor2_1
X_08885_ sig_norm.acc\[10\] _03590_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07055__B _01430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07836_ genblk2\[0\].wave_shpr.div.fin_quo\[4\] _02510_ _02512_ _02261_ VGND VGND
+ VPWR VPWR _02543_ sky130_fd_sc_hd__a31o_1
X_07767_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] _01309_ _01208_ genblk1\[0\].osc.clkdiv_C.cnt\[14\]
+ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__o22a_1
X_09506_ _02170_ genblk2\[1\].wave_shpr.div.busy _02157_ VGND VGND VPWR VPWR _04044_
+ sky130_fd_sc_hd__and3_1
X_06718_ _01605_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__inv_2
X_07698_ genblk2\[10\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09437_ _03956_ _03999_ _04000_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__a21oi_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06649_ genblk1\[3\].osc.clkdiv_C.cnt\[12\] _01543_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09368_ genblk2\[0\].wave_shpr.div.acc\[25\] _03802_ genblk2\[0\].wave_shpr.div.acc\[24\]
+ genblk2\[0\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__or4b_1
XFILLER_0_93_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08319_ genblk2\[9\].wave_shpr.div.fin_quo\[3\] _02303_ _02263_ _02316_ VGND VGND
+ VPWR VPWR _03026_ sky130_fd_sc_hd__a31o_1
XFILLER_0_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_113_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_113_clk sky130_fd_sc_hd__clkbuf_16
X_09299_ _03777_ _03756_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__or2b_1
XFILLER_0_90_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11321__A _05249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11330_ _05211_ _05166_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__or2b_1
XFILLER_0_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11261_ net534 _05245_ _05249_ genblk2\[7\].wave_shpr.div.quo\[23\] _05270_ VGND
+ VGND VPWR VPWR _00735_ sky130_fd_sc_hd__a221o_1
XANTENNA__08016__B1 _01739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10212_ net657 _04518_ _04522_ _04537_ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__a22o_1
X_13000_ clknet_leaf_132_clk _00329_ net63 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07568__A2_N _01349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11192_ _05235_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__clkbuf_1
X_10143_ genblk2\[3\].wave_shpr.div.acc\[1\] _04484_ _04420_ VGND VGND VPWR VPWR _04485_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09516__B1 _04047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10074_ _04447_ VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13764_ clknet_leaf_69_clk _01075_ net214 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10976_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12715_ clknet_leaf_54_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[10\] net175 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_85_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13695_ clknet_leaf_45_clk _01006_ net188 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12646_ clknet_leaf_24_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[13\] net92 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07058__A1 genblk1\[8\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_104_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_104_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_5_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07058__B2 genblk1\[8\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12577_ clknet_leaf_21_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[16\] net95 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11231__A _05074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11528_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold308 genblk2\[9\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__buf_1
XANTENNA__08007__B1 _01735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold319 genblk2\[1\].wave_shpr.div.quo\[12\] VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__dlygate4sd3_1
X_11459_ _05426_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08558__A1 genblk2\[8\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ clknet_leaf_3_clk _00454_ net46 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07156__A genblk1\[9\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1008 genblk2\[10\].wave_shpr.div.acc\[25\] VGND VGND VPWR VPWR net1226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1019 genblk1\[3\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR net1237 sky130_fd_sc_hd__dlygate4sd3_1
X_08670_ _03366_ _03376_ VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09371__A _02170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07621_ genblk1\[11\].osc.clkdiv_C.cnt\[6\] _01430_ _02326_ _02327_ VGND VGND VPWR
+ VPWR _02328_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_49_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07552_ _02259_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07603__B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06503_ genblk1\[2\].osc.clkdiv_C.cnt\[12\] _01411_ _01415_ _01419_ _01428_ VGND
+ VGND VPWR VPWR _01429_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_76_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12290__A1 _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07483_ _02208_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09222_ genblk2\[0\].wave_shpr.div.quo\[3\] _03836_ _03840_ net558 VGND VGND VPWR
+ VPWR _00126_ sky130_fd_sc_hd__a22o_1
X_06434_ _01374_ _01375_ _01376_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09153_ genblk2\[0\].wave_shpr.div.acc\[22\] genblk2\[0\].wave_shpr.div.acc\[21\]
+ genblk2\[0\].wave_shpr.div.acc\[20\] _03800_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__or4_1
XANTENNA__07049__A1 genblk1\[8\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06365_ _01171_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08104_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01323_ _01592_ genblk1\[4\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09084_ _03735_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__buf_8
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06235__A _01196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06296_ _01238_ _01257_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__or2_2
XFILLER_0_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08035_ _02221_ _02733_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__nor2_2
XFILLER_0_130_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold820 genblk2\[5\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR net1038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold831 genblk2\[0\].wave_shpr.div.acc\[8\] VGND VGND VPWR VPWR net1049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12345__A2 net1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold842 genblk2\[9\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR net1060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold853 genblk2\[4\].wave_shpr.div.b1\[0\] VGND VGND VPWR VPWR net1071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 genblk2\[0\].wave_shpr.div.acc\[25\] VGND VGND VPWR VPWR net1082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 genblk2\[6\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold886 genblk1\[6\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR net1104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold897 genblk1\[5\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ genblk2\[3\].wave_shpr.div.b1\[0\] _04380_ _04381_ VGND VGND VPWR VPWR _04382_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__07772__A2 _01190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08937_ _01098_ _03550_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__nor2_1
XANTENNA__06980__B1 _01574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10659__A2 _04853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08868_ _01156_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07819_ _02525_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08799_ _03500_ _03504_ _03427_ _03505_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__o211a_1
XANTENNA__11316__A _05245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10830_ genblk2\[6\].wave_shpr.div.acc\[9\] genblk2\[6\].wave_shpr.div.b1\[9\] VGND
+ VGND VPWR VPWR _04974_ sky130_fd_sc_hd__or2b_1
XFILLER_0_39_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10761_ _04806_ _04767_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__or2b_1
XANTENNA__12281__A1 _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06129__B net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12500_ clknet_leaf_102_clk net429 net156 VGND VGND VPWR VPWR sig_norm.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13480_ clknet_leaf_99_clk _00797_ net168 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10692_ genblk2\[5\].wave_shpr.div.quo\[20\] _04861_ _04862_ net233 _04873_ VGND
+ VGND VPWR VPWR _00563_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12431_ genblk2\[11\].wave_shpr.div.acc\[20\] _05978_ net20 VGND VGND VPWR VPWR _06095_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12362_ net985 _06039_ _06040_ _06043_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__a22o_1
XANTENNA__06145__A _01114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06799__B1 _01304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08063__C net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11313_ _05202_ _05308_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12293_ _06008_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11244_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08360__A _02885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10347__A1 _01658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07212__A1 _01308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11175_ genblk2\[7\].wave_shpr.div.fin_quo\[6\] net754 _00019_ VGND VGND VPWR VPWR
+ _05229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07763__A2 _02468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10126_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__and2_1
XANTENNA__06971__B1 _01805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10057_ net1225 _01329_ _04238_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07920__C1 _01441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11226__A _05245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13747_ clknet_leaf_51_clk net413 net111 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10959_ _05054_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__buf_2
XFILLER_0_70_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13678_ clknet_leaf_42_clk _00991_ net125 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12629_ clknet_leaf_120_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[14\] net82 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06150_ _01103_ _01111_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold105 _00311_ VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 genblk2\[10\].wave_shpr.div.quo\[21\] VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold127 _00638_ VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _01042_ VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _00245_ VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10338__A1 _03831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ genblk2\[2\].wave_shpr.div.quo\[22\] _04247_ _04259_ net261 _04271_ VGND
+ VGND VPWR VPWR _00313_ sky130_fd_sc_hd__a221o_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08400__B1 _01591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _04235_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__clkbuf_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06983_ _01436_ _01334_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__nand2_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _02588_ _02546_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__nor2_1
XANTENNA__07506__A2 _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08653_ _03313_ _03326_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07604_ genblk2\[9\].wave_shpr.div.fin_quo\[7\] _02309_ _02310_ VGND VGND VPWR VPWR
+ _02311_ sky130_fd_sc_hd__a21o_1
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _03289_ _03290_ _02419_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07535_ net279 _02249_ _01099_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12263__A1 _01263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07466_ _02195_ genblk2\[8\].wave_shpr.div.i\[1\] genblk2\[8\].wave_shpr.div.i\[0\]
+ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__or3b_1
XFILLER_0_147_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09205_ _03704_ net759 _03728_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06417_ _01360_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07397_ genblk1\[11\].osc.clkdiv_C.cnt\[16\] _02143_ VGND VGND VPWR VPWR _02145_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09136_ _03753_ _03782_ _03783_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06348_ _01269_ _01294_ _01295_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_60_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09067_ _02155_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__buf_2
X_06279_ _01237_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__buf_4
XANTENNA__06607__A2_N _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07993__A2 _01484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08018_ _01739_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold650 genblk2\[10\].wave_shpr.div.acc\[4\] VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 genblk2\[5\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 genblk2\[3\].wave_shpr.div.acc\[7\] VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 genblk2\[4\].wave_shpr.div.acc\[13\] VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 genblk2\[9\].wave_shpr.div.acc\[15\] VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06412__B _01355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout85_A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07745__A2 _01344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09969_ genblk2\[3\].wave_shpr.div.acc\[13\] genblk2\[3\].wave_shpr.div.b1\[13\]
+ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__or2b_1
X_12980_ clknet_leaf_14_clk _00309_ net72 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11931_ _05744_ _05751_ _05752_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__a21oi_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08170__A2 _01508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11862_ _05698_ _05603_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13601_ clknet_leaf_77_clk _00916_ net209 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10813_ genblk2\[5\].wave_shpr.div.i\[1\] genblk2\[5\].wave_shpr.div.i\[0\] genblk2\[5\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__nand3_1
X_11793_ _05610_ _05611_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13532_ clknet_leaf_97_clk _00023_ net166 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10804__A2 _04858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10744_ _04797_ _04909_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12006__A1 _01494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13463_ clknet_leaf_83_clk _00780_ net203 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10675_ net453 _04861_ _04862_ net500 _04864_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__a221o_1
X_12414_ _05926_ _05972_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13394_ clknet_leaf_116_clk net564 net145 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12345_ _03819_ net1220 _00004_ genblk2\[11\].wave_shpr.div.acc\[0\] _06030_ VGND
+ VGND VPWR VPWR _01059_ sky130_fd_sc_hd__o221a_1
XANTENNA__08630__B1 _02261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12309__A2 _03947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08090__A net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12276_ _05999_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09186__A1 _03704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11227_ _05074_ genblk1\[7\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06322__B genblk1\[0\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11158_ genblk2\[7\].wave_shpr.div.acc\[21\] genblk2\[7\].wave_shpr.div.acc\[20\]
+ genblk2\[7\].wave_shpr.div.acc\[19\] _05217_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__or4_1
X_10109_ _04268_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__clkbuf_2
X_11089_ net1043 _05057_ _05055_ _05154_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__a22o_1
XANTENNA__12340__A _03833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07434__A _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08449__B1 _02316_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12245__A1 _05982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07320_ genblk1\[11\].osc.clkdiv_C.cnt\[4\] _01513_ _02076_ _02079_ _02083_ VGND
+ VGND VPWR VPWR _02084_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_45_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09661__A2 _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07121__B1 _01855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07251_ _02031_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[1\] sky130_fd_sc_hd__clkbuf_1
X_06202_ PWM.counter\[6\] _01164_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07182_ _01953_ _01972_ _01973_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_42_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06133_ net8 net9 VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11220__A2 _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07609__A _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06513__A _01213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12181__B1 _05818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07727__A2 _02433_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09823_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__and2_1
XANTENNA__06593__A2_N _01498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09754_ _01436_ _01925_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__nand2_2
X_06966_ _01192_ _01245_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__nand2_1
X_08705_ _03361_ _03378_ _03411_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__a21o_1
X_09685_ genblk2\[2\].wave_shpr.div.acc\[8\] genblk2\[2\].wave_shpr.div.b1\[8\] VGND
+ VGND VPWR VPWR _04165_ sky130_fd_sc_hd__or2b_1
XFILLER_0_96_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06897_ genblk1\[6\].osc.clkdiv_C.cnt\[6\] _01367_ _01750_ genblk1\[6\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__o22ai_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08152__A2 _01500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _02216_ _02552_ genblk2\[8\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR
+ _03343_ sky130_fd_sc_hd__and3_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ _02946_ _03272_ _03268_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07998__B _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10909__S _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10247__B1 _04457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07518_ _02232_ PWM.final_sample_in\[3\] PWM.final_sample_in\[2\] _02234_ _02237_
+ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout44 net85 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
X_08498_ _03077_ _03203_ _03175_ _03202_ VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__a211oi_1
XANTENNA__09652__A2 _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout55 net58 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_147_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout66 net68 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout77 net84 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07663__A1 _01360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07449_ _02180_ _02153_ genblk2\[5\].wave_shpr.div.busy VGND VGND VPWR VPWR _02184_
+ sky130_fd_sc_hd__and3b_1
Xfanout88 net91 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_4
Xfanout99 net101 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10460_ _04599_ _04709_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11747__B1 _05624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09119_ _03761_ genblk2\[0\].wave_shpr.div.acc\[2\] _03766_ VGND VGND VPWR VPWR _03767_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10391_ _04058_ _01570_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12130_ genblk2\[10\].wave_shpr.div.acc\[13\] _05885_ _05865_ VGND VGND VPWR VPWR
+ _05886_ sky130_fd_sc_hd__mux2_1
XANTENNA__07966__A2 _01214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11739__A1_N _01099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12061_ _02155_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold480 genblk2\[4\].wave_shpr.div.quo\[23\] VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 genblk2\[8\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12172__B1 _05816_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11012_ _05097_ _04991_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12963_ clknet_leaf_111_clk _00292_ net130 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11278__A2 _05279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_84_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_16
X_11914_ genblk2\[10\].wave_shpr.div.acc\[12\] genblk2\[10\].wave_shpr.div.b1\[12\]
+ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__or2b_1
XFILLER_0_59_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ clknet_leaf_32_clk net427 net99 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _05596_ _05559_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__or2b_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10238__B1 _04454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ net513 _05628_ _05629_ net530 _05637_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__a221o_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13515_ clknet_leaf_78_clk _00832_ net206 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10727_ _04896_ _04789_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09909__A _04250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13446_ clknet_leaf_99_clk _00021_ net166 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12667__RESET_B net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10658_ genblk2\[5\].wave_shpr.div.quo\[2\] _04853_ _04857_ net879 VGND VGND VPWR
+ VPWR _00545_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13377_ clknet_leaf_81_clk _00696_ net199 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10589_ genblk2\[5\].wave_shpr.div.acc\[21\] genblk2\[5\].wave_shpr.div.acc\[20\]
+ genblk2\[5\].wave_shpr.div.acc\[19\] _04816_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__or4_1
XANTENNA__07429__A _02155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12328_ _03689_ genblk1\[11\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__and2_1
XANTENNA__09159__A1 genblk2\[0\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12259_ genblk2\[11\].wave_shpr.div.fin_quo\[7\] net1341 _00005_ VGND VGND VPWR VPWR
+ _05990_ sky130_fd_sc_hd__mux2_1
XANTENNA__08959__S _02248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08382__A2 _02336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06820_ _01656_ _01657_ _01664_ _01691_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__nor4_1
XANTENNA__12070__A _05815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07590__B1 _01923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07164__A genblk1\[9\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06751_ _01631_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_75_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09470_ _04022_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__clkbuf_1
X_06682_ genblk1\[4\].osc.clkdiv_C.cnt\[4\] _01439_ _01340_ genblk1\[4\].osc.clkdiv_C.cnt\[8\]
+ _01571_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__o221a_1
X_08421_ _03079_ _03127_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__or2b_1
XANTENNA__06696__A2 _01326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08352_ genblk2\[5\].wave_shpr.div.fin_quo\[5\] _02521_ _02791_ VGND VGND VPWR VPWR
+ _03059_ sky130_fd_sc_hd__a21o_1
XANTENNA__09095__A0 _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07303_ genblk1\[11\].osc.clkdiv_C.cnt\[13\] _01256_ _01595_ genblk1\[11\].osc.clkdiv_C.cnt\[6\]
+ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08283_ _02366_ _02976_ _02983_ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout135_A net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09819__A _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07234_ genblk1\[10\].osc.clkdiv_C.cnt\[15\] _01359_ VGND VGND VPWR VPWR _02016_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07165_ _01953_ _01960_ _01961_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__09538__B genblk1\[1\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06116_ net380 _01087_ VGND VGND VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.next_cnt\[4\]
+ sky130_fd_sc_hd__xor2_1
X_07096_ genblk1\[8\].osc.clkdiv_C.cnt\[10\] genblk1\[8\].osc.clkdiv_C.cnt\[9\] _01900_
+ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout201 net210 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_4
Xfanout212 net213 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10704__A1 _03819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09806_ net275 _04248_ _04252_ net449 VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07998_ genblk1\[6\].osc.clkdiv_C.cnt\[14\] _01361_ VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__nand2_1
XANTENNA__07581__B1 _01171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09737_ genblk2\[2\].wave_shpr.div.fin_quo\[1\] net1348 _00009_ VGND VGND VPWR VPWR
+ _04216_ sky130_fd_sc_hd__mux2_1
X_06949_ net1356 _01787_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_66_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08125__A2 _01870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09668_ genblk2\[1\].wave_shpr.div.i\[1\] genblk2\[1\].wave_shpr.div.i\[0\] genblk2\[1\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__and3_1
XANTENNA__09207__B1_N _03717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08530__C1 net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout48_A net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07802__A _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08619_ _03320_ _03325_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__xor2_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10639__S _04834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09599_ _03987_ _04100_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__xnor2_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ genblk2\[8\].wave_shpr.div.acc\[18\] genblk2\[8\].wave_shpr.div.acc\[19\]
+ _05529_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06418__A _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11561_ _05380_ _05372_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__or2b_1
XANTENNA__06137__B net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13300_ clknet_leaf_83_clk _00621_ net199 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10512_ genblk2\[4\].wave_shpr.div.acc\[25\] genblk2\[4\].wave_shpr.div.acc\[24\]
+ genblk2\[4\].wave_shpr.div.acc\[26\] _04621_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__o31a_1
XFILLER_0_80_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11492_ _05441_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13231_ clknet_leaf_11_clk _00554_ net73 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10443_ _04696_ _04591_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13162_ clknet_leaf_115_clk _00487_ net67 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10374_ net732 _04652_ _04656_ net793 VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__a22o_1
XANTENNA__10009__A_N genblk2\[3\].wave_shpr.div.b1\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_871 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12113_ net951 _05844_ _05850_ _05872_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__a22o_1
XANTENNA__11994__A _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13093_ clknet_leaf_139_clk _00420_ net39 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12044_ net521 _05823_ _05825_ net583 _05826_ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__a221o_1
XANTENNA__10403__A _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06600__B _01432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_57_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_16
X_12946_ clknet_leaf_125_clk _00275_ net69 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12877_ clknet_leaf_119_clk _00208_ net141 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11234__A _05249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11828_ _05612_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__buf_4
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11759_ net481 _03696_ _03694_ net557 _05627_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13429_ clknet_leaf_83_clk _00748_ net201 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08052__A1 _01489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06602__A2 _01484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08970_ _03656_ _03523_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__nor2_1
XANTENNA__08412__C_N net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07921_ genblk1\[8\].osc.clkdiv_C.cnt\[7\] _01430_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__or2_1
XANTENNA__10698__B1 _04856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12004__S _05802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07606__B net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07852_ genblk2\[1\].wave_shpr.div.fin_quo\[3\] _02309_ _02469_ VGND VGND VPWR VPWR
+ _02559_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07563__B1 _01801_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06803_ _01674_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__buf_4
XFILLER_0_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 pb[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
X_07783_ _01200_ genblk1\[0\].osc.clkdiv_C.cnt\[6\] genblk1\[0\].osc.clkdiv_C.cnt\[7\]
+ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_48_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08107__A2 _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09522_ _03853_ genblk1\[1\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__and2_1
X_06734_ _01600_ _01617_ _01618_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07315__B1 _02077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09453_ _04014_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__clkbuf_1
X_06665_ net436 _01554_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08404_ _01201_ genblk1\[2\].osc.clkdiv_C.cnt\[16\] _01362_ _03109_ _03110_ VGND
+ VGND VPWR VPWR _03111_ sky130_fd_sc_hd__o311a_1
XFILLER_0_19_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09384_ _03944_ _03948_ _03950_ _03947_ net741 VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__a32o_1
XFILLER_0_52_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06596_ genblk1\[3\].osc.clkdiv_C.cnt\[17\] _01493_ _01495_ _01503_ VGND VGND VPWR
+ VPWR _01504_ sky130_fd_sc_hd__or4b_1
XANTENNA__06238__A _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08335_ _02604_ _03034_ _03040_ _02648_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__a22o_1
XANTENNA__10983__A _05074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08266_ _02349_ _02351_ _02354_ genblk2\[11\].wave_shpr.div.fin_quo\[4\] VGND VGND
+ VPWR VPWR _02973_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07217_ _01995_ _01996_ _01997_ _01342_ _01998_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09268__B genblk1\[0\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08197_ genblk2\[11\].wave_shpr.div.fin_quo\[6\] _02361_ VGND VGND VPWR VPWR _02904_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07148_ genblk1\[9\].osc.clkdiv_C.cnt\[1\] _01947_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07079_ _01887_ _01892_ _01893_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__10922__S _05042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10090_ genblk2\[3\].wave_shpr.div.quo\[3\] _04452_ _04456_ net737 VGND VGND VPWR
+ VPWR _00378_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12800_ clknet_leaf_59_clk _00133_ net192 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10992_ _05081_ _05082_ net1122 _05052_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_96_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09846__A2 _04247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12731_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[8\] net115 VGND VGND
+ VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09059__A0 _01229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12941__RESET_B net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12662_ clknet_leaf_25_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[11\] net87 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _05403_ _05520_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12593_ clknet_leaf_13_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[14\] net70 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11544_ net445 _05441_ _05458_ net505 _05469_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11475_ net1236 net34 _05433_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13214_ clknet_leaf_6_clk _00537_ net48 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10426_ genblk2\[4\].wave_shpr.div.b1\[0\] _04583_ _04584_ VGND VGND VPWR VPWR _04684_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_111_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10916__A1 _01797_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13145_ clknet_leaf_121_clk net603 net81 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10357_ _03708_ _01441_ _01367_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__and3_4
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07707__A _02316_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13076_ clknet_leaf_136_clk _00403_ net62 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ genblk2\[4\].wave_shpr.div.b1\[9\] genblk2\[4\].wave_shpr.div.acc\[9\] VGND
+ VGND VPWR VPWR _04600_ sky130_fd_sc_hd__and2b_1
X_12027_ net555 _05813_ _05817_ net723 VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__a22o_1
XANTENNA__11229__A _05074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10133__A _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10144__A2 _04452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11892__A2 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12929_ clknet_leaf_123_clk _00008_ net76 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11644__A2 _05448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06450_ genblk1\[1\].osc.clkdiv_C.cnt\[6\] _01385_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__nor2_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06381_ _01324_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08120_ _01224_ _01249_ genblk1\[4\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _02827_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_154_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08051_ genblk1\[5\].osc.clkdiv_C.cnt\[10\] _01667_ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07002_ genblk1\[7\].osc.clkdiv_C.cnt\[6\] _01830_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__and2_1
XANTENNA__09222__B1 _03840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08953_ _03559_ _03642_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__xnor2_1
X_07904_ genblk1\[8\].osc.clkdiv_C.cnt\[11\] _01869_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__nor2_1
X_08884_ sig_norm.acc\[9\] _03589_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07835_ _02510_ _02512_ genblk2\[0\].wave_shpr.div.fin_quo\[4\] VGND VGND VPWR VPWR
+ _02542_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10978__A _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07766_ genblk1\[0\].osc.clkdiv_C.cnt\[13\] _01255_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__and2_1
XANTENNA__09043__S _03708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09505_ _04042_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__buf_4
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06717_ genblk1\[4\].osc.clkdiv_C.cnt\[2\] genblk1\[4\].osc.clkdiv_C.cnt\[1\] genblk1\[4\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__and3_1
X_07697_ _02403_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__buf_2
XFILLER_0_63_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08167__B _01231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09436_ genblk2\[1\].wave_shpr.div.b1\[15\] genblk2\[1\].wave_shpr.div.acc\[15\]
+ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__and2b_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07071__B genblk1\[8\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06648_ _01486_ _01542_ _01544_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__a21oi_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09367_ genblk2\[0\].wave_shpr.div.acc\[24\] _03802_ genblk2\[0\].wave_shpr.div.acc\[25\]
+ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06579_ _01172_ _01182_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__nand2_4
XANTENNA__12225__A_N genblk2\[11\].wave_shpr.div.b1\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08318_ _02303_ _02263_ genblk2\[9\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR
+ _03025_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09298_ net964 _03870_ _03877_ _03886_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10071__A1 _01595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08249_ genblk2\[8\].wave_shpr.div.fin_quo\[6\] _02309_ _02636_ VGND VGND VPWR VPWR
+ _02956_ sky130_fd_sc_hd__a21o_1
XANTENNA__06814__A2 _01242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12348__B1 _03947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11260_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__and2_1
XANTENNA__13558__RESET_B net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10211_ genblk2\[3\].wave_shpr.div.acc\[17\] _04536_ _04507_ VGND VGND VPWR VPWR
+ _04537_ sky130_fd_sc_hd__mux2_1
XANTENNA__09764__A1 _01794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11191_ net1280 _01556_ _05042_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10142_ _04382_ _04483_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11049__A _05054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09516__A1 net292 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10073_ net1262 _04242_ _04440_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__mux2_1
X_13763_ clknet_leaf_69_clk _01074_ net214 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10975_ genblk2\[6\].wave_shpr.div.quo\[20\] _05062_ _05064_ net313 _05072_ VGND
+ VGND VPWR VPWR _00647_ sky130_fd_sc_hd__a221o_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12714_ clknet_leaf_54_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[9\] net175 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_2
X_13694_ clknet_leaf_45_clk _01005_ net122 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12645_ clknet_leaf_24_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[12\] net92 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09189__A _03701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07058__A2 _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08255__B2 _02539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12576_ clknet_leaf_29_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[15\] net95 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__06606__A _01234_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10062__A1 _01240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11527_ net502 _05454_ _05458_ net611 _05460_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12339__B1 _03941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold309 genblk2\[7\].wave_shpr.div.quo\[20\] VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11458_ genblk2\[9\].wave_shpr.div.b1\[0\] _02064_ _05237_ VGND VGND VPWR VPWR _05426_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09755__A1 _04225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08558__A2 genblk2\[8\].wave_shpr.div.fin_quo\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10409_ genblk2\[4\].wave_shpr.div.quo\[21\] _04661_ _04663_ net626 _04673_ VGND
+ VGND VPWR VPWR _00480_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11389_ genblk2\[8\].wave_shpr.div.acc\[10\] genblk2\[8\].wave_shpr.div.b1\[10\]
+ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ clknet_leaf_3_clk _00453_ net46 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ clknet_leaf_24_clk _00386_ net92 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07156__B genblk1\[9\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1009 genblk2\[4\].wave_shpr.div.b1\[17\] VGND VGND VPWR VPWR net1227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07620_ genblk1\[11\].osc.clkdiv_C.cnt\[6\] _01430_ _01595_ genblk1\[11\].osc.clkdiv_C.cnt\[5\]
+ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07551_ net1142 net1128 PWM.start VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06502_ genblk1\[2\].osc.clkdiv_C.cnt\[11\] _01420_ _01421_ _01422_ _01427_ VGND
+ VGND VPWR VPWR _01428_ sky130_fd_sc_hd__o221a_1
XFILLER_0_124_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07482_ _02147_ _02207_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09221_ net558 _03836_ _03840_ net655 VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06433_ genblk1\[1\].osc.clkdiv_C.cnt\[1\] genblk1\[1\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09152_ genblk2\[0\].wave_shpr.div.acc\[19\] _03799_ VGND VGND VPWR VPWR _03800_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_146_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06364_ _01178_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__inv_4
XANTENNA__06254__A2_N _01215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06516__A _01200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08103_ genblk1\[4\].osc.clkdiv_C.cnt\[11\] _01574_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06295_ _01188_ _01187_ _01173_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__o21ba_1
X_09083_ _02170_ _01201_ _01363_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__or3_4
XANTENNA_fanout215_A net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08034_ _02739_ _02740_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__and2b_1
XFILLER_0_141_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09827__A _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold810 _00043_ VGND VGND VPWR VPWR net1028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold821 genblk2\[9\].wave_shpr.div.i\[1\] VGND VGND VPWR VPWR net1039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 genblk2\[0\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR net1050 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11568__S _05417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold843 genblk2\[5\].wave_shpr.div.acc\[11\] VGND VGND VPWR VPWR net1061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09546__B genblk1\[1\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold854 genblk1\[5\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR net1072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 sig_norm.quo\[0\] VGND VGND VPWR VPWR net1083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 genblk2\[2\].wave_shpr.div.acc\[25\] VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 genblk1\[5\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR net1105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 genblk2\[8\].wave_shpr.div.acc\[1\] VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09985_ genblk2\[3\].wave_shpr.div.b1\[1\] genblk2\[3\].wave_shpr.div.acc\[1\] VGND
+ VGND VPWR VPWR _04381_ sky130_fd_sc_hd__xor2_1
XANTENNA__06251__A _01174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08936_ _03529_ _03547_ _03549_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__a21o_1
X_08867_ net1131 _02260_ _03573_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__a21o_1
XANTENNA__08182__B1 _02224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07818_ _02524_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__clkbuf_4
X_08798_ _03425_ _03426_ _03423_ _03424_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_79_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07082__A genblk1\[8\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07749_ _02426_ _02454_ _02428_ _02451_ _02455_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__a221o_1
X_10760_ _04856_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07810__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09419_ _03965_ genblk2\[1\].wave_shpr.div.acc\[6\] _03982_ VGND VGND VPWR VPWR _03983_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10691_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_124_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12430_ net931 _06072_ _06073_ _06094_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12361_ genblk2\[11\].wave_shpr.div.acc\[3\] _06042_ _05982_ VGND VGND VPWR VPWR
+ _06043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11792__A1 _03819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11312_ _05203_ _05170_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__or2b_1
XFILLER_0_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12292_ net1270 _01327_ _05994_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_139_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11243_ net550 _05255_ _05256_ net613 _05261_ VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11174_ _05228_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__clkbuf_1
X_10125_ genblk2\[3\].wave_shpr.div.quo\[21\] _04461_ _04462_ net545 _04473_ VGND
+ VGND VPWR VPWR _00396_ sky130_fd_sc_hd__a221o_1
XANTENNA__09472__A _03701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10056_ _04437_ VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11507__A _05441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07920__B1 genblk1\[8\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10807__A0 _04856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13746_ clknet_leaf_51_clk net435 net110 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10958_ genblk2\[6\].wave_shpr.div.quo\[12\] _05062_ _05055_ net623 _05063_ VGND
+ VGND VPWR VPWR _00639_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13677_ clknet_leaf_42_clk _00990_ net125 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10889_ _05028_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12338__A _03833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12628_ clknet_leaf_18_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[13\] net81 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08228__B2 _02362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12024__A2 _05813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11232__B1 _05248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12559_ clknet_leaf_56_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[16\] net181 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_102_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold106 genblk2\[5\].wave_shpr.div.quo\[24\] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 _00971_ VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 genblk2\[8\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 genblk2\[10\].wave_shpr.div.quo\[15\] VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07167__A genblk1\[9\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ genblk2\[3\].wave_shpr.div.b1\[7\] _02077_ _04039_ VGND VGND VPWR VPWR _04235_
+ sky130_fd_sc_hd__mux2_1
X_06982_ _01800_ _01804_ _01807_ _01817_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__and4_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _03408_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__inv_2
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07506__A3 _02224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08652_ _03334_ _03335_ _03357_ _03358_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__a211oi_4
X_07603_ _02221_ net32 VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__nor2_2
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08583_ genblk2\[10\].wave_shpr.div.fin_quo\[2\] _02308_ _02416_ VGND VGND VPWR VPWR
+ _03290_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout165_A net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07534_ _01151_ _02245_ _02250_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07465_ genblk2\[8\].wave_shpr.div.i\[2\] genblk2\[8\].wave_shpr.div.i\[3\] genblk2\[8\].wave_shpr.div.i\[4\]
+ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_9_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09204_ _03830_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06416_ _01359_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__buf_4
XFILLER_0_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07396_ genblk1\[11\].osc.clkdiv_C.cnt\[16\] _02143_ VGND VGND VPWR VPWR _02144_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07690__A2 _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08164__C _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09135_ genblk2\[0\].wave_shpr.div.b1\[10\] genblk2\[0\].wave_shpr.div.acc\[10\]
+ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__and2b_1
XANTENNA__11223__B1 _05250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06347_ genblk1\[0\].osc.clkdiv_C.cnt\[14\] genblk1\[0\].osc.clkdiv_C.cnt\[13\] _01291_
+ VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09557__A _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09066_ _03724_ VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06278_ _01238_ _01239_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__nor2_8
X_08017_ _02720_ _02722_ _02723_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__o21ai_1
Xhold640 genblk2\[10\].wave_shpr.div.acc\[13\] VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 _00979_ VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 _00545_ VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07077__A genblk1\[8\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold673 genblk2\[4\].wave_shpr.div.acc\[8\] VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 genblk2\[5\].wave_shpr.div.acc\[14\] VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 genblk2\[0\].wave_shpr.div.acc\[14\] VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06402__B1 _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09968_ genblk2\[3\].wave_shpr.div.acc\[14\] genblk2\[3\].wave_shpr.div.b1\[14\]
+ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__or2b_1
X_08919_ sig_norm.acc\[6\] _03614_ net612 VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__o21ai_1
X_09899_ net857 _04282_ _04289_ _04314_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__a22o_1
XANTENNA__08155__B1 _01494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11930_ genblk2\[10\].wave_shpr.div.b1\[3\] genblk2\[10\].wave_shpr.div.acc\[3\]
+ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__and2b_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _05604_ _05555_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13600_ clknet_leaf_76_clk _00915_ net208 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10812_ genblk2\[5\].wave_shpr.div.i\[1\] genblk2\[5\].wave_shpr.div.i\[0\] genblk2\[5\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__a21o_1
XANTENNA__09655__B1 _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11792_ _03819_ genblk1\[9\].osc.clkdiv_C.cnt\[17\] _00022_ net1209 _05645_ VGND
+ VGND VPWR VPWR _00891_ sky130_fd_sc_hd__o221a_1
XANTENNA__08636__A _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13531_ clknet_leaf_84_clk _00022_ net202 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10743_ _04798_ _04771_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13462_ clknet_leaf_83_clk _00779_ net203 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10674_ _04672_ genblk1\[5\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12413_ net1125 _06072_ _06073_ _06082_ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13393_ clknet_leaf_118_clk _00712_ net139 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12344_ genblk2\[11\].wave_shpr.div.acc_next\[0\] _03941_ VGND VGND VPWR VPWR _06030_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_51_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12275_ genblk2\[1\].wave_shpr.div.b1\[6\] _01311_ _05994_ VGND VGND VPWR VPWR _05999_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08090__B _02364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11226_ _05245_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11157_ genblk2\[7\].wave_shpr.div.acc\[18\] _05216_ VGND VGND VPWR VPWR _05217_
+ sky130_fd_sc_hd__or2_1
X_10108_ genblk2\[3\].wave_shpr.div.quo\[13\] _04461_ _04462_ net387 _04464_ VGND
+ VGND VPWR VPWR _00388_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11088_ _05152_ _05153_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__nand2_1
XANTENNA__11237__A _05074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10039_ genblk2\[3\].wave_shpr.div.fin_quo\[6\] net1346 _04422_ VGND VGND VPWR VPWR
+ _04429_ sky130_fd_sc_hd__mux2_1
XANTENNA__08449__A1 genblk2\[8\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07450__A _02184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13729_ clknet_leaf_74_clk _01040_ net212 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11185__A2_N _01432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07121__A1 genblk1\[9\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07121__B2 genblk1\[9\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07250_ _02028_ _02029_ _02030_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__and3_1
XFILLER_0_144_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06201_ _01164_ net811 VGND VGND VPWR VPWR PWM.next_counter\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_0_155_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07181_ genblk1\[9\].osc.clkdiv_C.cnt\[7\] _01967_ genblk1\[9\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06132_ net8 net9 VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08385__B1 _01418_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12181__A1 _05816_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09822_ genblk2\[2\].wave_shpr.div.quo\[14\] _04257_ _04259_ net457 _04261_ VGND
+ VGND VPWR VPWR _00305_ sky130_fd_sc_hd__a221o_1
X_09753_ _04224_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__clkbuf_1
X_06965_ _01213_ _01344_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__nand2_2
X_08704_ _03362_ _03377_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__and2b_1
X_09684_ genblk2\[2\].wave_shpr.div.acc\[9\] genblk2\[2\].wave_shpr.div.b1\[9\] VGND
+ VGND VPWR VPWR _04164_ sky130_fd_sc_hd__or2b_1
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06896_ _01342_ _01439_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__nand2_2
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ genblk2\[8\].wave_shpr.div.fin_quo\[2\] _03341_ VGND VGND VPWR VPWR _03342_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _02946_ _03268_ _03272_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__or3_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10247__A1 _04454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11444__A0 genblk2\[8\].wave_shpr.div.fin_quo\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07517_ _02234_ PWM.final_sample_in\[2\] PWM.final_sample_in\[1\] _02235_ _02236_
+ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08497_ _03175_ _03202_ _03077_ _03203_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout45 net47 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_4
Xfanout56 net58 VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11995__A1 _02805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout67 net68 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07448_ _02183_ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__inv_2
Xfanout78 net79 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07663__A2 _01224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout89 net90 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07379_ genblk1\[11\].osc.clkdiv_C.cnt\[12\] _02130_ VGND VGND VPWR VPWR _02131_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_72_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09118_ _03764_ _03765_ _03762_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10390_ _04654_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__buf_2
XFILLER_0_115_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09049_ _03713_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12060_ net334 _05823_ _05825_ net383 _05834_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__a221o_1
Xhold470 genblk2\[0\].wave_shpr.div.acc\[19\] VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 genblk2\[8\].wave_shpr.div.acc\[2\] VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 genblk2\[3\].wave_shpr.div.acc\[22\] VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ _04992_ _04978_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__or2b_1
X_12962_ clknet_leaf_130_clk _00291_ net65 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11913_ genblk2\[10\].wave_shpr.div.acc\[13\] genblk2\[10\].wave_shpr.div.b1\[13\]
+ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__or2b_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ clknet_leaf_28_clk _00224_ net91 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _03693_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__clkbuf_4
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _04676_ _01930_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__nor2_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11986__A1 _01811_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _04790_ _04775_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13514_ clknet_leaf_78_clk _00831_ net207 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13445_ clknet_leaf_81_clk _00020_ net199 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
X_10657_ net879 _04853_ _04857_ net1056 VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13376_ clknet_leaf_96_clk _00695_ net167 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10588_ genblk2\[5\].wave_shpr.div.acc\[18\] _04815_ VGND VGND VPWR VPWR _04816_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09800__B1 _04252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06614__B1 _01484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12327_ net510 _06014_ _06015_ net571 _06021_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12258_ _05989_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12636__RESET_B net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11209_ _02171_ net1191 VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__and2_1
X_12189_ genblk2\[11\].wave_shpr.div.acc\[15\] genblk2\[11\].wave_shpr.div.b1\[15\]
+ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__or2b_1
XANTENNA__12351__A _05982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06750_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01627_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__and2_1
X_06681_ genblk1\[4\].osc.clkdiv_C.cnt\[15\] _01362_ _01248_ _01570_ VGND VGND VPWR
+ VPWR _01571_ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08420_ _03079_ _03125_ _03126_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08351_ genblk2\[5\].wave_shpr.div.fin_quo\[4\] _03056_ _03057_ VGND VGND VPWR VPWR
+ _03058_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09095__A1 _01556_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07302_ genblk1\[11\].osc.clkdiv_C.cnt\[13\] _01256_ _02064_ genblk1\[11\].osc.clkdiv_C.cnt\[5\]
+ _02065_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08282_ _02987_ _02988_ _02314_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07233_ genblk1\[10\].osc.clkdiv_C.cnt\[16\] _01363_ genblk1\[10\].osc.clkdiv_C.cnt\[15\]
+ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_6_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07164_ genblk1\[9\].osc.clkdiv_C.cnt\[3\] _01958_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06115_ _01087_ _01091_ VGND VGND VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.next_cnt\[3\]
+ sky130_fd_sc_hd__nor2_1
X_07095_ _01887_ _01902_ _01903_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09835__A _02147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout202 net204 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_4
Xfanout213 net217 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_4
X_09805_ net449 _04248_ _04252_ net716 VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__a22o_1
X_07997_ genblk1\[6\].osc.clkdiv_C.cnt\[14\] _01360_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09736_ _04215_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__clkbuf_1
X_06948_ genblk1\[6\].osc.clkdiv_C.cnt\[15\] genblk1\[6\].osc.clkdiv_C.cnt\[14\] _01783_
+ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09667_ genblk2\[1\].wave_shpr.div.i\[1\] genblk2\[1\].wave_shpr.div.i\[0\] genblk2\[1\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__a21o_1
X_06879_ genblk1\[6\].osc.clkdiv_C.cnt\[4\] _01730_ _01732_ genblk1\[6\].osc.clkdiv_C.cnt\[9\]
+ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08530__B1 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08618_ _03323_ _03324_ _02846_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__o21ai_2
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07802__B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09598_ _03988_ _03962_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__or2b_1
XANTENNA__08186__A net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13165__RESET_B net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08549_ _03253_ _03255_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__xnor2_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11968__A1 genblk2\[10\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11560_ net872 _05447_ _05446_ _05480_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10511_ net787 _04657_ _04722_ _04747_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11491_ _02198_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13230_ clknet_leaf_11_clk net311 net73 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10442_ _04592_ _04577_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__or2b_1
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13161_ clknet_leaf_122_clk _00486_ net79 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10373_ genblk2\[4\].wave_shpr.div.quo\[2\] _04652_ _04656_ net464 VGND VGND VPWR
+ VPWR _00461_ sky130_fd_sc_hd__a22o_1
XANTENNA__08061__A2 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12112_ genblk2\[10\].wave_shpr.div.acc\[9\] _05871_ _05865_ VGND VGND VPWR VPWR
+ _05872_ sky130_fd_sc_hd__mux2_1
XANTENNA__10943__A2 _05052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13092_ clknet_leaf_137_clk _00419_ net39 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12043_ _04676_ _01993_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11656__B1 _05448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12945_ clknet_leaf_13_clk _00274_ net69 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07324__B2 _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08096__A _01174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12876_ clknet_leaf_49_clk _00207_ net113 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10224__A2_N _04480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11827_ _05587_ _05671_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__xnor2_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11758_ _05464_ genblk1\[9\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__and2_1
XANTENNA__07627__A2 _01209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10709_ genblk2\[5\].wave_shpr.div.b1\[0\] _04781_ _04782_ VGND VGND VPWR VPWR _04883_
+ sky130_fd_sc_hd__and3_1
X_11689_ _05569_ _05580_ _05567_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13428_ clknet_leaf_82_clk net798 net201 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13359_ clknet_leaf_91_clk _00018_ net143 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07920_ genblk1\[8\].osc.clkdiv_C.cnt\[7\] _01430_ genblk1\[8\].osc.clkdiv_C.cnt\[6\]
+ _01441_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__a211o_1
X_07851_ _02556_ _02557_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__or2_1
XANTENNA__11895__A0 _03838_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06802_ _01238_ net36 VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__nor2_1
X_07782_ genblk1\[0\].osc.clkdiv_C.cnt\[4\] _01241_ _02483_ VGND VGND VPWR VPWR _02489_
+ sky130_fd_sc_hd__o21a_1
Xinput2 pb[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12439__A2 _03947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09521_ net517 _04048_ _04045_ net460 _04049_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__a221o_1
X_06733_ genblk1\[4\].osc.clkdiv_C.cnt\[4\] genblk1\[4\].osc.clkdiv_C.cnt\[3\] _01605_
+ genblk1\[4\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__a31o_1
XANTENNA__07903__A genblk1\[8\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09452_ genblk2\[1\].wave_shpr.div.fin_quo\[2\] net1312 _00007_ VGND VGND VPWR VPWR
+ _04014_ sky130_fd_sc_hd__mux2_1
X_06664_ _01555_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[16\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__07622__B _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08403_ _03103_ _03105_ _03106_ _03107_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09383_ _03949_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06595_ genblk1\[3\].osc.clkdiv_C.cnt\[15\] _01363_ _01499_ _01501_ _01502_ VGND
+ VGND VPWR VPWR _01503_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08334_ _02604_ _02648_ _03034_ _03040_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__nand4_2
XFILLER_0_129_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08265_ _02971_ _02914_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07216_ genblk1\[10\].osc.clkdiv_C.cnt\[13\] _01442_ VGND VGND VPWR VPWR _01998_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08196_ genblk2\[11\].wave_shpr.div.fin_quo\[5\] net33 _02350_ _02355_ _02222_ VGND
+ VGND VPWR VPWR _02903_ sky130_fd_sc_hd__a41o_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07147_ _01241_ _01946_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10386__B1 _04655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07078_ genblk1\[8\].osc.clkdiv_C.cnt\[3\] _01890_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07085__A genblk1\[8\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout60_A net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09719_ genblk2\[2\].wave_shpr.div.b1\[13\] genblk2\[2\].wave_shpr.div.acc\[13\]
+ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__and2b_1
X_10991_ genblk2\[6\].wave_shpr.div.b1\[0\] genblk2\[6\].wave_shpr.div.acc\[0\] _05023_
+ _05079_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__a31o_1
XANTENNA__07306__A1 _01223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12730_ clknet_leaf_39_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[7\] net115 VGND VGND
+ VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ clknet_leaf_26_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[10\] net88 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _05404_ _05360_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ clknet_leaf_13_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[13\] net70 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_108_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11543_ _05464_ genblk1\[8\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12981__RESET_B net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11474_ _05434_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13213_ clknet_leaf_7_clk _00536_ net49 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10425_ _04651_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13144_ clknet_leaf_121_clk net673 net81 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07242__B1 _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10356_ _04646_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ clknet_leaf_2_clk _00402_ net42 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10287_ _04574_ _04597_ _04598_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__a21o_1
XANTENNA__10129__B1 _04455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10414__A _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12026_ genblk2\[10\].wave_shpr.div.quo\[4\] _05813_ _05817_ net682 VGND VGND VPWR
+ VPWR _00953_ sky130_fd_sc_hd__a22o_1
XANTENNA__08019__A2_N _01732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12928_ clknet_leaf_35_clk _00259_ net118 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ clknet_leaf_132_clk _00190_ net64 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06380_ _01178_ _01176_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__and2_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08050_ genblk1\[5\].osc.clkdiv_C.cnt\[11\] _01355_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07001_ _01823_ _01830_ _01831_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06802__A _01238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08952_ _03564_ _03563_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__or2b_1
XANTENNA__07228__A2_N _01235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07903_ genblk1\[8\].osc.clkdiv_C.cnt\[11\] _01360_ _02011_ VGND VGND VPWR VPWR _02610_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09525__A2 _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08883_ sig_norm.acc\[8\] _03588_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout195_A net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07834_ _02537_ _02538_ _02540_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__o21a_1
X_07765_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] _01309_ _01208_ genblk1\[0\].osc.clkdiv_C.cnt\[14\]
+ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06716_ _01604_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[1\] sky130_fd_sc_hd__clkbuf_1
X_09504_ _02159_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07696_ _02398_ _02402_ genblk1\[10\].osc.clkdiv_C.cnt\[16\] genblk1\[10\].osc.clkdiv_C.cnt\[17\]
+ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__a211o_4
XANTENNA__06249__A _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09435_ _03957_ _03997_ _03998_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__a21o_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06647_ _01522_ _01543_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09366_ net1082 _03841_ _03839_ _03936_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06578_ genblk1\[3\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08317_ _03018_ _03023_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09297_ genblk2\[0\].wave_shpr.div.acc\[6\] _03885_ _03804_ VGND VGND VPWR VPWR _03886_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08248_ _02953_ _02954_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_887 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12348__A1 _03944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08179_ genblk2\[3\].wave_shpr.div.fin_quo\[0\] genblk2\[3\].wave_shpr.div.fin_quo\[1\]
+ genblk2\[3\].wave_shpr.div.fin_quo\[2\] genblk2\[3\].wave_shpr.div.fin_quo\[3\]
+ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__or4_1
XFILLER_0_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10210_ _04412_ _04535_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__xnor2_1
X_11190_ _03831_ net768 _04241_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_101_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10141_ genblk2\[3\].wave_shpr.div.b1\[0\] _04380_ _04381_ VGND VGND VPWR VPWR _04483_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_30_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13598__RESET_B net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold574_A genblk2\[6\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09516__A2 _04043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10072_ _04446_ VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13180__RESET_B net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13762_ clknet_leaf_69_clk net994 net214 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10974_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__and2_1
XANTENNA__06159__A _01114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12713_ clknet_leaf_55_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[8\] net175 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_1
X_13693_ clknet_leaf_45_clk _01004_ net122 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12036__B1 _05816_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12644_ clknet_leaf_10_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[11\] net57 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12575_ clknet_leaf_29_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[14\] net95 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08093__B _01360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11004__S _05023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11526_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11457_ _05425_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10408_ _04672_ genblk1\[4\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07718__A _01360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11388_ genblk2\[8\].wave_shpr.div.acc\[11\] genblk2\[8\].wave_shpr.div.b1\[11\]
+ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__or2b_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10339_ _03732_ net708 _03717_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__o21a_1
X_13127_ clknet_leaf_3_clk _00452_ net46 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13268__RESET_B net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ clknet_leaf_24_clk _00385_ net92 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12009_ _05809_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08268__B _02361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07550_ _02258_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06501_ genblk1\[2\].osc.clkdiv_C.cnt\[15\] _01424_ _01425_ _01426_ VGND VGND VPWR
+ VPWR _01427_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07481_ genblk2\[10\].wave_shpr.div.busy _02206_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09220_ net655 _03836_ _03840_ net804 VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__a22o_1
X_06432_ genblk1\[1\].osc.clkdiv_C.cnt\[1\] genblk1\[1\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01375_ sky130_fd_sc_hd__or2_1
XANTENNA__12027__B1 _05817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09151_ genblk2\[0\].wave_shpr.div.acc\[18\] _03798_ VGND VGND VPWR VPWR _03799_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_134_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06363_ genblk1\[1\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_8_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08102_ genblk1\[4\].osc.clkdiv_C.cnt\[11\] _01574_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__and2_1
XANTENNA__06516__B _01441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09082_ net702 VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06294_ _01255_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08033_ _02699_ _02734_ _02738_ genblk2\[6\].wave_shpr.div.fin_quo\[6\] VGND VGND
+ VPWR VPWR _02740_ sky130_fd_sc_hd__a31o_1
Xhold800 genblk2\[8\].wave_shpr.div.acc\[21\] VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 genblk2\[7\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold822 _00072_ VGND VGND VPWR VPWR net1040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 genblk1\[2\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR net1051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 genblk2\[5\].wave_shpr.div.acc\[1\] VGND VGND VPWR VPWR net1062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 sig_norm.b1\[2\] VGND VGND VPWR VPWR net1073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 genblk2\[0\].wave_shpr.div.b1\[11\] VGND VGND VPWR VPWR net1084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 genblk1\[3\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold888 genblk2\[0\].wave_shpr.div.i\[1\] VGND VGND VPWR VPWR net1106 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ genblk2\[3\].wave_shpr.div.acc\[0\] VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__inv_2
Xhold899 genblk2\[5\].wave_shpr.div.i\[1\] VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09843__A _04269_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08935_ net1083 _02260_ _03596_ _03574_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__a22o_1
XANTENNA__06980__A2 _01578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08866_ net428 _02248_ _00024_ _03572_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07817_ net17 net18 VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__and2b_2
X_08797_ _03501_ _03502_ _03500_ _03503_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_98_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07082__B genblk1\[8\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07748_ genblk1\[1\].osc.clkdiv_C.cnt\[16\] _01576_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07679_ _01489_ genblk1\[10\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR _02386_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07810__B net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09418_ _03965_ genblk2\[1\].wave_shpr.div.acc\[6\] _03981_ VGND VGND VPWR VPWR _03982_
+ sky130_fd_sc_hd__o21a_1
X_10690_ net233 _04861_ _04862_ net507 _04872_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__a221o_1
XANTENNA__08194__A net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09349_ _03924_ _03925_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12360_ _05946_ _06041_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06799__A2 _01210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11311_ net894 _05279_ _05283_ _05307_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11792__A2 genblk1\[9\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12291_ _06007_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__clkbuf_1
X_11242_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11544__A2 _05441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11173_ genblk2\[7\].wave_shpr.div.fin_quo\[5\] genblk2\[7\].wave_shpr.div.quo\[4\]
+ _00019_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10124_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__and2_1
X_10055_ net1178 _04436_ _04238_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__mux2_1
XANTENNA__09370__B1 _03839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07920__A1 genblk1\[8\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10807__A1 _02183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13745_ clknet_leaf_51_clk net439 net110 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10957_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11523__A _05444_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07684__A0 _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06487__B2 _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11480__A1 _01732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13676_ clknet_leaf_42_clk _00989_ net124 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10888_ genblk2\[6\].wave_shpr.div.fin_quo\[4\] net1319 _00017_ VGND VGND VPWR VPWR
+ _05028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12627_ clknet_leaf_120_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[12\] net81 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12558_ clknet_leaf_55_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[15\] net176 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_112_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11509_ _04268_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12489_ clknet_leaf_107_clk _00051_ net151 VGND VGND VPWR VPWR sig_norm.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold107 _00568_ VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 genblk2\[2\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold129 _00799_ VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07448__A _02183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07739__A1 genblk1\[1\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07739__B2 genblk1\[1\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08978__S _02248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08400__A2 _02425_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _01809_ _01810_ _01812_ _01816_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__and4b_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _03423_ _03424_ _03425_ _03426_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__a211o_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ _03351_ _03352_ _03356_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__a21oi_2
X_07602_ _02308_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__buf_4
X_08582_ genblk2\[10\].wave_shpr.div.fin_quo\[1\] _03286_ _03288_ VGND VGND VPWR VPWR
+ _03289_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07533_ _02248_ _02249_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout158_A net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07464_ _02194_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07630__B _02336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09203_ net1251 _01302_ _03822_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06415_ _01358_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__buf_4
XFILLER_0_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07395_ _02080_ _02140_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09134_ _03754_ _03780_ _03781_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__a21o_1
X_06346_ genblk1\[0\].osc.clkdiv_C.cnt\[13\] _01291_ genblk1\[0\].osc.clkdiv_C.cnt\[14\]
+ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09065_ net1184 _01185_ _03722_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__mux2_1
XANTENNA__10483__S _04704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06277_ _01173_ _01188_ _01191_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_130_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10982__B1 _05054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08016_ genblk1\[6\].osc.clkdiv_C.cnt\[6\] _01750_ _01739_ genblk1\[6\].osc.clkdiv_C.cnt\[7\]
+ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold630 genblk1\[7\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold641 genblk2\[10\].wave_shpr.div.acc\[17\] VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold652 genblk2\[10\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 genblk2\[4\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold674 genblk2\[9\].wave_shpr.div.acc\[23\] VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 genblk2\[2\].wave_shpr.div.acc\[8\] VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 genblk2\[2\].wave_shpr.div.acc_next\[0\] VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__dlygate4sd3_1
X_09967_ genblk2\[3\].wave_shpr.div.acc\[15\] genblk2\[3\].wave_shpr.div.b1\[15\]
+ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__or2b_1
X_08918_ net612 _02260_ _03617_ _03574_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__a22o_1
X_09898_ genblk2\[2\].wave_shpr.div.acc\[11\] _04313_ _04301_ VGND VGND VPWR VPWR
+ _04314_ sky130_fd_sc_hd__mux2_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08849_ _03498_ _03553_ _03554_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08384__A_N _01437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07902__A1 genblk1\[8\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11860_ net1060 _05684_ _05685_ _05697_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__a22o_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10811_ _04855_ _04957_ _04958_ _04858_ net1117 VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__a32o_1
X_11791_ genblk2\[9\].wave_shpr.div.acc_next\[0\] _03693_ VGND VGND VPWR VPWR _05645_
+ sky130_fd_sc_hd__or2b_1
XANTENNA__09037__B1_N _03705_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09655__A1 _04045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06469__A1 genblk1\[1\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13530_ clknet_leaf_98_clk _00847_ net169 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11462__A1 _01797_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10742_ net772 _04886_ _04890_ _04908_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10673_ net500 _04861_ _04862_ net572 _04863_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__a221o_1
X_13461_ clknet_leaf_84_clk _00778_ net203 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12412_ genblk2\[11\].wave_shpr.div.acc\[15\] _06081_ _06055_ VGND VGND VPWR VPWR
+ _06082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13392_ clknet_leaf_91_clk _00711_ net143 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12343_ genblk2\[11\].wave_shpr.div.acc_next\[0\] _03942_ _03941_ net412 _06029_
+ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08630__A2 _02733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12274_ _05998_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08090__C _02365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11225_ genblk2\[7\].wave_shpr.div.quo\[8\] _05246_ _05250_ net421 VGND VGND VPWR
+ VPWR _00719_ sky130_fd_sc_hd__a22o_1
X_11156_ _05164_ _05214_ _05215_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10107_ _04269_ genblk1\[3\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__and2_1
X_11087_ genblk2\[6\].wave_shpr.div.acc\[25\] _05021_ genblk2\[6\].wave_shpr.div.acc\[24\]
+ genblk2\[6\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__or4b_1
X_10038_ _04428_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08449__A2 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11989_ _05799_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13728_ clknet_leaf_97_clk _01039_ net167 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06347__A genblk1\[0\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13659_ clknet_leaf_47_clk net475 net120 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06200_ PWM.counter\[4\] _01161_ net810 VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11205__A1 _03831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07180_ genblk1\[9\].osc.clkdiv_C.cnt\[8\] genblk1\[9\].osc.clkdiv_C.cnt\[7\] _01967_
+ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06131_ net3 _01102_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12084__A _05815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09821_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09752_ genblk2\[3\].wave_shpr.div.b1\[0\] _04223_ _04039_ VGND VGND VPWR VPWR _04224_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_123_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10332__A _03717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06964_ genblk1\[7\].osc.clkdiv_C.cnt\[4\] _01799_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__xnor2_1
X_08703_ _02586_ _03409_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__nand2_1
X_09683_ genblk2\[2\].wave_shpr.div.acc\[10\] genblk2\[2\].wave_shpr.div.b1\[10\]
+ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__or2b_1
X_06895_ genblk1\[6\].osc.clkdiv_C.cnt\[15\] _01362_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__nor2_1
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ genblk2\[8\].wave_shpr.div.fin_quo\[0\] genblk2\[8\].wave_shpr.div.fin_quo\[1\]
+ _02638_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_138_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _02261_ _03270_ _03271_ _02950_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07516_ PWM.final_sample_in\[1\] _02235_ PWM.counter\[1\] VGND VGND VPWR VPWR _02236_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08496_ _03054_ _03076_ _03075_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout46 net47 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07447_ _02182_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__clkbuf_4
Xfanout57 net58 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout68 net85 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout79 net84 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07378_ _02128_ _02127_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11747__A2 _05623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11135__A_N genblk2\[7\].wave_shpr.div.b1\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06329_ net592 _01281_ _01283_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__a21oi_1
X_09117_ genblk2\[0\].wave_shpr.div.acc\[0\] genblk2\[0\].wave_shpr.div.b1\[0\] VGND
+ VGND VPWR VPWR _03765_ sky130_fd_sc_hd__and2b_1
XFILLER_0_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08612__A2 _02521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10955__B1 _05055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06704__B _01592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09048_ genblk2\[0\].wave_shpr.div.b1\[4\] _03712_ _03708_ VGND VGND VPWR VPWR _03713_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold460 sig_norm.acc\[8\] VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold471 _00168_ VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout90_A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold482 genblk2\[9\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ net907 _05086_ _05093_ _05096_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12172__A2 _05818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold493 genblk2\[2\].wave_shpr.div.i\[2\] VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06387__B1 _01329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11380__B1 _03855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12961_ clknet_leaf_139_clk _00290_ net39 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11912_ genblk2\[10\].wave_shpr.div.acc\[14\] genblk2\[10\].wave_shpr.div.b1\[14\]
+ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__or2b_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ clknet_leaf_28_clk net463 net91 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _02203_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__clkbuf_4
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10238__A2 _04457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ genblk2\[9\].wave_shpr.div.quo\[17\] _05628_ _05629_ net349 _05636_ VGND
+ VGND VPWR VPWR _00882_ sky130_fd_sc_hd__a221o_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13513_ clknet_leaf_78_clk _00830_ net205 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10725_ net885 _04886_ _04890_ _04895_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__a22o_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11801__A _02203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13444_ clknet_leaf_95_clk net382 net149 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10656_ _04856_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12108__S _05865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10587_ _04763_ _04813_ _04814_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__a21o_1
XANTENNA__08603__A2 _02885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13375_ clknet_leaf_86_clk _00694_ net179 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_106_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10946__B1 _05056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10417__A _04672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12326_ _03689_ genblk1\[11\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12257_ genblk2\[11\].wave_shpr.div.fin_quo\[6\] net1332 _00005_ VGND VGND VPWR VPWR
+ _05989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12163__A2 _05818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11208_ _03726_ _05243_ _03736_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07726__A _01342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12188_ genblk2\[11\].wave_shpr.div.b1\[16\] genblk2\[11\].wave_shpr.div.acc\[16\]
+ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__xor2_1
X_11139_ genblk2\[7\].wave_shpr.div.b1\[9\] genblk2\[7\].wave_shpr.div.acc\[9\] VGND
+ VGND VPWR VPWR _05199_ sky130_fd_sc_hd__and2b_1
XANTENNA__07590__A2 _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06680_ genblk1\[4\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__inv_2
XANTENNA__07461__A _02155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08350_ genblk2\[5\].wave_shpr.div.fin_quo\[4\] _03056_ _02527_ VGND VGND VPWR VPWR
+ _03057_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07301_ genblk1\[11\].osc.clkdiv_C.cnt\[6\] _01595_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__nor2_1
X_08281_ genblk2\[9\].wave_shpr.div.fin_quo\[5\] _02521_ _02310_ VGND VGND VPWR VPWR
+ _02988_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07232_ genblk1\[10\].osc.clkdiv_C.cnt\[0\] _01321_ _02013_ genblk1\[10\].osc.clkdiv_C.cnt\[3\]
+ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07163_ genblk1\[9\].osc.clkdiv_C.cnt\[3\] _01958_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06114_ net368 _01086_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07094_ genblk1\[8\].osc.clkdiv_C.cnt\[9\] _01900_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10046__B _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout203 net204 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09555__B1 _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout214 net217 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09804_ genblk2\[2\].wave_shpr.div.quo\[5\] _04248_ _04252_ net696 VGND VGND VPWR
+ VPWR _00296_ sky130_fd_sc_hd__a22o_1
X_07996_ _02701_ _02702_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__or2b_1
XANTENNA__07581__A2 _01437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09735_ genblk2\[2\].wave_shpr.div.fin_quo\[0\] _04214_ _00009_ VGND VGND VPWR VPWR
+ _04215_ sky130_fd_sc_hd__mux2_1
X_06947_ net1104 _01783_ _01786_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10997__A _05051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09666_ _04045_ _04148_ _04149_ _04048_ net1091 VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__a32o_1
X_06878_ _01731_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__buf_4
X_08617_ genblk2\[4\].wave_shpr.div.fin_quo\[2\] _02362_ _02838_ VGND VGND VPWR VPWR
+ _03324_ sky130_fd_sc_hd__a21o_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ net847 _04076_ _04080_ _04099_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07090__B genblk1\[8\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08548_ _02742_ _03254_ _02745_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__o21a_1
X_08479_ _02838_ _03185_ _02846_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__o21a_1
X_10510_ _04745_ _04619_ genblk2\[4\].wave_shpr.div.acc\[22\] VGND VGND VPWR VPWR
+ _04747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11490_ _05440_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10441_ net970 _04683_ _04690_ _04695_ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__a22o_1
XANTENNA__08046__B1 _01666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10372_ genblk2\[4\].wave_shpr.div.quo\[1\] _04652_ _04656_ net418 VGND VGND VPWR
+ VPWR _00460_ sky130_fd_sc_hd__a22o_1
X_13160_ clknet_leaf_122_clk _00485_ net78 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12111_ _05763_ _05870_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13091_ clknet_leaf_137_clk _00418_ net39 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12042_ _05815_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__clkbuf_4
Xhold290 genblk2\[4\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09761__A _01436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12944_ clknet_leaf_2_clk _00273_ net42 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11656__A1 _05449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07324__A2 _01334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ clknet_leaf_138_clk _00206_ net39 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _05588_ _05563_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__or2b_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07088__A1 genblk1\[8\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_134_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_134_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ genblk2\[9\].wave_shpr.div.quo\[10\] _03696_ _03694_ net290 _05626_ VGND
+ VGND VPWR VPWR _00875_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10092__B1 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10708_ _04855_ _04881_ _04882_ _04858_ net1062 VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__a32o_1
X_11688_ _05570_ _05578_ _05579_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13427_ clknet_leaf_87_clk _00746_ net201 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10639_ net1248 _04225_ _04834_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13358_ clknet_leaf_4_clk _00679_ net46 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08052__A3 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12309_ genblk2\[11\].wave_shpr.div.quo\[9\] _03947_ _03944_ net355 _06011_ VGND
+ VGND VPWR VPWR _01042_ sky130_fd_sc_hd__a221o_1
X_13289_ clknet_leaf_92_clk _00610_ net147 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_07850_ genblk2\[1\].wave_shpr.div.fin_quo\[2\] _02461_ _02462_ _02316_ VGND VGND
+ VPWR VPWR _02557_ sky130_fd_sc_hd__a31o_1
XANTENNA__10698__A2 _02183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07563__A2 _01556_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06801_ _01669_ _01559_ _01671_ _01436_ _01672_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__a221o_1
X_07781_ genblk1\[0\].osc.clkdiv_C.cnt\[5\] _02483_ _02484_ _02486_ _02487_ VGND VGND
+ VPWR VPWR _02488_ sky130_fd_sc_hd__a2111o_1
Xinput3 pb[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_4
X_09520_ _03855_ _01330_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06732_ _01616_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__inv_2
XANTENNA__07903__B _01360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07315__A2 _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09451_ _04013_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__clkbuf_1
X_06663_ _01524_ _01553_ _01554_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08402_ genblk1\[2\].osc.clkdiv_C.cnt\[11\] _01411_ _03102_ _03106_ _03108_ VGND
+ VGND VPWR VPWR _03109_ sky130_fd_sc_hd__a2111o_1
X_06594_ genblk1\[3\].osc.clkdiv_C.cnt\[6\] _01500_ _01496_ genblk1\[3\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__o2bb2a_1
X_09382_ genblk2\[11\].wave_shpr.div.i\[1\] genblk2\[11\].wave_shpr.div.i\[0\] genblk2\[11\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__and3_1
XFILLER_0_148_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08333_ _03037_ _03038_ _03039_ _02694_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__a211o_1
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_125_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_125_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout140_A net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08264_ _02915_ _02910_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__or2b_1
XFILLER_0_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07215_ _01490_ _01993_ genblk1\[10\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR _01997_
+ sky130_fd_sc_hd__o21ai_1
X_08195_ _02349_ _02351_ _02355_ genblk2\[11\].wave_shpr.div.fin_quo\[5\] VGND VGND
+ VPWR VPWR _02902_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_61_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07146_ _01336_ _01496_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__nor2_4
XFILLER_0_30_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10491__S _04704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07077_ genblk1\[8\].osc.clkdiv_C.cnt\[3\] _01890_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07979_ genblk2\[7\].wave_shpr.div.fin_quo\[0\] genblk2\[7\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__nor2_1
X_09718_ _04161_ _04196_ _04197_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__a21o_1
X_10990_ genblk2\[6\].wave_shpr.div.b1\[0\] _05023_ genblk2\[6\].wave_shpr.div.acc\[0\]
+ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout53_A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07306__A2 _01678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09649_ genblk2\[1\].wave_shpr.div.acc\[22\] _04109_ _04113_ _04138_ VGND VGND VPWR
+ VPWR _00255_ sky130_fd_sc_hd__a22o_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ clknet_leaf_26_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[9\] net87 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ net947 _05507_ _05445_ _05519_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08267__B1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_116_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_116_clk sky130_fd_sc_hd__clkbuf_16
X_12591_ clknet_leaf_13_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[12\] net70 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11542_ genblk2\[8\].wave_shpr.div.quo\[23\] _05441_ _05458_ net229 _05468_ VGND
+ VGND VPWR VPWR _00818_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11473_ genblk2\[9\].wave_shpr.div.b1\[7\] _04230_ _05433_ VGND VGND VPWR VPWR _05434_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09767__B1 _04233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13212_ clknet_leaf_25_clk _00535_ net86 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10424_ _04681_ _04682_ net1129 _04652_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_104_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08660__A _02789_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13143_ clknet_leaf_121_clk net252 net81 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10355_ genblk2\[5\].wave_shpr.div.b1\[13\] _04645_ _04637_ VGND VGND VPWR VPWR _04646_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10286_ genblk2\[4\].wave_shpr.div.b1\[8\] genblk2\[4\].wave_shpr.div.acc\[8\] VGND
+ VGND VPWR VPWR _04598_ sky130_fd_sc_hd__and2b_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ clknet_leaf_11_clk net437 net56 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_12025_ net682 _05813_ _05817_ net724 VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__a22o_1
XANTENNA__12121__S _05865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12927_ clknet_leaf_35_clk _00258_ net106 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06505__B1 _01196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12858_ clknet_leaf_134_clk _00189_ net60 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08835__A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__13056__RESET_B net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11809_ genblk2\[9\].wave_shpr.div.acc\[3\] _05658_ _05613_ VGND VGND VPWR VPWR _05659_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_107_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_107_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12789_ clknet_leaf_43_clk _00122_ net124 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12357__A _03942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06355__A genblk1\[0\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07000_ genblk1\[7\].osc.clkdiv_C.cnt\[4\] _01827_ genblk1\[7\].osc.clkdiv_C.cnt\[5\]
+ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09222__A2 _03836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06802__B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12109__A2 _05844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08951_ _03641_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07902_ genblk1\[8\].osc.clkdiv_C.cnt\[12\] _01328_ _02607_ _02608_ VGND VGND VPWR
+ VPWR _02609_ sky130_fd_sc_hd__a211o_1
X_08882_ sig_norm.acc\[7\] sig_norm.acc\[6\] sig_norm.acc\[5\] _03587_ VGND VGND VPWR
+ VPWR _03588_ sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_4_4_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07833_ genblk2\[1\].wave_shpr.div.fin_quo\[5\] _02539_ _02469_ VGND VGND VPWR VPWR
+ _02540_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout188_A net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07764_ _02465_ _02466_ _02470_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09503_ _03714_ _04041_ _03736_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__o21ai_1
X_06715_ _01600_ _01602_ _01603_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07695_ _02016_ _02390_ _02393_ _02400_ _02401_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__a221oi_2
X_09434_ genblk2\[1\].wave_shpr.div.b1\[14\] genblk2\[1\].wave_shpr.div.acc\[14\]
+ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__and2b_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06646_ _01486_ _01542_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09365_ _03934_ _03802_ genblk2\[0\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR
+ _03936_ sky130_fd_sc_hd__mux2_1
X_06577_ genblk1\[3\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__inv_2
XANTENNA__12267__A _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08316_ _02419_ _03022_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06265__A _01224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09296_ _03774_ _03884_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08247_ genblk2\[8\].wave_shpr.div.fin_quo\[5\] _02638_ _02952_ _02223_ VGND VGND
+ VPWR VPWR _02954_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10359__A1 _01365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08178_ _02853_ _02878_ _02884_ genblk1\[3\].osc.clkdiv_C.cnt\[17\] genblk1\[3\].osc.clkdiv_C.cnt\[16\]
+ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__a311o_4
XANTENNA__11556__B1 _05448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07129_ genblk1\[9\].osc.clkdiv_C.cnt\[9\] _01801_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10140_ _04454_ _04481_ _04482_ _04457_ net1067 VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__a32o_1
XANTENNA__07775__A2 _01227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10234__B _04480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10071_ net1281 _01595_ _04440_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__mux2_1
XANTENNA__10250__A _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_cap21 net1350 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
XFILLER_0_97_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13761_ clknet_leaf_70_clk _01072_ net214 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10973_ net313 _05062_ _05064_ net486 _05071_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12712_ clknet_leaf_55_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[7\] net175 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13692_ clknet_leaf_44_clk _01003_ net122 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12643_ clknet_leaf_10_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[10\] net56 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12574_ clknet_leaf_29_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[13\] net89 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11525_ genblk2\[8\].wave_shpr.div.quo\[15\] _05454_ _05458_ net237 _05459_ VGND
+ VGND VPWR VPWR _00810_ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12339__A2 _03942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11456_ genblk2\[8\].wave_shpr.div.fin_quo\[7\] net1335 _00021_ VGND VGND VPWR VPWR
+ _05425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07215__A1 _01490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10407_ _04268_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__buf_2
XANTENNA__12116__S _05865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07718__B _01302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10425__A _04651_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11387_ genblk2\[8\].wave_shpr.div.acc\[12\] genblk2\[8\].wave_shpr.div.b1\[12\]
+ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13126_ clknet_leaf_3_clk _00451_ net51 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10338_ _03831_ net625 _03733_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__a21bo_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ clknet_leaf_24_clk net539 net92 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10269_ genblk2\[4\].wave_shpr.div.acc\[3\] genblk2\[4\].wave_shpr.div.b1\[3\] VGND
+ VGND VPWR VPWR _04581_ sky130_fd_sc_hd__or2b_1
XFILLER_0_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12008_ genblk2\[11\].wave_shpr.div.b1\[13\] _01483_ _05802_ VGND VGND VPWR VPWR
+ _05809_ sky130_fd_sc_hd__mux2_1
XANTENNA__12275__A1 _01311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06500_ genblk1\[2\].osc.clkdiv_C.cnt\[13\] genblk1\[2\].osc.clkdiv_C.cnt\[0\] net35
+ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__and3_1
X_07480_ genblk2\[10\].wave_shpr.div.i\[1\] _02205_ genblk2\[10\].wave_shpr.div.i\[4\]
+ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__or3b_1
XFILLER_0_124_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06431_ net29 VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09150_ _03746_ _03796_ _03797_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06362_ genblk1\[1\].osc.clkdiv_C.cnt\[5\] _01305_ VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11786__B1 _03693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08101_ _02804_ _02807_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__or2_1
X_09081_ _03704_ net396 _03717_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__a21bo_1
X_06293_ _01196_ _01254_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08032_ _02699_ genblk2\[6\].wave_shpr.div.fin_quo\[6\] _02734_ _02738_ _02261_ VGND
+ VGND VPWR VPWR _02739_ sky130_fd_sc_hd__a41o_1
XFILLER_0_114_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06813__A genblk1\[5\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold801 genblk2\[1\].wave_shpr.div.acc\[14\] VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold812 genblk2\[7\].wave_shpr.div.acc\[5\] VGND VGND VPWR VPWR net1030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 genblk2\[5\].wave_shpr.div.acc\[25\] VGND VGND VPWR VPWR net1041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold834 genblk2\[8\].wave_shpr.div.acc\[25\] VGND VGND VPWR VPWR net1052 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11387__B_N genblk2\[8\].wave_shpr.div.b1\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold845 genblk1\[6\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR net1063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold856 genblk2\[4\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR net1074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 genblk2\[9\].wave_shpr.div.quo\[7\] VGND VGND VPWR VPWR net1085 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold878 genblk2\[6\].wave_shpr.div.b1\[16\] VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 genblk2\[1\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ genblk2\[3\].wave_shpr.div.b1\[1\] VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08934_ _01099_ _00024_ _03627_ _03628_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__a31o_1
XANTENNA__07644__A _02350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08865_ _03009_ _03134_ _03571_ _02248_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__o31ai_2
X_07816_ genblk2\[1\].wave_shpr.div.fin_quo\[3\] _02522_ VGND VGND VPWR VPWR _02523_
+ sky130_fd_sc_hd__xor2_1
X_08796_ _03395_ _03499_ _03484_ _03498_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__a211oi_2
X_07747_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] _01172_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07678_ genblk1\[10\].osc.clkdiv_C.cnt\[9\] _01215_ _01991_ _02003_ VGND VGND VPWR
+ VPWR _02385_ sky130_fd_sc_hd__a2bb2o_1
X_09417_ _03966_ _03979_ _03980_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__o21bai_1
X_06629_ net1077 _01530_ _01532_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08194__B net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09348_ _03798_ net23 genblk2\[0\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR _03925_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09279_ _03766_ _03871_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__xnor2_1
X_11310_ genblk2\[7\].wave_shpr.div.acc\[10\] _05306_ _05300_ VGND VGND VPWR VPWR
+ _05307_ sky130_fd_sc_hd__mux2_1
XANTENNA__07819__A _02525_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12290_ net1299 _01249_ _05994_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11241_ _04268_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_120_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11172_ _05227_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10792__A2_N _04880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06956__B1 _01732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10123_ genblk2\[3\].wave_shpr.div.quo\[20\] _04461_ _04462_ net296 _04472_ VGND
+ VGND VPWR VPWR _00395_ sky130_fd_sc_hd__a221o_1
XANTENNA__06420__A2 _01363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07554__A _02223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10054_ _01557_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__inv_2
XANTENNA__07920__A2 _01430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13330__RESET_B net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13744_ clknet_leaf_51_clk _01055_ net110 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10956_ _05051_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__buf_2
XANTENNA__09205__B1_N _03728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13675_ clknet_leaf_42_clk _00988_ net125 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10887_ _05027_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12626_ clknet_leaf_16_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[11\] net74 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12557_ clknet_leaf_55_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[14\] net175 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11508_ _05444_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12488_ clknet_leaf_107_clk _00050_ net151 VGND VGND VPWR VPWR sig_norm.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold108 genblk2\[3\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold119 _00295_ VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ genblk2\[8\].wave_shpr.div.acc\[25\] genblk2\[8\].wave_shpr.div.acc\[26\]
+ _05414_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06352__B genblk1\[0\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07739__A2 _01334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ clknet_leaf_114_clk _00434_ net133 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ genblk1\[7\].osc.clkdiv_C.cnt\[16\] _01578_ _01574_ genblk1\[7\].osc.clkdiv_C.cnt\[7\]
+ _01815_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08650_ _03351_ _03352_ _03356_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__and3_2
X_07601_ _02307_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__buf_4
XANTENNA__07911__A2 _01308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08581_ _03285_ _03287_ _02404_ _02525_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__o31a_1
XFILLER_0_88_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07532_ _01151_ _02245_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__nor2_1
XANTENNA__13000__RESET_B net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07463_ _02191_ _02153_ genblk2\[7\].wave_shpr.div.busy VGND VGND VPWR VPWR _02194_
+ sky130_fd_sc_hd__and3b_1
XANTENNA__07630__C net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09202_ _03829_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06414_ _01178_ freq_div.state\[2\] VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07394_ _02080_ _02140_ _02142_ _02092_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11759__B1 _03694_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09133_ genblk2\[0\].wave_shpr.div.b1\[9\] genblk2\[0\].wave_shpr.div.acc\[9\] VGND
+ VGND VPWR VPWR _03781_ sky130_fd_sc_hd__and2b_1
XANTENNA__11223__A2 _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06345_ genblk1\[0\].osc.clkdiv_C.cnt\[13\] _01291_ _01293_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06276_ _01237_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__clkbuf_8
X_09064_ _03723_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08015_ _02721_ _02719_ genblk1\[6\].osc.clkdiv_C.cnt\[6\] _01750_ VGND VGND VPWR
+ VPWR _02722_ sky130_fd_sc_hd__a2bb2o_1
Xhold620 genblk2\[6\].wave_shpr.div.acc\[12\] VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 genblk2\[3\].wave_shpr.div.quo\[4\] VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold642 _00992_ VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold653 genblk2\[8\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 genblk2\[5\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 genblk2\[7\].wave_shpr.div.acc\[7\] VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 genblk2\[3\].wave_shpr.div.acc\[19\] VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 _00317_ VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06402__A2 _01340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09966_ _04245_ genblk2\[3\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR _04362_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09065__S _03722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08917_ sig_norm.acc\[6\] _03614_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__xnor2_1
X_09897_ _04194_ _04312_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__xnor2_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08155__A2 _01483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08848_ _03498_ _03553_ _03554_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__or3_1
XANTENNA__07902__A2 _01328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ _02518_ _02566_ _02570_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__a21oi_1
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ genblk2\[5\].wave_shpr.div.i\[1\] genblk2\[5\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _04958_ sky130_fd_sc_hd__nand2_1
X_11790_ genblk2\[9\].wave_shpr.div.acc_next\[0\] _02203_ _03693_ net306 _05644_ VGND
+ VGND VPWR VPWR _00890_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08636__C genblk2\[8\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10741_ genblk2\[5\].wave_shpr.div.acc\[8\] _04906_ _04907_ VGND VGND VPWR VPWR _04908_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07666__B2 _01190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13460_ clknet_leaf_84_clk _00777_ net203 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_10672_ _04672_ genblk1\[5\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12411_ _05970_ _06080_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08615__B1 _02223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13391_ clknet_leaf_79_clk _00710_ net206 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_105_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12342_ _03689_ genblk1\[11\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR _06029_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_51_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06453__A genblk1\[1\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12273_ net1272 _05997_ _05994_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_12_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11224_ genblk2\[7\].wave_shpr.div.quo\[7\] _05246_ _05250_ net317 VGND VGND VPWR
+ VPWR _00718_ sky130_fd_sc_hd__a22o_1
X_11155_ genblk2\[7\].wave_shpr.div.b1\[17\] genblk2\[7\].wave_shpr.div.acc\[17\]
+ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__and2b_1
X_10106_ net387 _04461_ _04462_ net525 _04463_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__a221o_1
X_11086_ genblk2\[6\].wave_shpr.div.acc\[24\] _05021_ genblk2\[6\].wave_shpr.div.acc\[25\]
+ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_87_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_16
X_10037_ genblk2\[3\].wave_shpr.div.fin_quo\[5\] genblk2\[3\].wave_shpr.div.quo\[4\]
+ _04422_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__mux2_1
XANTENNA__11534__A _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09774__B1_N _03733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11988_ net1265 _01946_ _05433_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13727_ clknet_leaf_97_clk _01038_ net167 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10939_ _05054_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10661__B1 _04857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13658_ clknet_leaf_44_clk net335 net120 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12609_ clknet_leaf_22_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[12\] net94 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_144_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06880__A2 _01684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13589_ clknet_leaf_72_clk _00904_ net215 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06130_ _01100_ _01101_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10413__B1 _04654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08989__S _01155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12166__B1 _05818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09820_ net457 _04257_ _04259_ net553 _04260_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__a221o_1
XANTENNA__08385__A2 _01439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06810__B _01326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07194__A genblk1\[9\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09751_ _01211_ _01302_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__nor2_2
X_06963_ _01229_ _01230_ _01238_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__a21oi_4
Xclkbuf_leaf_78_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_16
X_08702_ _02561_ _02585_ _02548_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09682_ genblk2\[2\].wave_shpr.div.acc\[11\] genblk2\[2\].wave_shpr.div.b1\[11\]
+ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__or2b_1
X_06894_ genblk1\[6\].osc.clkdiv_C.cnt\[5\] _01747_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09613__S _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08633_ _02742_ _03338_ _03339_ _02745_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout170_A net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ genblk2\[7\].wave_shpr.div.fin_quo\[2\] _02521_ VGND VGND VPWR VPWR _03271_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07515_ PWM.next_counter\[0\] PWM.final_sample_in\[0\] VGND VGND VPWR VPWR _02235_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_65_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08495_ _03175_ _03200_ _03201_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__nor3_2
XFILLER_0_9_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout47 net50 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
XFILLER_0_9_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07446_ _02147_ _02181_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__nor2_1
Xfanout58 net85 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06320__A1 genblk1\[0\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout69 net75 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07377_ _02128_ _02127_ _02129_ _02092_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09116_ _03762_ _03763_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06328_ genblk1\[0\].osc.clkdiv_C.cnt\[7\] _01281_ _01270_ VGND VGND VPWR VPWR _01283_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__06273__A _01231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09047_ _01248_ _02374_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__nor2_2
XFILLER_0_142_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06259_ _01194_ _01175_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_130_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold450 genblk2\[6\].wave_shpr.div.quo\[24\] VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 genblk2\[7\].wave_shpr.div.acc\[21\] VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 genblk2\[8\].wave_shpr.div.acc\[20\] VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 genblk2\[1\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 genblk2\[9\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout83_A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09949_ _04349_ _04350_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_69_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_16
X_12960_ clknet_leaf_137_clk _00289_ net39 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11911_ genblk2\[10\].wave_shpr.div.acc\[15\] genblk2\[10\].wave_shpr.div.b1\[15\]
+ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__or2b_1
XANTENNA__07832__A _02309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ clknet_leaf_28_clk net512 net91 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ net1046 _05652_ _05653_ _05683_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _04676_ _01928_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ clknet_leaf_78_clk _00829_ net205 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ genblk2\[5\].wave_shpr.div.acc\[4\] _04894_ _04821_ VGND VGND VPWR VPWR _04895_
+ sky130_fd_sc_hd__mux2_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13443_ clknet_leaf_92_clk _00762_ net149 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10655_ _04854_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13374_ clknet_leaf_96_clk _00693_ net167 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10586_ genblk2\[5\].wave_shpr.div.b1\[17\] genblk2\[5\].wave_shpr.div.acc\[17\]
+ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09800__A2 _04248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12325_ genblk2\[11\].wave_shpr.div.quo\[16\] _06014_ _06015_ net351 _06020_ VGND
+ VGND VPWR VPWR _01049_ sky130_fd_sc_hd__a221o_1
XANTENNA__06614__A2 _01483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12256_ _05988_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__clkbuf_1
X_11207_ net703 VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__inv_2
XANTENNA__07726__B _01241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12187_ genblk2\[11\].wave_shpr.div.acc\[17\] genblk2\[11\].wave_shpr.div.b1\[17\]
+ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__or2b_1
X_11138_ _05173_ _05196_ _05197_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__a21o_1
X_11069_ net622 _05119_ _05126_ _05141_ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10882__A0 genblk2\[6\].wave_shpr.div.fin_quo\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08827__B1 _02468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07300_ _01182_ _01226_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__nor2_4
XFILLER_0_128_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08280_ _02985_ _02986_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07231_ _01225_ _01354_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__nor2_2
XFILLER_0_128_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06805__B _01362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08055__A1 _01309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07162_ _01953_ _01958_ _01959_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06113_ _01086_ net360 VGND VGND VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.next_cnt\[2\]
+ sky130_fd_sc_hd__nor2_1
X_07093_ genblk1\[8\].osc.clkdiv_C.cnt\[9\] _01900_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__and2_1
XANTENNA__09608__S _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout204 net210 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__buf_2
Xfanout215 net217 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_4
X_09803_ genblk2\[2\].wave_shpr.div.quo\[4\] _04248_ _04252_ net336 VGND VGND VPWR
+ VPWR _00295_ sky130_fd_sc_hd__a22o_1
X_07995_ genblk1\[6\].osc.clkdiv_C.cnt\[10\] _01484_ _01742_ genblk1\[6\].osc.clkdiv_C.cnt\[9\]
+ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__a22oi_1
X_09734_ _04213_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07581__A3 _01226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06946_ net1356 _01785_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__nor2_1
XANTENNA__08748__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12311__B1 _03944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07652__A _02316_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09665_ genblk2\[1\].wave_shpr.div.i\[1\] genblk2\[1\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _04149_ sky130_fd_sc_hd__nand2_1
X_06877_ _01177_ _01249_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08616_ _03321_ _03322_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__nor2_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ genblk2\[1\].wave_shpr.div.acc\[8\] _04098_ _04095_ VGND VGND VPWR VPWR _04099_
+ sky130_fd_sc_hd__mux2_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08186__C _02365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ genblk2\[6\].wave_shpr.div.fin_quo\[0\] _02527_ _02309_ genblk2\[6\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08478_ _03183_ _03184_ genblk2\[4\].wave_shpr.div.fin_quo\[4\] _02308_ VGND VGND
+ VPWR VPWR _03185_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_53_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07429_ _02155_ _02168_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07099__A genblk1\[8\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10440_ genblk2\[4\].wave_shpr.div.acc\[4\] _04694_ _04623_ VGND VGND VPWR VPWR _04695_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06882__A2_N _01732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10371_ _04654_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__buf_2
XFILLER_0_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12110_ _05764_ _05739_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13090_ clknet_leaf_137_clk _00417_ net39 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12041_ genblk2\[10\].wave_shpr.div.quo\[12\] _05823_ _05816_ net223 _05824_ VGND
+ VGND VPWR VPWR _00961_ sky130_fd_sc_hd__a221o_1
Xhold280 genblk2\[6\].wave_shpr.div.quo\[14\] VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 genblk2\[11\].wave_shpr.div.quo\[18\] VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09761__B _04229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12302__B1 _06010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12943_ clknet_leaf_111_clk _00272_ net130 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12874_ clknet_leaf_136_clk _00205_ net42 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08096__C _01359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ net839 _05652_ _05653_ _05670_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__a22o_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _05464_ genblk1\[9\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_79_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ genblk2\[5\].wave_shpr.div.b1\[0\] _04821_ genblk2\[5\].wave_shpr.div.acc\[0\]
+ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11687_ genblk2\[9\].wave_shpr.div.b1\[3\] genblk2\[9\].wave_shpr.div.acc\[3\] VGND
+ VGND VPWR VPWR _05579_ sky130_fd_sc_hd__and2b_1
XFILLER_0_153_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_122_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12346__C _05982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13426_ clknet_leaf_82_clk _00745_ net201 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10638_ _04846_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09234__B1 _03839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09785__A1 _04242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13357_ clknet_leaf_4_clk _00678_ net45 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10569_ _04772_ _04795_ _04796_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07737__A genblk1\[1\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12308_ _05835_ genblk1\[11\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__and2_1
X_13288_ clknet_leaf_90_clk _00609_ net147 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_137_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12239_ genblk2\[11\].wave_shpr.div.acc\[18\] _05976_ VGND VGND VPWR VPWR _05977_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07456__B _02153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06800_ genblk1\[5\].osc.clkdiv_C.cnt\[11\] _01667_ _01666_ genblk1\[5\].osc.clkdiv_C.cnt\[13\]
+ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08760__A2 _02521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07563__A3 _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07780_ genblk1\[0\].osc.clkdiv_C.cnt\[5\] _02483_ _01215_ genblk1\[0\].osc.clkdiv_C.cnt\[3\]
+ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput4 pb[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_06731_ genblk1\[4\].osc.clkdiv_C.cnt\[5\] genblk1\[4\].osc.clkdiv_C.cnt\[4\] _01609_
+ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__and3_1
XANTENNA__11647__A2 _05448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07903__C _02011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09450_ genblk2\[1\].wave_shpr.div.fin_quo\[1\] genblk2\[1\].wave_shpr.div.quo\[0\]
+ _00007_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__mux2_1
X_06662_ genblk1\[3\].osc.clkdiv_C.cnt\[16\] _01551_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07720__B1 _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08401_ genblk1\[2\].osc.clkdiv_C.cnt\[12\] _01591_ _03107_ VGND VGND VPWR VPWR _03108_
+ sky130_fd_sc_hd__a21bo_1
X_09381_ genblk2\[11\].wave_shpr.div.i\[1\] genblk2\[11\].wave_shpr.div.i\[0\] genblk2\[11\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__a21o_1
X_06593_ genblk1\[3\].osc.clkdiv_C.cnt\[14\] _01498_ _01500_ genblk1\[3\].osc.clkdiv_C.cnt\[6\]
+ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_59_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08332_ _02217_ _02553_ genblk2\[7\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR
+ _03039_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08263_ _02899_ _02923_ VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_4_0_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07214_ _01181_ _01187_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__nor2_4
XFILLER_0_27_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08194_ net3 net163 _02312_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__and3_1
XANTENNA__09225__B1 _03840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07145_ genblk1\[9\].osc.clkdiv_C.cnt\[8\] _01514_ _01513_ genblk1\[9\].osc.clkdiv_C.cnt\[7\]
+ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10386__A2 _04657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07076_ _01887_ _01890_ _01891_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07978_ genblk2\[7\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__inv_2
X_09717_ genblk2\[2\].wave_shpr.div.b1\[12\] genblk2\[2\].wave_shpr.div.acc\[12\]
+ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__and2b_1
X_06929_ _01761_ _01773_ _01774_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_97_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08197__B _02361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09648_ genblk2\[1\].wave_shpr.div.acc\[21\] _04136_ VGND VGND VPWR VPWR _04138_
+ sky130_fd_sc_hd__xor2_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ genblk2\[1\].wave_shpr.div.acc\[4\] _04085_ _04011_ VGND VGND VPWR VPWR _04086_
+ sky130_fd_sc_hd__mux2_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11610_ net846 _05518_ _05493_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__mux2_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ clknet_leaf_13_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[11\] net70 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11541_ _05464_ genblk1\[8\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11472_ _03707_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__clkbuf_4
X_13211_ clknet_leaf_25_clk _00534_ net86 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10423_ genblk2\[4\].wave_shpr.div.b1\[0\] genblk2\[4\].wave_shpr.div.acc\[0\] _04623_
+ _04679_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__a31o_1
XANTENNA__09767__A1 _03704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13142_ clknet_leaf_115_clk _00467_ net135 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10354_ _01490_ _01242_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ clknet_leaf_23_clk net562 net98 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10285_ _04575_ _04595_ _04596_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__a21o_1
XANTENNA__10129__A2 _04451_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12024_ genblk2\[10\].wave_shpr.div.quo\[2\] _05813_ _05817_ net220 VGND VGND VPWR
+ VPWR _00951_ sky130_fd_sc_hd__a22o_1
XANTENNA__11526__B genblk1\[8\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12926_ clknet_leaf_35_clk _00257_ net106 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06505__A1 _01362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ clknet_leaf_91_clk _00188_ net146 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _05578_ _05657_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__xnor2_1
X_12788_ clknet_leaf_43_clk _00121_ net124 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11739_ _01099_ _01147_ _05622_ net1161 VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_83_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09758__A1 _04227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13409_ clknet_leaf_90_clk net549 net144 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07769__B1 _01240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07233__A2 _01363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08950_ sig_norm.quo\[3\] _03640_ _00024_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__mux2_1
X_07901_ genblk1\[8\].osc.clkdiv_C.cnt\[13\] _01246_ _01328_ genblk1\[8\].osc.clkdiv_C.cnt\[12\]
+ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__o22ai_1
X_08881_ sig_norm.acc\[4\] _03586_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07832_ _02309_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07763_ genblk2\[1\].wave_shpr.div.fin_quo\[6\] _02468_ _02469_ VGND VGND VPWR VPWR
+ _02470_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09502_ net761 VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06714_ genblk1\[4\].osc.clkdiv_C.cnt\[1\] genblk1\[4\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01603_ sky130_fd_sc_hd__nand2_1
X_07694_ _02386_ _02392_ _02387_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__and3_1
XFILLER_0_154_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09433_ _03958_ _03995_ _03996_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06645_ genblk1\[3\].osc.clkdiv_C.cnt\[10\] _01540_ _01542_ _01524_ VGND VGND VPWR
+ VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o211a_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09364_ net1305 _03841_ _03910_ _03935_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06576_ _01182_ _01302_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__or2_2
X_08315_ _03019_ _03020_ _03021_ _02416_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__a211o_1
XFILLER_0_129_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09295_ _03775_ _03757_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__or2b_1
XANTENNA__06265__B _01226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09857__A _04247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08246_ _02638_ _02952_ genblk2\[8\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR
+ _02953_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08761__A net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11005__B1 _05056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08177_ _02868_ _02879_ _02883_ _02864_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11556__A1 _05449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07128_ genblk1\[9\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__inv_2
X_07059_ genblk1\[8\].osc.clkdiv_C.cnt\[4\] _01866_ _01869_ genblk1\[8\].osc.clkdiv_C.cnt\[12\]
+ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10070_ _04445_ VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__clkbuf_1
Xmax_cap22 net1351 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_1
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13760_ clknet_leaf_70_clk _01071_ net213 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10972_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12711_ clknet_leaf_56_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[6\] net175 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
X_13691_ clknet_leaf_44_clk _01002_ net122 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_69_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12642_ clknet_leaf_10_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[9\] net56 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12036__A2 _05818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06456__A genblk1\[1\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10047__B2 _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12573_ clknet_leaf_29_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[12\] net89 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11524_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11455_ _05424_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10706__A _04880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06903__B _01327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10406_ net626 _04661_ _04663_ net658 _04671_ VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11386_ genblk2\[8\].wave_shpr.div.acc\[13\] genblk2\[8\].wave_shpr.div.b1\[13\]
+ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__or2b_1
X_13125_ clknet_leaf_3_clk _00450_ net51 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10337_ _04636_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ clknet_leaf_134_clk _00383_ net63 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_10268_ _04578_ _04579_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__nand2_1
X_12007_ _05808_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__clkbuf_1
X_10199_ genblk2\[3\].wave_shpr.div.acc\[14\] _04527_ _04507_ VGND VGND VPWR VPWR
+ _04528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12909_ clknet_leaf_31_clk _00240_ net100 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_06430_ net718 _01373_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12027__A2 _05813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06366__A _01308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06361_ _01223_ _01226_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__or2_2
XANTENNA__13206__RESET_B net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08100_ genblk1\[4\].osc.clkdiv_C.cnt\[12\] _02805_ _02806_ VGND VGND VPWR VPWR _02807_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_127_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09080_ _03732_ net577 _03733_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__o21a_1
X_06292_ _01176_ _01178_ _01194_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__and3b_2
XFILLER_0_140_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08031_ genblk2\[6\].wave_shpr.div.fin_quo\[4\] _02737_ VGND VGND VPWR VPWR _02738_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06813__B _01684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold802 genblk2\[11\].wave_shpr.div.acc\[3\] VGND VGND VPWR VPWR net1020 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07197__A genblk1\[9\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold813 genblk2\[6\].wave_shpr.div.acc\[22\] VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold824 genblk2\[9\].wave_shpr.div.b1\[9\] VGND VGND VPWR VPWR net1042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold835 genblk2\[7\].wave_shpr.div.acc\[25\] VGND VGND VPWR VPWR net1053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 genblk2\[3\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR net1064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 genblk2\[4\].wave_shpr.div.b1\[2\] VGND VGND VPWR VPWR net1075 sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ genblk2\[3\].wave_shpr.div.acc\[2\] genblk2\[3\].wave_shpr.div.b1\[2\] VGND
+ VGND VPWR VPWR _04378_ sky130_fd_sc_hd__or2b_1
Xhold868 genblk2\[11\].wave_shpr.div.b1\[16\] VGND VGND VPWR VPWR net1086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 genblk2\[5\].wave_shpr.div.b1\[7\] VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__dlygate4sd3_1
X_08933_ sig_norm.acc\[12\] _01157_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08864_ _03135_ _03225_ _03570_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__nor3_1
XANTENNA__10351__A _01355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07815_ genblk2\[1\].wave_shpr.div.fin_quo\[2\] _02462_ _02461_ VGND VGND VPWR VPWR
+ _02522_ sky130_fd_sc_hd__o21a_1
X_08795_ _03489_ _03496_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__or2_1
X_07746_ _02447_ _02446_ _02448_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07677_ _02377_ _02381_ _02368_ _02382_ _02383_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_66_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09416_ genblk2\[1\].wave_shpr.div.b1\[5\] genblk2\[1\].wave_shpr.div.acc\[5\] VGND
+ VGND VPWR VPWR _03980_ sky130_fd_sc_hd__and2b_1
XFILLER_0_137_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06628_ genblk1\[3\].osc.clkdiv_C.cnt\[4\] _01530_ _01524_ VGND VGND VPWR VPWR _01532_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__10029__A1 genblk2\[3\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09347_ _03799_ net23 VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__or2_1
X_06559_ _01451_ _01472_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09278_ genblk2\[0\].wave_shpr.div.b1\[2\] genblk2\[0\].wave_shpr.div.acc\[2\] VGND
+ VGND VPWR VPWR _03871_ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08229_ _02838_ _02935_ _02846_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11240_ net613 _05255_ _05256_ net640 _05259_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11171_ genblk2\[7\].wave_shpr.div.fin_quo\[4\] net1318 _00019_ VGND VGND VPWR VPWR
+ _05227_ sky130_fd_sc_hd__mux2_1
XANTENNA__12582__RESET_B net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10122_ _04058_ _01486_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__nor2_1
XANTENNA__08158__B1 _01858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10053_ _04435_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09370__A2 _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09658__B1 _04045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10955_ genblk2\[6\].wave_shpr.div.quo\[11\] _05057_ _05055_ net344 _05061_ VGND
+ VGND VPWR VPWR _00638_ sky130_fd_sc_hd__a221o_1
X_13743_ clknet_leaf_51_clk net240 net110 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13674_ clknet_leaf_41_clk _00987_ net125 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10886_ genblk2\[6\].wave_shpr.div.fin_quo\[3\] net1320 _00017_ VGND VGND VPWR VPWR
+ _05027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12625_ clknet_leaf_16_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[10\] net74 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__06892__B1 _01666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09497__A _03701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12556_ clknet_leaf_55_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[13\] net175 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11507_ _05441_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12487_ clknet_leaf_108_clk _00049_ net151 VGND VGND VPWR VPWR sig_norm.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold109 _00377_ VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__dlygate4sd3_1
X_11438_ genblk2\[8\].wave_shpr.div.acc\[24\] _05413_ VGND VGND VPWR VPWR _05414_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08397__B1 _02425_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_775 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11369_ _05349_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__clkbuf_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ clknet_leaf_127_clk _00433_ net133 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ clknet_leaf_126_clk _00366_ net61 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09361__A2 _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07600_ net17 net18 VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__and2_2
X_08580_ genblk2\[10\].wave_shpr.div.fin_quo\[1\] VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__inv_2
XANTENNA__07911__A3 _01440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07531_ _01155_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__buf_4
XFILLER_0_44_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06808__B _01359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07462_ _02193_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__inv_2
X_09201_ net1199 _01183_ _03822_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11208__B1 _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06413_ genblk1\[1\].osc.clkdiv_C.cnt\[9\] _01356_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07393_ genblk1\[11\].osc.clkdiv_C.cnt\[15\] _02139_ VGND VGND VPWR VPWR _02142_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_91_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09132_ _03755_ _03778_ _03779_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__a21o_1
X_06344_ genblk1\[0\].osc.clkdiv_C.cnt\[13\] _01291_ _01269_ VGND VGND VPWR VPWR _01293_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09063_ net1276 _03721_ _03722_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__mux2_1
X_06275_ _01178_ _01176_ _01194_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__nor3b_1
XANTENNA_fanout213_A net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10982__A2 _05051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08014_ genblk1\[6\].osc.clkdiv_C.cnt\[5\] _01367_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold610 genblk2\[5\].wave_shpr.div.acc\[17\] VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 genblk2\[9\].wave_shpr.div.acc\[8\] VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold632 genblk2\[4\].wave_shpr.div.acc\[14\] VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 genblk2\[0\].wave_shpr.div.b1\[0\] VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 genblk2\[8\].wave_shpr.div.acc\[3\] VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 genblk2\[6\].wave_shpr.div.acc\[13\] VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 genblk2\[7\].wave_shpr.div.acc\[11\] VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 genblk2\[1\].wave_shpr.div.acc\[15\] VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07655__A _02361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold698 genblk2\[7\].wave_shpr.div.acc\[9\] VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ genblk2\[3\].wave_shpr.div.acc\[17\] genblk2\[3\].wave_shpr.div.b1\[17\]
+ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__or2b_1
XANTENNA__11486__B1_N _03717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08916_ net1155 _02260_ _03616_ _03574_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__a22o_1
X_09896_ _04195_ _04162_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__or2b_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _03536_ _03537_ _03531_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__a21boi_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08778_ _03333_ _03483_ _03465_ _03482_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__a211oi_2
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ _01360_ net37 genblk1\[1\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _02436_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10740_ _04820_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__buf_4
XFILLER_0_138_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10671_ _04854_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12410_ _05971_ _05927_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__or2b_1
XANTENNA__08933__B _01157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13390_ clknet_leaf_79_clk _00709_ net205 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09812__B1 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12341_ net412 _03942_ _03941_ net434 _06028_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12272_ _01305_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__inv_2
X_11223_ net317 _05246_ _05250_ net754 VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11154_ _05165_ _05212_ _05213_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_101_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10105_ _04269_ genblk1\[3\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__and2_1
X_11085_ net1076 _05057_ _05055_ _05151_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__a22o_1
X_10036_ _04427_ VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__clkbuf_1
X_11987_ _05798_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__clkbuf_1
X_13726_ clknet_leaf_97_clk _01037_ net166 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10938_ net792 _05052_ _05023_ _05055_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13657_ clknet_leaf_48_clk _00970_ net120 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10869_ _04968_ _05011_ _05012_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12608_ clknet_leaf_23_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[11\] net94 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09803__B1 _04252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13588_ clknet_leaf_72_clk _00903_ net215 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09020__A _02152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12539_ clknet_leaf_62_clk _00091_ net189 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12166__A1 _05816_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07475__A _02155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09750_ net1198 VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__clkbuf_1
X_06962_ genblk1\[7\].osc.clkdiv_C.cnt\[9\] _01797_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__xnor2_1
X_08701_ _03359_ _03381_ _03406_ _03407_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__o211ai_2
X_09681_ genblk2\[2\].wave_shpr.div.acc\[12\] genblk2\[2\].wave_shpr.div.b1\[12\]
+ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__or2b_1
XFILLER_0_146_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06893_ _01308_ _01577_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__nand2_2
XANTENNA__08542__B1 _02308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08632_ _02217_ _02553_ genblk2\[6\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR
+ _03339_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08563_ genblk2\[7\].wave_shpr.div.fin_quo\[1\] _03269_ VGND VGND VPWR VPWR _03270_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout163_A net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07514_ PWM.counter\[2\] VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__inv_2
X_08494_ _03051_ _03174_ _03154_ _03173_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07445_ genblk2\[5\].wave_shpr.div.busy _02180_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout48 net50 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
Xfanout59 net63 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07376_ _02128_ _02127_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_889 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09115_ genblk2\[0\].wave_shpr.div.acc\[1\] genblk2\[0\].wave_shpr.div.b1\[1\] VGND
+ VGND VPWR VPWR _03763_ sky130_fd_sc_hd__or2b_1
X_06327_ _01269_ _01281_ _01282_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_17_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06273__B _01234_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10955__A2 _05057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09046_ _03711_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__clkbuf_1
X_06258_ freq_div.state\[1\] _01176_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__xor2_4
XFILLER_0_103_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold440 genblk2\[4\].wave_shpr.div.quo\[19\] VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__dlygate4sd3_1
X_06189_ net361 VGND VGND VPWR VPWR PWM.next_counter\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_102_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold451 genblk2\[9\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09076__S _03722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10707__A2 _04821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold462 genblk2\[4\].wave_shpr.div.quo\[16\] VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 genblk1\[8\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 genblk2\[0\].wave_shpr.div.b1\[17\] VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 genblk2\[9\].wave_shpr.div.b1\[16\] VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07584__A1 genblk1\[9\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06387__A2 _01323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07584__B2 genblk1\[9\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09948_ genblk2\[2\].wave_shpr.div.acc\[25\] _04212_ genblk2\[2\].wave_shpr.div.acc\[24\]
+ genblk2\[2\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout76_A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09879_ _04187_ _04166_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__or2b_1
X_11910_ _03832_ genblk2\[10\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR _05732_
+ sky130_fd_sc_hd__nor2_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10340__B1 _04432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12890_ clknet_leaf_28_clk _00221_ net91 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ genblk2\[9\].wave_shpr.div.acc\[11\] _05682_ _05673_ VGND VGND VPWR VPWR
+ _05683_ sky130_fd_sc_hd__mux2_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ genblk2\[9\].wave_shpr.div.quo\[16\] _05628_ _05629_ net304 _05635_ VGND
+ VGND VPWR VPWR _00881_ sky130_fd_sc_hd__a221o_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _04778_ _04788_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__xor2_1
XFILLER_0_55_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13511_ clknet_leaf_78_clk _00828_ net205 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10654_ net1342 _04853_ _04821_ _04855_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__a22o_1
X_13442_ clknet_leaf_92_clk _00761_ net149 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13373_ clknet_leaf_117_clk _00692_ net140 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10585_ _04764_ _04811_ _04812_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__o21bai_1
XANTENNA__10946__A2 _05052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12324_ _03689_ genblk1\[11\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12255_ genblk2\[11\].wave_shpr.div.fin_quo\[5\] net767 _00005_ VGND VGND VPWR VPWR
+ _05988_ sky130_fd_sc_hd__mux2_1
X_11206_ _03831_ net391 _03717_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__a21bo_1
X_12186_ net289 _05923_ _05924_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07575__A1 genblk1\[9\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold4_A modein.delay_in\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11137_ genblk2\[7\].wave_shpr.div.b1\[8\] genblk2\[7\].wave_shpr.div.acc\[8\] VGND
+ VGND VPWR VPWR _05197_ sky130_fd_sc_hd__and2b_1
X_11068_ _05139_ _05140_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__nand2_1
XANTENNA__08838__B _03544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10019_ genblk2\[3\].wave_shpr.div.acc\[18\] _04414_ VGND VGND VPWR VPWR _04415_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_149_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10882__A1 genblk2\[6\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13709_ clknet_leaf_31_clk _01020_ net103 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07230_ genblk1\[10\].osc.clkdiv_C.cnt\[6\] _01432_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12614__RESET_B net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06805__C _01226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07161_ genblk1\[9\].osc.clkdiv_C.cnt\[1\] genblk1\[9\].osc.clkdiv_C.cnt\[0\] genblk1\[9\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08055__A2 _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06112_ smpl_rt_clkdiv.clkDiv_inst.cnt\[1\] net338 net359 VGND VGND VPWR VPWR _01090_
+ sky130_fd_sc_hd__a21oi_1
X_07092_ _01887_ _01900_ _01901_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_10_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09555__A2 _04042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout205 net209 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_4
Xfanout216 net217 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_4
X_09802_ net336 _04248_ _04252_ net719 VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__a22o_1
X_07994_ genblk1\[6\].osc.clkdiv_C.cnt\[8\] _01732_ _01742_ genblk1\[6\].osc.clkdiv_C.cnt\[9\]
+ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__o22a_1
XANTENNA__07933__A genblk2\[8\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09733_ genblk2\[2\].wave_shpr.div.acc\[25\] genblk2\[2\].wave_shpr.div.acc\[24\]
+ genblk2\[2\].wave_shpr.div.acc\[26\] _04212_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__or4_2
X_06945_ genblk1\[6\].osc.clkdiv_C.cnt\[14\] _01783_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__and2_1
X_06876_ _01336_ net37 VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__or2_1
X_09664_ genblk2\[1\].wave_shpr.div.i\[1\] genblk2\[1\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _04148_ sky130_fd_sc_hd__or2_1
X_08615_ genblk2\[4\].wave_shpr.div.fin_quo\[0\] genblk2\[4\].wave_shpr.div.fin_quo\[1\]
+ _02932_ _02223_ VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__a31o_1
X_09595_ _03985_ _04097_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__xnor2_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _03251_ _03252_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__and2b_1
X_08477_ genblk2\[4\].wave_shpr.div.fin_quo\[3\] _02932_ _02840_ _02222_ VGND VGND
+ VPWR VPWR _03184_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07428_ genblk2\[3\].wave_shpr.div.busy _02167_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07359_ genblk1\[11\].osc.clkdiv_C.cnt\[7\] _02112_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10389__B1 _04655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10370_ net418 _04652_ _04623_ _04655_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09029_ _03694_ _03697_ _03699_ _03696_ net789 VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__a32o_1
XFILLER_0_131_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12040_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__and2_1
Xhold270 _00734_ VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _00641_ VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 genblk2\[11\].wave_shpr.div.quo\[17\] VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12942_ clknet_leaf_111_clk _00271_ net130 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06459__A genblk1\[1\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ clknet_leaf_138_clk _00204_ net39 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ genblk2\[9\].wave_shpr.div.acc\[7\] _05669_ _05613_ VGND VGND VPWR VPWR _05670_
+ sky130_fd_sc_hd__mux2_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09482__A1 _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ net290 _03696_ _03694_ net526 _05625_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10092__A2 _04452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10706_ _04880_ _04781_ genblk2\[5\].wave_shpr.div.b1\[0\] VGND VGND VPWR VPWR _04881_
+ sky130_fd_sc_hd__or3b_1
X_11686_ _05571_ _05576_ _05577_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13425_ clknet_leaf_87_clk _00744_ net201 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10637_ net1233 _04223_ _04834_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10568_ genblk2\[5\].wave_shpr.div.b1\[8\] genblk2\[5\].wave_shpr.div.acc\[8\] VGND
+ VGND VPWR VPWR _04796_ sky130_fd_sc_hd__and2b_1
X_13356_ clknet_leaf_4_clk _00677_ net45 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_2
X_12307_ net355 _06009_ _06010_ net358 VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10499_ net591 _04715_ _04722_ _04739_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__a22o_1
X_13287_ clknet_leaf_118_clk _00608_ net138 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12238_ _05925_ _05974_ _05975_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__a21o_1
X_12169_ net1226 _05818_ _05816_ _05913_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__a22o_1
XANTENNA__07753__A _02458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput5 pb[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_06730_ _01615_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06369__A _01192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06661_ genblk1\[3\].osc.clkdiv_C.cnt\[16\] _01551_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08400_ genblk1\[2\].osc.clkdiv_C.cnt\[13\] _02425_ _01591_ genblk1\[2\].osc.clkdiv_C.cnt\[12\]
+ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__o22a_1
XANTENNA__07720__B2 genblk1\[1\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09380_ _03944_ _03945_ _03946_ _03947_ net1124 VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__a32o_1
X_06592_ _01233_ _01437_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__nor2_2
X_08331_ _03036_ _02682_ _03035_ _02526_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__o31a_1
XANTENNA__09473__A1 _04023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06816__B _01355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08262_ _02945_ _02967_ _02968_ VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07213_ genblk1\[10\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__inv_2
X_08193_ _02423_ _02601_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09225__A1 net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout126_A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07144_ _01933_ _01941_ _01942_ _01943_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__and4b_1
XANTENNA__07236__B1 _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07075_ _01879_ _01889_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10354__A _01490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08200__A2 _02403_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07977_ genblk2\[7\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__inv_2
X_09716_ _04162_ _04194_ _04195_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__a21o_1
X_06928_ genblk1\[6\].osc.clkdiv_C.cnt\[7\] _01770_ genblk1\[6\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09647_ net1109 _04109_ _04113_ _04137_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06859_ _01693_ _01717_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__nor2_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09578_ _04084_ _03977_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__xnor2_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout39_A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ genblk2\[11\].wave_shpr.div.fin_quo\[0\] _02524_ _02307_ genblk2\[11\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09464__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08267__A2 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11540_ net229 _05441_ _05458_ net575 _05467_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11471_ _05432_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10422_ genblk2\[4\].wave_shpr.div.b1\[0\] _04623_ genblk2\[4\].wave_shpr.div.acc\[0\]
+ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__a21oi_1
X_13210_ clknet_leaf_25_clk _00533_ net86 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07778__A1 _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13141_ clknet_leaf_115_clk _00466_ net135 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10353_ _04644_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold874_A genblk1\[8\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13072_ clknet_leaf_23_clk net491 net94 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10284_ genblk2\[4\].wave_shpr.div.b1\[7\] genblk2\[4\].wave_shpr.div.acc\[7\] VGND
+ VGND VPWR VPWR _04596_ sky130_fd_sc_hd__and2b_1
X_12023_ net220 _05813_ _05817_ net740 VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__a22o_1
XANTENNA__07950__A1 _01556_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10203__S _04507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12925_ clknet_leaf_35_clk _00256_ net106 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06505__A2 _01430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ clknet_leaf_91_clk _00187_ net146 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _05579_ _05570_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__or2b_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12787_ clknet_leaf_43_clk _00120_ net124 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _02248_ _01150_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09207__A1 _03831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11669_ genblk2\[9\].wave_shpr.div.acc\[10\] genblk2\[9\].wave_shpr.div.b1\[10\]
+ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__or2b_1
XFILLER_0_114_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13408_ clknet_leaf_90_clk _00727_ net142 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07218__B1 _01442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_784 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13339_ clknet_leaf_7_clk _00660_ net49 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07900_ genblk1\[8\].osc.clkdiv_C.cnt\[14\] _01172_ _02605_ _02606_ VGND VGND VPWR
+ VPWR _02607_ sky130_fd_sc_hd__a211o_1
X_08880_ _03575_ sig_norm.acc\[3\] _03585_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__a21o_1
XANTENNA__10525__B1 _04657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09174__S _03722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07831_ genblk2\[1\].wave_shpr.div.fin_quo\[4\] _02461_ _02463_ _02224_ VGND VGND
+ VPWR VPWR _02538_ sky130_fd_sc_hd__a31o_1
X_07762_ _02458_ _02459_ _02220_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09501_ _03831_ net1025 _03717_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__a21bo_1
X_06713_ genblk1\[4\].osc.clkdiv_C.cnt\[1\] genblk1\[4\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01602_ sky130_fd_sc_hd__or2_1
X_07693_ _02399_ _02394_ _02385_ _02396_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09432_ genblk2\[1\].wave_shpr.div.b1\[13\] genblk2\[1\].wave_shpr.div.acc\[13\]
+ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__and2b_1
X_06644_ genblk1\[3\].osc.clkdiv_C.cnt\[10\] _01540_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09363_ genblk2\[0\].wave_shpr.div.acc\[23\] _03801_ _03934_ VGND VGND VPWR VPWR
+ _03935_ sky130_fd_sc_hd__a21o_1
X_06575_ _01196_ _01327_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__or2_4
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08249__A2 _02309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08314_ _02216_ _02552_ genblk2\[10\].wave_shpr.div.fin_quo\[4\] VGND VGND VPWR VPWR
+ _03021_ sky130_fd_sc_hd__and3_1
X_09294_ net866 _03870_ _03877_ _03883_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10068__B _01226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08245_ _02641_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08176_ _02880_ _02882_ _02870_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__a21o_1
X_07127_ genblk1\[9\].osc.clkdiv_C.cnt\[2\] _01920_ _01923_ genblk1\[9\].osc.clkdiv_C.cnt\[11\]
+ _01926_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__a221oi_1
XANTENNA_clkbuf_leaf_63_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06281__B _01242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07058_ genblk1\[8\].osc.clkdiv_C.cnt\[0\] _01211_ _01246_ genblk1\[8\].osc.clkdiv_C.cnt\[14\]
+ _01875_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_121_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_cap23 net1352 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
X_10971_ net486 _05062_ _05064_ net582 _05070_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap34 _01794_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_4
X_12710_ clknet_leaf_56_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[5\] net181 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
X_13690_ clknet_leaf_97_clk _00005_ net166 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_136_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12641_ clknet_leaf_10_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[8\] net56 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_109_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06456__B genblk1\[1\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12572_ clknet_leaf_28_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[11\] net89 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__12441__B1 _03944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07999__A1 _01200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11795__A2 _05613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11523_ _05444_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11454_ genblk2\[8\].wave_shpr.div.fin_quo\[6\] net1325 _00021_ VGND VGND VPWR VPWR
+ _05424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10405_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__and2_1
X_11385_ genblk2\[8\].wave_shpr.div.acc\[14\] genblk2\[8\].wave_shpr.div.b1\[14\]
+ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__or2b_1
XFILLER_0_104_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13124_ clknet_leaf_3_clk _00449_ net51 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10336_ net1287 _01256_ _04440_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__mux2_1
XANTENNA__07620__B1 _01595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_10267_ genblk2\[4\].wave_shpr.div.acc\[4\] genblk2\[4\].wave_shpr.div.b1\[4\] VGND
+ VGND VPWR VPWR _04579_ sky130_fd_sc_hd__or2b_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ clknet_leaf_113_clk _00382_ net128 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12006_ genblk2\[11\].wave_shpr.div.b1\[12\] _01494_ _05802_ VGND VGND VPWR VPWR
+ _05808_ sky130_fd_sc_hd__mux2_1
XANTENNA__11537__B genblk1\[8\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10198_ _04406_ _04526_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12908_ clknet_leaf_36_clk _00239_ net103 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07151__A2 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12839_ clknet_leaf_65_clk _00172_ net197 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06366__B _01309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06360_ _01303_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__clkbuf_4
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11786__A2 _02203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06291_ genblk1\[0\].osc.clkdiv_C.cnt\[13\] _01240_ _01243_ _01244_ _01252_ VGND
+ VGND VPWR VPWR _01253_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08030_ genblk2\[6\].wave_shpr.div.fin_quo\[3\] _02736_ VGND VGND VPWR VPWR _02737_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07478__A _02204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06382__A _01229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold803 genblk2\[3\].wave_shpr.div.acc\[25\] VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 genblk2\[0\].wave_shpr.div.acc\[21\] VGND VGND VPWR VPWR net1032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 genblk2\[6\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold836 genblk2\[2\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net1054 sky130_fd_sc_hd__buf_1
XFILLER_0_101_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold847 sig_norm.acc\[3\] VGND VGND VPWR VPWR net1065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 genblk2\[6\].wave_shpr.div.acc\[25\] VGND VGND VPWR VPWR net1076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 genblk2\[10\].wave_shpr.div.acc\[21\] VGND VGND VPWR VPWR net1087 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ genblk2\[3\].wave_shpr.div.acc\[3\] genblk2\[3\].wave_shpr.div.b1\[3\] VGND
+ VGND VPWR VPWR _04377_ sky130_fd_sc_hd__or2b_1
XFILLER_0_40_787 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08932_ _03625_ _03591_ sig_norm.acc\[11\] VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__mux2_1
X_08863_ _03525_ _03568_ _03569_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07914__A1 genblk1\[8\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07914__B2 _01489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07814_ _02308_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08794_ _03491_ _03495_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07745_ genblk1\[1\].osc.clkdiv_C.cnt\[12\] _01344_ _01337_ genblk1\[1\].osc.clkdiv_C.cnt\[11\]
+ _02451_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_79_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07678__B1 _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07676_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _01190_ _01992_ genblk1\[10\].osc.clkdiv_C.cnt\[4\]
+ _02371_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__a221o_1
X_09415_ _03967_ _03977_ _03978_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_149_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06627_ _01523_ _01530_ _01531_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_137_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10079__A _03833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09346_ genblk2\[0\].wave_shpr.div.acc\[25\] genblk2\[0\].wave_shpr.div.acc\[24\]
+ genblk2\[0\].wave_shpr.div.acc\[26\] _03802_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__nor4_1
XFILLER_0_47_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06558_ genblk1\[2\].osc.clkdiv_C.cnt\[12\] genblk1\[2\].osc.clkdiv_C.cnt\[11\] _01468_
+ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09277_ _03835_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__clkbuf_4
X_06489_ genblk1\[2\].osc.clkdiv_C.cnt\[15\] _01414_ _01210_ VGND VGND VPWR VPWR _01415_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08228_ _02933_ _02934_ genblk2\[4\].wave_shpr.div.fin_quo\[6\] _02362_ VGND VGND
+ VPWR VPWR _02935_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07850__B1 _02316_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08159_ _01489_ genblk1\[3\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11170_ _05226_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06956__A2 _01311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10121_ net296 _04461_ _04462_ net451 _04471_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__a221o_1
X_10052_ genblk2\[4\].wave_shpr.div.b1\[5\] _01870_ _04238_ VGND VGND VPWR VPWR _04435_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13742_ clknet_leaf_46_clk _01053_ net121 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10954_ _04676_ _01729_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06467__A genblk1\[1\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07133__A2 _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13673_ clknet_leaf_40_clk _00986_ net117 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13757__RESET_B net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10885_ _05026_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12624_ clknet_leaf_19_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[9\] net109 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08094__B1 _01498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12555_ clknet_leaf_55_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[12\] net175 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11506_ genblk2\[8\].wave_shpr.div.quo\[8\] _05447_ _05446_ net404 VGND VGND VPWR
+ VPWR _00803_ sky130_fd_sc_hd__a22o_1
X_12486_ clknet_leaf_107_clk _00048_ net151 VGND VGND VPWR VPWR sig_norm.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10991__A3 _05023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11437_ genblk2\[8\].wave_shpr.div.acc\[23\] _05412_ VGND VGND VPWR VPWR _05413_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11368_ _05249_ _05245_ genblk2\[7\].wave_shpr.div.i\[0\] VGND VGND VPWR VPWR _05349_
+ sky130_fd_sc_hd__mux2_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ clknet_leaf_13_clk _00432_ net53 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11548__A _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10319_ _04627_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _05197_ _05173_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__or2b_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ clknet_leaf_126_clk _00365_ net66 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07761__A _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09452__S _00007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10598__S _00015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07530_ _02247_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07461_ _02155_ _02192_ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09200_ _03828_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06412_ _01226_ _01355_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__or2_2
XANTENNA__11208__A1 _03726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07392_ _02141_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11759__A2 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06343_ genblk1\[0\].osc.clkdiv_C.cnt\[12\] _01290_ _01292_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__o21a_1
X_09131_ genblk2\[0\].wave_shpr.div.b1\[8\] genblk2\[0\].wave_shpr.div.acc\[8\] VGND
+ VGND VPWR VPWR _03779_ sky130_fd_sc_hd__and2b_1
XFILLER_0_115_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06824__B genblk1\[5\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09062_ _03701_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__buf_4
X_06274_ genblk1\[0\].osc.clkdiv_C.cnt\[3\] _01227_ _01235_ genblk1\[0\].osc.clkdiv_C.cnt\[1\]
+ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13080__RESET_B net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08013_ genblk1\[6\].osc.clkdiv_C.cnt\[5\] _01367_ _02716_ _02718_ _02719_ VGND VGND
+ VPWR VPWR _02720_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold600 genblk2\[6\].wave_shpr.div.acc\[15\] VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 genblk2\[1\].wave_shpr.div.acc\[4\] VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold622 genblk2\[0\].wave_shpr.div.acc\[15\] VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 genblk1\[4\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 genblk2\[3\].wave_shpr.div.acc\[14\] VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold655 genblk2\[7\].wave_shpr.div.acc\[23\] VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold666 genblk2\[9\].wave_shpr.div.acc\[10\] VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 genblk2\[2\].wave_shpr.div.acc\[9\] VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 genblk2\[10\].wave_shpr.div.acc\[23\] VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ net282 _04359_ _04360_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__a21oi_1
Xhold699 genblk2\[8\].wave_shpr.div.acc\[11\] VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08915_ _03614_ _03615_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__nand2_1
X_09895_ net830 _04282_ _04289_ _04311_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__a22o_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _03484_ _03485_ _03497_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__o21ba_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08560__A1 genblk2\[8\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07671__A _01308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08777_ _03465_ _03482_ _03333_ _03483_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ _01342_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07659_ net3 _02364_ _02365_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__nand3_2
XFILLER_0_94_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10670_ _02182_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09329_ _03838_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10958__B1 _05055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12340_ _03833_ _02080_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12271_ _05996_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11222_ genblk2\[7\].wave_shpr.div.quo\[5\] _05246_ _05250_ net661 VGND VGND VPWR
+ VPWR _00716_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11153_ _05049_ genblk2\[7\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR _05213_
+ sky130_fd_sc_hd__and2_1
X_10104_ _04455_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__buf_2
X_11084_ _05149_ _05021_ genblk2\[6\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR
+ _05151_ sky130_fd_sc_hd__mux2_1
X_10035_ genblk2\[3\].wave_shpr.div.fin_quo\[4\] genblk2\[3\].wave_shpr.div.quo\[3\]
+ _04422_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10211__S _04507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11986_ genblk2\[11\].wave_shpr.div.b1\[2\] _01811_ _05433_ VGND VGND VPWR VPWR _05798_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09500__B1 _03733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13725_ clknet_leaf_97_clk net403 net166 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10937_ _05054_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__buf_4
XFILLER_0_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13656_ clknet_leaf_44_clk _00969_ net116 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10661__A2 _04853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10868_ genblk2\[6\].wave_shpr.div.b1\[15\] genblk2\[6\].wave_shpr.div.acc\[15\]
+ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12607_ clknet_leaf_22_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[10\] net94 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_143_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12138__S _05865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13587_ clknet_leaf_73_clk _00902_ net215 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10799_ _04949_ _04950_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12538_ clknet_leaf_63_clk _00090_ net190 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10413__A2 _04651_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12469_ clknet_leaf_33_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[3\] net101 VGND VGND
+ VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.cnt\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06961_ _01432_ _01221_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__nand2_2
X_08700_ _03405_ _03404_ _03401_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__a21bo_1
X_09680_ genblk2\[2\].wave_shpr.div.acc\[13\] genblk2\[2\].wave_shpr.div.b1\[13\]
+ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__or2b_1
X_06892_ genblk1\[6\].osc.clkdiv_C.cnt\[14\] _01675_ _01666_ genblk1\[6\].osc.clkdiv_C.cnt\[13\]
+ _01745_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__o221ai_2
XANTENNA__09182__S _03722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08542__A1 genblk2\[7\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08631_ _03336_ _03337_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08562_ _02676_ _02679_ _02680_ genblk2\[7\].wave_shpr.div.fin_quo\[0\] VGND VGND
+ VPWR VPWR _03269_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07513_ _02232_ PWM.final_sample_in\[3\] VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08493_ _03196_ _03199_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout38 net44 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_4
X_07444_ genblk2\[5\].wave_shpr.div.i\[1\] _02179_ genblk2\[5\].wave_shpr.div.i\[4\]
+ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__or3b_1
XFILLER_0_18_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13261__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout49 net50 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09211__A _03833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10357__A _03708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07375_ genblk1\[11\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09114_ genblk2\[0\].wave_shpr.div.b1\[1\] genblk2\[0\].wave_shpr.div.acc\[1\] VGND
+ VGND VPWR VPWR _03762_ sky130_fd_sc_hd__or2b_1
XFILLER_0_60_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06326_ genblk1\[0\].osc.clkdiv_C.cnt\[6\] _01279_ VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09270__A2 _03804_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06257_ genblk1\[0\].osc.clkdiv_C.cnt\[10\] _01184_ _01206_ _01218_ VGND VGND VPWR
+ VPWR _01219_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09045_ net1238 _01991_ _03708_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09558__B1 _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06188_ _01158_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__clkbuf_4
Xhold430 genblk2\[2\].wave_shpr.div.acc\[20\] VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 genblk2\[6\].wave_shpr.div.acc\[23\] VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11365__B1 _05248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold452 genblk2\[7\].wave_shpr.div.quo\[12\] VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 _00475_ VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold474 genblk2\[5\].wave_shpr.div.b1\[2\] VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 genblk2\[8\].wave_shpr.div.b1\[16\] VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 genblk2\[4\].wave_shpr.div.quo\[24\] VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07584__A2 _01234_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09947_ genblk2\[2\].wave_shpr.div.acc\[24\] _04212_ genblk2\[2\].wave_shpr.div.acc\[25\]
+ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__o21ai_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ net836 _04282_ _04289_ _04298_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__a22o_1
Xhold1130 genblk2\[2\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net1348 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout69_A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08829_ _03533_ _03535_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10340__A1 _03714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10340__B2 _03727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _05593_ _05681_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__xnor2_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13510_ clknet_leaf_80_clk _00827_ net205 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ net888 _04886_ _04890_ _04893_ VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13441_ clknet_leaf_95_clk _00760_ net162 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10653_ _04854_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13372_ clknet_leaf_115_clk _00691_ net140 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10584_ _04649_ genblk2\[5\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR _04812_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_2_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12323_ net351 _06014_ _06015_ net489 _06019_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12254_ _05987_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11205_ _03831_ net722 _03728_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__a21bo_1
X_12185_ net289 _05923_ _03855_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07575__A2 _01925_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09791__A _03833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11136_ _05174_ _05194_ _05195_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__a21o_1
X_11067_ _05017_ net21 genblk2\[6\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR _05140_
+ sky130_fd_sc_hd__o21ai_1
X_10018_ _04361_ _04412_ _04413_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__a21o_1
XANTENNA__11545__B genblk1\[8\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10331__A1 _01304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_137_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_137_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08827__A2 _02592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11969_ _05789_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10095__B1 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13708_ clknet_leaf_36_clk _01019_ net104 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09031__A _02155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11485__B1_N _03728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13639_ clknet_leaf_94_clk _00952_ net159 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07160_ genblk1\[9\].osc.clkdiv_C.cnt\[2\] genblk1\[9\].osc.clkdiv_C.cnt\[1\] genblk1\[9\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06111_ net364 net338 VGND VGND VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.next_cnt\[1\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07091_ genblk1\[8\].osc.clkdiv_C.cnt\[7\] _01897_ genblk1\[8\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout206 net209 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_4
Xfanout217 net218 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__buf_2
X_09801_ net719 _04248_ _04252_ net812 VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07993_ genblk1\[6\].osc.clkdiv_C.cnt\[10\] _01484_ _01519_ genblk1\[6\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__o22a_1
X_09732_ genblk2\[2\].wave_shpr.div.acc\[23\] _04211_ VGND VGND VPWR VPWR _04212_
+ sky130_fd_sc_hd__or2_2
X_06944_ net1146 _01781_ _01784_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__12311__A2 _03947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08748__C _02365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09206__A _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09663_ _04147_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__clkbuf_1
X_06875_ genblk1\[6\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__inv_2
X_08614_ genblk2\[4\].wave_shpr.div.fin_quo\[0\] _02932_ genblk2\[4\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__a21oi_1
X_09594_ _03986_ _03963_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__or2b_1
XFILLER_0_89_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ _02604_ _03248_ _03250_ _03247_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__a22o_1
XANTENNA__08279__B1 _02223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_128_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_128_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__12075__B2 _05813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08476_ _02932_ _02840_ genblk2\[4\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR
+ _03183_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07427_ genblk2\[3\].wave_shpr.div.i\[1\] _02166_ genblk2\[3\].wave_shpr.div.i\[4\]
+ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__or3b_1
XFILLER_0_135_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10087__A _04455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07358_ _02115_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06309_ _01268_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07289_ genblk1\[10\].osc.clkdiv_C.cnt\[14\] genblk1\[10\].osc.clkdiv_C.cnt\[13\]
+ _02053_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09028_ _03698_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__inv_2
XANTENNA__12452__D net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold260 genblk2\[9\].wave_shpr.div.b1\[13\] VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 genblk2\[11\].wave_shpr.div.quo\[14\] VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 genblk2\[5\].wave_shpr.div.quo\[11\] VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09951__A0 _04250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold293 genblk2\[1\].wave_shpr.div.quo\[14\] VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08506__B2 _02468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12302__A2 _06009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12941_ clknet_leaf_111_clk _00270_ net136 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06517__B1 _01442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12872_ clknet_leaf_134_clk _00203_ net59 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _05585_ _05668_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__xnor2_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_119_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _05464_ genblk1\[9\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__and2_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _04818_ _04819_ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__nor2_2
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11685_ genblk2\[9\].wave_shpr.div.b1\[2\] genblk2\[9\].wave_shpr.div.acc\[2\] VGND
+ VGND VPWR VPWR _05577_ sky130_fd_sc_hd__and2b_1
XFILLER_0_102_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13424_ clknet_leaf_87_clk _00743_ net179 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10636_ _04845_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09234__A2 _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13355_ clknet_leaf_4_clk _00676_ net45 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10567_ _04773_ _04793_ _04794_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12306_ net358 _06009_ _06010_ net397 VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13286_ clknet_leaf_118_clk _00607_ net137 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10498_ genblk2\[4\].wave_shpr.div.acc\[18\] _04738_ VGND VGND VPWR VPWR _04739_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12237_ genblk2\[11\].wave_shpr.div.b1\[17\] genblk2\[11\].wave_shpr.div.acc\[17\]
+ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__and2b_1
X_12168_ _05785_ _05899_ _05912_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07753__B _02459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11119_ _05177_ _05178_ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__nand2_1
X_12099_ genblk2\[10\].wave_shpr.div.acc\[6\] _05861_ _05787_ VGND VGND VPWR VPWR
+ _05862_ sky130_fd_sc_hd__mux2_1
Xinput6 pb[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06508__B1 _01432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11501__B1 _05446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06369__B _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06660_ net1237 _01549_ _01552_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09460__S _00007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07720__A2 _01309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06591_ genblk1\[3\].osc.clkdiv_C.cnt\[2\] _01496_ _01498_ genblk1\[3\].osc.clkdiv_C.cnt\[14\]
+ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08330_ _02682_ _03035_ _03036_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06385__A _01326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08261_ _02966_ _02965_ VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__and2b_1
XFILLER_0_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07212_ _01308_ genblk1\[10\].osc.clkdiv_C.cnt\[2\] _01214_ _01993_ genblk1\[10\].osc.clkdiv_C.cnt\[17\]
+ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__a221o_1
X_08192_ _02897_ _02898_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09225__A2 _03836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07143_ genblk1\[9\].osc.clkdiv_C.cnt\[3\] _01514_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07074_ _01879_ _01889_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10354__B _01242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07976_ genblk2\[7\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__inv_2
X_09715_ genblk2\[2\].wave_shpr.div.b1\[11\] genblk2\[2\].wave_shpr.div.acc\[11\]
+ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__and2b_1
XANTENNA__12296__A1 _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06927_ genblk1\[6\].osc.clkdiv_C.cnt\[8\] genblk1\[6\].osc.clkdiv_C.cnt\[7\] _01770_
+ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__and3_1
X_09646_ genblk2\[1\].wave_shpr.div.acc\[20\] _04133_ _04136_ VGND VGND VPWR VPWR
+ _04137_ sky130_fd_sc_hd__a21o_1
X_06858_ genblk1\[5\].osc.clkdiv_C.cnt\[13\] genblk1\[5\].osc.clkdiv_C.cnt\[12\] _01714_
+ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__and3_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _03978_ _03967_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__nor2_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06789_ genblk1\[5\].osc.clkdiv_C.cnt\[2\] _01660_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12297__A _03942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _03230_ _03234_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08267__A3 _02350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08459_ genblk2\[6\].wave_shpr.div.fin_quo\[3\] _02734_ _02736_ _02261_ VGND VGND
+ VPWR VPWR _03166_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11470_ net1187 _01946_ _05237_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10421_ genblk2\[4\].wave_shpr.div.acc\[0\] _00012_ _04679_ net643 _04680_ VGND VGND
+ VPWR VPWR _00485_ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13140_ clknet_leaf_115_clk _00465_ net133 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10352_ net1279 _04643_ _04637_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13071_ clknet_leaf_24_clk _00398_ net92 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10283_ _04576_ _04593_ _04594_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__a21o_1
X_12022_ _05815_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__buf_4
XANTENNA__07950__A2 _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12924_ clknet_leaf_35_clk _00255_ net105 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_88_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09280__S _03804_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12855_ clknet_leaf_91_clk _00186_ net146 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ net1006 _05652_ _05653_ _05656_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__a22o_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ clknet_leaf_43_clk _00119_ net124 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _05621_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__clkbuf_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11668_ genblk2\[9\].wave_shpr.div.acc\[11\] genblk2\[9\].wave_shpr.div.b1\[11\]
+ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13407_ clknet_leaf_90_clk _00726_ net144 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10619_ _04835_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07748__B _01576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11599_ net909 _05507_ _05484_ _05510_ VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07769__A2 _01256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13338_ clknet_leaf_8_clk _00659_ net50 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13188__D _00015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13269_ clknet_leaf_1_clk _00592_ net41 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10525__A1 _04655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07830_ _02461_ _02463_ genblk2\[1\].wave_shpr.div.fin_quo\[4\] VGND VGND VPWR VPWR
+ _02537_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07761_ _02467_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__clkbuf_4
X_09500_ _03732_ net369 _03733_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__o21a_1
X_06712_ _01601_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[0\] sky130_fd_sc_hd__clkbuf_1
X_07692_ genblk1\[10\].osc.clkdiv_C.cnt\[11\] _02011_ VGND VGND VPWR VPWR _02399_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09190__S _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09431_ _03959_ _03993_ _03994_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06643_ net1145 _01538_ _01541_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09362_ _03802_ _03923_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__nor2_1
X_06574_ _01452_ _01482_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__nor2_1
X_08313_ _02406_ _02404_ _02408_ _02525_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__o31a_1
XFILLER_0_75_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09293_ genblk2\[0\].wave_shpr.div.acc\[5\] _03882_ _03804_ VGND VGND VPWR VPWR _03883_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08244_ _02947_ _02948_ _02949_ _02950_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08175_ _02872_ _02881_ _02877_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07126_ genblk1\[9\].osc.clkdiv_C.cnt\[5\] _01925_ _01855_ genblk1\[9\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07057_ genblk1\[8\].osc.clkdiv_C.cnt\[14\] _01246_ genblk1\[8\].osc.clkdiv_C.cnt\[17\]
+ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_2_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07959_ genblk1\[7\].osc.clkdiv_C.cnt\[10\] _01311_ _01925_ genblk1\[7\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__a22o_1
Xmax_cap24 net1353 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
X_10970_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__and2_1
XANTENNA__07145__B1 _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09629_ _04123_ _04001_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12640_ clknet_leaf_15_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[7\] net73 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12571_ clknet_leaf_28_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[10\] net89 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_50_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_136_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11522_ net237 _05454_ _05449_ net312 _05457_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__a221o_1
XFILLER_0_150_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11453_ _05423_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10404_ genblk2\[4\].wave_shpr.div.quo\[19\] _04661_ _04663_ net255 _04670_ VGND
+ VGND VPWR VPWR _00478_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11384_ genblk2\[8\].wave_shpr.div.acc\[15\] genblk2\[8\].wave_shpr.div.b1\[15\]
+ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13123_ clknet_leaf_124_clk _00448_ net77 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_10335_ _04635_ VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__clkbuf_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ clknet_leaf_113_clk net815 net128 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10266_ genblk2\[4\].wave_shpr.div.b1\[4\] genblk2\[4\].wave_shpr.div.acc\[4\] VGND
+ VGND VPWR VPWR _04578_ sky130_fd_sc_hd__or2b_1
X_12005_ _05807_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__clkbuf_1
X_10197_ _04407_ _04364_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__or2b_1
XFILLER_0_88_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12907_ clknet_leaf_36_clk _00238_ net102 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12838_ clknet_leaf_65_clk _00171_ net196 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12769_ clknet_leaf_93_clk _00102_ net148 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08100__A2 _02805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06290_ genblk1\[0\].osc.clkdiv_C.cnt\[11\] _01251_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold804 genblk2\[9\].wave_shpr.div.acc\[2\] VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 genblk2\[0\].wave_shpr.div.acc\[4\] VGND VGND VPWR VPWR net1033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold826 genblk2\[11\].wave_shpr.div.acc\[1\] VGND VGND VPWR VPWR net1044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 genblk2\[3\].wave_shpr.div.acc\[20\] VGND VGND VPWR VPWR net1055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold848 genblk2\[0\].wave_shpr.div.acc\[1\] VGND VGND VPWR VPWR net1066 sky130_fd_sc_hd__dlygate4sd3_1
X_09980_ _04374_ _04375_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold859 genblk1\[3\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR net1077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07494__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08931_ net1141 _02260_ _03626_ _03574_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08862_ _03136_ _03224_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08102__B _01574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07813_ _02424_ _02471_ _02519_ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__nor3_2
X_08793_ _03484_ _03498_ _03395_ _03499_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__o211a_1
XANTENNA__11744__A _03693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07744_ genblk1\[1\].osc.clkdiv_C.cnt\[13\] _02425_ _01344_ genblk1\[1\].osc.clkdiv_C.cnt\[12\]
+ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__o22ai_2
XANTENNA__07127__B1 _01923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09081__B1_N _03717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07675_ _02369_ _02370_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09414_ genblk2\[1\].wave_shpr.div.b1\[4\] genblk2\[1\].wave_shpr.div.acc\[4\] VGND
+ VGND VPWR VPWR _03978_ sky130_fd_sc_hd__and2b_1
XFILLER_0_149_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06626_ genblk1\[3\].osc.clkdiv_C.cnt\[3\] _01528_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09345_ net604 _03903_ _03910_ _03922_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06557_ net1213 _01468_ _01471_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__07669__A _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09276_ _03839_ _03867_ _03869_ _03841_ net1139 VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06488_ genblk1\[2\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08227_ genblk2\[4\].wave_shpr.div.fin_quo\[5\] _02932_ _02842_ _02316_ VGND VGND
+ VPWR VPWR _02934_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08158_ genblk1\[3\].osc.clkdiv_C.cnt\[7\] _01483_ _01858_ _01486_ _02864_ VGND VGND
+ VPWR VPWR _02865_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07109_ _01886_ _01912_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__nor2_1
X_08089_ genblk2\[5\].wave_shpr.div.fin_quo\[7\] _02309_ _02795_ _02527_ VGND VGND
+ VPWR VPWR _02796_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10120_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_99_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08158__A2 _01483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10051_ _04434_ VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12938__RESET_B net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09658__A2 _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13741_ clknet_leaf_46_clk _01052_ net121 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10953_ net344 _05057_ _05055_ net477 _05060_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13672_ clknet_leaf_40_clk _00985_ net117 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10884_ genblk2\[6\].wave_shpr.div.fin_quo\[2\] net1338 _00017_ VGND VGND VPWR VPWR
+ _05026_ sky130_fd_sc_hd__mux2_1
X_12623_ clknet_leaf_16_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[8\] net74 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06892__A2 _01675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12554_ clknet_leaf_55_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[11\] net175 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11505_ _05441_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12485_ clknet_leaf_106_clk _00047_ net151 VGND VGND VPWR VPWR sig_norm.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09794__A _04247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11436_ genblk2\[8\].wave_shpr.div.acc\[22\] _05411_ VGND VGND VPWR VPWR _05412_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_80_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08397__A2 _01209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11367_ net381 _05251_ _05248_ _05348_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13106_ clknet_leaf_12_clk _00431_ net52 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10318_ genblk2\[4\].wave_shpr.div.fin_quo\[3\] genblk2\[4\].wave_shpr.div.quo\[2\]
+ _00013_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__mux2_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ net1009 _05279_ _05283_ _05297_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__a22o_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ clknet_leaf_125_clk _00364_ net72 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10249_ genblk2\[3\].wave_shpr.div.i\[3\] _02168_ _04560_ VGND VGND VPWR VPWR _04563_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_119_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10900__A1 _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_62_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10664__B1 _04857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07460_ genblk2\[7\].wave_shpr.div.busy _02191_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06411_ _01354_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__buf_4
XFILLER_0_57_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06883__A2 _01484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07391_ _02091_ _02138_ _02140_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_146_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10416__B1 _04654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09130_ _03756_ _03776_ _03777_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06342_ _01268_ _01291_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__nor2_1
XANTENNA__07489__A _02147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06393__A _01336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09061_ _01193_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__inv_2
X_06273_ _01231_ _01234_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__nor2_4
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12169__B1 _05816_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_120_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08012_ genblk1\[6\].osc.clkdiv_C.cnt\[4\] _01747_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__or2_1
XANTENNA__07134__A1_N genblk1\[9\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold601 genblk2\[6\].wave_shpr.div.acc\[6\] VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold612 genblk2\[2\].wave_shpr.div.acc\[11\] VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold623 genblk2\[11\].wave_shpr.div.acc\[6\] VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 genblk2\[7\].wave_shpr.div.acc\[12\] VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 genblk2\[5\].wave_shpr.div.acc\[6\] VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout101_A net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold656 genblk2\[1\].wave_shpr.div.acc\[20\] VGND VGND VPWR VPWR net874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 genblk2\[5\].wave_shpr.div.acc\[5\] VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold678 genblk2\[5\].wave_shpr.div.acc\[19\] VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ net282 _04359_ _03855_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_135_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold689 genblk2\[6\].wave_shpr.div.acc\[5\] VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ sig_norm.acc\[5\] _03611_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__nand2_1
X_09894_ genblk2\[2\].wave_shpr.div.acc\[10\] _04310_ _04301_ VGND VGND VPWR VPWR
+ _04311_ sky130_fd_sc_hd__mux2_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12341__B1 _03941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _03533_ _03535_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__and2b_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08560__A2 _02362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08776_ _03298_ _03332_ _03331_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__a21bo_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07727_ genblk1\[1\].osc.clkdiv_C.cnt\[5\] _02433_ _01305_ genblk1\[1\].osc.clkdiv_C.cnt\[4\]
+ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__o22ai_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06287__B _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07658_ _02312_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06323__A1 genblk1\[0\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06609_ genblk1\[3\].osc.clkdiv_C.cnt\[4\] _01514_ _01513_ genblk1\[3\].osc.clkdiv_C.cnt\[3\]
+ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07589_ _02282_ _02286_ _02292_ _02295_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__o31a_1
X_09328_ net913 _03903_ _03877_ _03909_ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__a22o_1
XANTENNA__09812__A2 _04253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09259_ _03853_ genblk1\[0\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09025__B1 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12270_ net1267 _04229_ _05994_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__mux2_1
XANTENNA__11907__B1 _03855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11221_ genblk2\[7\].wave_shpr.div.quo\[4\] _05246_ _05250_ net331 VGND VGND VPWR
+ VPWR _00715_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07587__B1 _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11152_ _05166_ _05210_ _05211_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__a21oi_1
X_10103_ _04451_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__buf_2
X_11083_ genblk2\[6\].wave_shpr.div.acc\[24\] _05057_ _05126_ _05150_ VGND VGND VPWR
+ VPWR _00677_ sky130_fd_sc_hd__a22o_1
X_10034_ _04426_ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10894__A0 genblk2\[6\].wave_shpr.div.fin_quo\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11985_ _05797_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09500__A1 _03732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10936_ _05053_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__clkbuf_4
X_13724_ clknet_leaf_96_clk _01035_ net160 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13655_ clknet_leaf_41_clk _00968_ net116 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10867_ _04969_ _05009_ _05010_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12606_ clknet_leaf_22_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[9\] net92 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_2
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13586_ clknet_leaf_72_clk _00901_ net215 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09264__B1 _03838_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10798_ genblk2\[5\].wave_shpr.div.acc\[23\] _04818_ VGND VGND VPWR VPWR _04950_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09803__A2 _04248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07102__A genblk1\[8\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12537_ clknet_leaf_41_clk _00089_ net123 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12468_ clknet_leaf_34_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[2\] net99 VGND VGND
+ VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.cnt\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11419_ _05365_ _05393_ _05394_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__a21o_1
X_12399_ net949 _06039_ _06040_ _06071_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__a22o_1
XANTENNA__07042__A2 _01436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06250__B1 _01210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06960_ genblk1\[7\].osc.clkdiv_C.cnt\[10\] genblk1\[7\].osc.clkdiv_C.cnt\[0\] _01514_
+ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__and3b_1
Xclkbuf_leaf_3_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_16
X_06891_ genblk1\[6\].osc.clkdiv_C.cnt\[13\] _01666_ _01484_ genblk1\[6\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08542__A2 _02526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08630_ genblk2\[6\].wave_shpr.div.fin_quo\[2\] _02733_ _02735_ _02261_ VGND VGND
+ VPWR VPWR _03337_ sky130_fd_sc_hd__a31o_1
XANTENNA__07491__B _02152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08561_ _03266_ _03267_ _02604_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07512_ PWM.counter\[3\] VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__inv_2
X_08492_ _03197_ _03198_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07443_ genblk2\[5\].wave_shpr.div.i\[2\] genblk2\[5\].wave_shpr.div.i\[3\] genblk2\[5\].wave_shpr.div.i\[0\]
+ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__nand3b_1
Xfanout39 net44 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13648__RESET_B net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout149_A net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07374_ net1269 _02123_ _02127_ _02092_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[10\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10357__B _01441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09113_ genblk2\[0\].wave_shpr.div.b1\[2\] VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06325_ genblk1\[0\].osc.clkdiv_C.cnt\[6\] _01279_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09044_ _03710_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06256_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] _01210_ _01212_ _01217_ VGND VGND VPWR
+ VPWR _01218_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_142_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold420 _00472_ VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__dlygate4sd3_1
X_06187_ _01157_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__inv_2
Xhold431 genblk2\[9\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold442 genblk2\[8\].wave_shpr.div.quo\[20\] VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold453 genblk2\[6\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold464 genblk2\[10\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 genblk2\[7\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08136__C_N _02837_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold486 genblk2\[8\].wave_shpr.div.acc\[23\] VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold497 genblk2\[0\].wave_shpr.div.acc\[0\] VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__dlygate4sd3_1
X_09946_ net1094 _04253_ _04251_ _04348_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__a22o_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ genblk2\[2\].wave_shpr.div.acc\[6\] _04297_ _04214_ VGND VGND VPWR VPWR _04298_
+ sky130_fd_sc_hd__mux2_1
Xhold1120 genblk2\[6\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net1338 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 genblk2\[6\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net1349 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ net8 _02744_ _03534_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__and3_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ genblk2\[5\].wave_shpr.div.fin_quo\[0\] _02467_ _02791_ VGND VGND VPWR VPWR
+ _03466_ sky130_fd_sc_hd__a21o_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ net304 _05628_ _05629_ net485 _05634_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__a221o_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ genblk2\[5\].wave_shpr.div.acc\[3\] _04892_ _04821_ VGND VGND VPWR VPWR _04893_
+ sky130_fd_sc_hd__mux2_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13440_ clknet_leaf_95_clk _00759_ net162 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10652_ _02170_ genblk2\[5\].wave_shpr.div.busy _02180_ VGND VGND VPWR VPWR _04854_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_76_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08018__A _01739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13371_ clknet_leaf_117_clk _00690_ net140 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10583_ _04765_ _04809_ _04810_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12322_ _05835_ genblk1\[11\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__and2_1
XANTENNA__10800__B1 _04858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11379__A _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12253_ genblk2\[11\].wave_shpr.div.fin_quo\[4\] genblk2\[11\].wave_shpr.div.quo\[3\]
+ _00005_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11204_ _03727_ _01490_ _03687_ net1005 VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12184_ _03690_ _05922_ _05923_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__nor3_1
XFILLER_0_102_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11135_ genblk2\[7\].wave_shpr.div.b1\[7\] genblk2\[7\].wave_shpr.div.acc\[7\] VGND
+ VGND VPWR VPWR _05195_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12305__B1 _06010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11066_ _05018_ net21 VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__or2_1
X_10017_ genblk2\[3\].wave_shpr.div.b1\[17\] genblk2\[3\].wave_shpr.div.acc\[17\]
+ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11968_ genblk2\[10\].wave_shpr.div.fin_quo\[1\] genblk2\[10\].wave_shpr.div.quo\[0\]
+ _00003_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10095__A1 genblk2\[3\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10095__B2 net401 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13707_ clknet_leaf_37_clk _01018_ net104 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10919_ _05044_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11899_ _03839_ _05723_ _05724_ _03841_ net1106 VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__a32o_1
XFILLER_0_67_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13638_ clknet_leaf_94_clk net221 net159 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09237__B1 _03839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13569_ clknet_leaf_55_clk _00884_ net182 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07799__B1 _01577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09458__S _00007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06110_ net338 VGND VGND VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.next_cnt\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07090_ genblk1\[8\].osc.clkdiv_C.cnt\[8\] genblk1\[8\].osc.clkdiv_C.cnt\[7\] _01897_
+ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09800_ net812 _04248_ _04252_ net1054 VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__a22o_1
Xfanout207 net208 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_4
Xfanout218 net16 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_4
X_07992_ genblk2\[6\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12623__RESET_B net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09731_ genblk2\[2\].wave_shpr.div.acc\[22\] genblk2\[2\].wave_shpr.div.acc\[21\]
+ genblk2\[2\].wave_shpr.div.acc\[20\] _04210_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__or4_1
X_06943_ net28 _01783_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__nor2_1
X_09662_ _04046_ _04042_ genblk2\[1\].wave_shpr.div.i\[0\] VGND VGND VPWR VPWR _04147_
+ sky130_fd_sc_hd__mux2_1
X_06874_ genblk1\[6\].osc.clkdiv_C.cnt\[16\] _01578_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__xnor2_1
X_08613_ _03318_ _03319_ _02797_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__a21bo_1
X_09593_ net827 _04076_ _04080_ _04096_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08544_ _02603_ _03247_ _03248_ _03250_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__and4_1
XFILLER_0_49_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11283__B1 _05283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08475_ _03180_ _03181_ _02797_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__o21a_1
XANTENNA__06829__A2 genblk1\[5\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07426_ genblk2\[3\].wave_shpr.div.i\[2\] genblk2\[3\].wave_shpr.div.i\[3\] genblk2\[3\].wave_shpr.div.i\[0\]
+ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_92_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07357_ _02092_ _02113_ _02114_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06308_ net1089 _01269_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07288_ genblk1\[10\].osc.clkdiv_C.cnt\[13\] _02053_ genblk1\[10\].osc.clkdiv_C.cnt\[14\]
+ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09027_ genblk2\[9\].wave_shpr.div.i\[1\] genblk2\[9\].wave_shpr.div.i\[0\] genblk2\[9\].wave_shpr.div.i\[2\]
+ genblk2\[9\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06239_ _01200_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09559__B_N _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold250 _01044_ VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold261 genblk2\[11\].wave_shpr.div.quo\[9\] VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold272 genblk2\[3\].wave_shpr.div.quo\[23\] VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _00555_ VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09951__A1 _04247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold294 _00222_ VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__dlygate4sd3_1
X_09929_ _04336_ _04337_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__nand2_1
X_12940_ clknet_leaf_110_clk _00269_ net136 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ clknet_leaf_134_clk _00202_ net59 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11822_ _05586_ _05564_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__or2b_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ net526 _05623_ _05624_ net1085 VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__a22o_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _03819_ net493 _00014_ genblk2\[5\].wave_shpr.div.acc\[0\] _04879_ VGND VGND
+ VPWR VPWR _00569_ sky130_fd_sc_hd__o221a_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _05572_ genblk2\[9\].wave_shpr.div.acc\[1\] _05575_ VGND VGND VPWR VPWR _05576_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13423_ clknet_leaf_87_clk _00742_ net179 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10635_ genblk2\[6\].wave_shpr.div.b1\[10\] _04844_ _04834_ VGND VGND VPWR VPWR _04845_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13354_ clknet_leaf_4_clk _00675_ net45 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10566_ genblk2\[5\].wave_shpr.div.b1\[7\] genblk2\[5\].wave_shpr.div.acc\[7\] VGND
+ VGND VPWR VPWR _04794_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12305_ net397 _06009_ _06010_ net731 VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__a22o_1
X_13285_ clknet_leaf_117_clk _00606_ net137 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_10497_ _04617_ _04622_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__nand2b_1
X_12236_ _05810_ genblk2\[11\].wave_shpr.div.acc\[16\] _05973_ VGND VGND VPWR VPWR
+ _05974_ sky130_fd_sc_hd__a21o_1
X_12167_ genblk2\[10\].wave_shpr.div.acc\[24\] _05784_ VGND VGND VPWR VPWR _05912_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07953__B1 _02656_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11118_ genblk2\[7\].wave_shpr.div.acc\[4\] genblk2\[7\].wave_shpr.div.b1\[4\] VGND
+ VGND VPWR VPWR _05178_ sky130_fd_sc_hd__or2b_1
X_12098_ _05757_ _05860_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__xnor2_1
X_11049_ _05054_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__06508__A1 _01201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput7 pb[1] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_4
XFILLER_0_79_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09741__S _00009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06590_ _01497_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06385__B _01328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08260_ _02965_ _02966_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07211_ genblk1\[10\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08191_ _02697_ _02747_ _02896_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07142_ genblk1\[9\].osc.clkdiv_C.cnt\[3\] _01514_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07073_ _01862_ _01885_ _01888_ _01889_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[1\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08105__B _01192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10651__A _02183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07944__B1 _01514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09217__A _03838_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07975_ _02681_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__buf_2
X_09714_ _04163_ _04192_ _04193_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__a21o_1
X_06926_ _01761_ _01772_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09645_ _04007_ _04129_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__nor2_1
X_06857_ genblk1\[5\].osc.clkdiv_C.cnt\[12\] _01714_ _01716_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__o21a_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ net829 _04076_ _04080_ _04083_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__a22o_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06788_ _01179_ _01262_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__nor2_1
XANTENNA__06576__A _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10059__A1 _01263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _03232_ _03233_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08458_ _02734_ _02736_ genblk2\[6\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR
+ _03165_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07409_ _02149_ _02153_ genblk2\[0\].wave_shpr.div.busy VGND VGND VPWR VPWR _02154_
+ sky130_fd_sc_hd__and3b_1
X_08389_ _03086_ _03095_ genblk1\[2\].osc.clkdiv_C.cnt\[7\] _02011_ VGND VGND VPWR
+ VPWR _03096_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_107_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10420_ _03719_ genblk1\[4\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07200__A genblk1\[9\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10351_ _01355_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10782__A2 _04880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13070_ clknet_leaf_24_clk _00397_ net92 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10282_ genblk2\[4\].wave_shpr.div.b1\[6\] genblk2\[4\].wave_shpr.div.acc\[6\] VGND
+ VGND VPWR VPWR _04594_ sky130_fd_sc_hd__and2b_1
X_12021_ genblk2\[10\].wave_shpr.div.quo\[0\] _05813_ _05787_ _05816_ VGND VGND VPWR
+ VPWR _00949_ sky130_fd_sc_hd__a22o_1
XANTENNA__07935__B1 _02223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12923_ clknet_leaf_35_clk _00254_ net105 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ clknet_leaf_119_clk _00185_ net139 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ genblk2\[9\].wave_shpr.div.acc\[2\] _05655_ _05613_ VGND VGND VPWR VPWR _05656_
+ sky130_fd_sc_hd__mux2_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ clknet_leaf_41_clk _00118_ net123 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09797__A _04250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11736_ net1259 genblk2\[9\].wave_shpr.div.quo\[6\] _00023_ VGND VGND VPWR VPWR _05621_
+ sky130_fd_sc_hd__mux2_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11667_ genblk2\[9\].wave_shpr.div.acc\[12\] genblk2\[9\].wave_shpr.div.b1\[12\]
+ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__or2b_1
XFILLER_0_142_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13406_ clknet_leaf_90_clk _00725_ net144 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10618_ genblk2\[6\].wave_shpr.div.b1\[3\] _01758_ _04834_ VGND VGND VPWR VPWR _04835_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07218__A2 _01246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11598_ genblk2\[8\].wave_shpr.div.acc\[11\] _05509_ _05493_ VGND VGND VPWR VPWR
+ _05510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06426__B1 _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10549_ genblk2\[5\].wave_shpr.div.acc\[4\] genblk2\[5\].wave_shpr.div.b1\[4\] VGND
+ VGND VPWR VPWR _04777_ sky130_fd_sc_hd__or2b_1
XFILLER_0_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13337_ clknet_leaf_8_clk _00658_ net49 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13268_ clknet_leaf_1_clk _00591_ net44 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12219_ genblk2\[11\].wave_shpr.div.b1\[8\] genblk2\[11\].wave_shpr.div.acc\[8\]
+ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__and2b_1
X_13199_ clknet_leaf_114_clk _00522_ net134 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11722__A1 _05613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07760_ _02362_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__clkbuf_4
X_06711_ genblk1\[4\].osc.clkdiv_C.cnt\[0\] _01600_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__and2b_1
X_07691_ _02373_ _02384_ _02385_ _02397_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__a211o_1
X_09430_ genblk2\[1\].wave_shpr.div.b1\[12\] genblk2\[1\].wave_shpr.div.acc\[12\]
+ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__and2b_1
X_06642_ _01523_ _01540_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06396__A _01238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09361_ net653 _03841_ _03910_ _03933_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__a22o_1
X_06573_ genblk1\[2\].osc.clkdiv_C.cnt\[17\] _01480_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08312_ _02404_ _02408_ _02406_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09292_ _03881_ _03772_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08243_ _02225_ _02682_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout131_A net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08174_ _02873_ _02874_ _02871_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07125_ _01924_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07056_ genblk1\[8\].osc.clkdiv_C.cnt\[3\] _01498_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10381__A _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07958_ _02655_ _02663_ _02664_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06909_ genblk1\[6\].osc.clkdiv_C.cnt\[1\] net837 VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11477__B1 _04233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07889_ genblk2\[0\].wave_shpr.div.fin_quo\[6\] _02595_ VGND VGND VPWR VPWR _02596_
+ sky130_fd_sc_hd__xnor2_1
Xmax_cap36 _01423_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_2
X_09628_ _04002_ _03955_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout44_A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09559_ net588 _04046_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__or2b_1
XFILLER_0_65_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12570_ clknet_leaf_28_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[9\] net90 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09842__B1 _04250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12441__A2 _03947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07999__A3 _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11521_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11452_ genblk2\[8\].wave_shpr.div.fin_quo\[5\] genblk2\[8\].wave_shpr.div.quo\[4\]
+ _00021_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10403_ _04058_ _01588_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__nor2_1
X_11383_ _05243_ genblk2\[8\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR _05359_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_21_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13122_ clknet_leaf_136_clk _00447_ net43 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10334_ net1212 _01240_ _04440_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__mux2_1
XANTENNA__07865__A _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07620__A2 _01430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ clknet_leaf_113_clk _00380_ net128 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10265_ genblk2\[4\].wave_shpr.div.acc\[5\] genblk2\[4\].wave_shpr.div.b1\[5\] VGND
+ VGND VPWR VPWR _04577_ sky130_fd_sc_hd__or2b_1
X_12004_ genblk2\[11\].wave_shpr.div.b1\[11\] _01500_ _05802_ VGND VGND VPWR VPWR
+ _05807_ sky130_fd_sc_hd__mux2_1
X_10196_ net862 _04518_ _04522_ _04525_ VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08581__B1 _02525_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12906_ clknet_leaf_36_clk _00237_ net104 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07687__A2 _02011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10140__B1 _04457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ clknet_leaf_65_clk _00170_ net196 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ clknet_leaf_93_clk _00101_ net148 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11719_ genblk2\[9\].wave_shpr.div.acc\[23\] genblk2\[9\].wave_shpr.div.acc\[25\]
+ genblk2\[9\].wave_shpr.div.acc\[24\] genblk2\[9\].wave_shpr.div.acc\[26\] VGND VGND
+ VPWR VPWR _05611_ sky130_fd_sc_hd__or4_2
XFILLER_0_25_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12699_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[12\] net172 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_116_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput10 pb[4] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold805 genblk2\[9\].wave_shpr.div.acc\[19\] VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold816 genblk2\[2\].wave_shpr.div.acc\[21\] VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09466__S _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold827 genblk2\[9\].wave_shpr.div.acc\[25\] VGND VGND VPWR VPWR net1045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 genblk2\[5\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net1056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 genblk2\[3\].wave_shpr.div.acc\[1\] VGND VGND VPWR VPWR net1067 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07611__A2 _01437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08930_ sig_norm.acc\[10\] _03590_ _03625_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__a21o_1
XANTENNA__09364__A2 _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08861_ _03565_ _03567_ _03519_ _03523_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__or4_1
X_07812_ _02509_ _02516_ _02518_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__o21ai_1
X_08792_ _03384_ _03394_ _03393_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07743_ _02440_ _02443_ _02449_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07127__A1 genblk1\[9\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07674_ _02378_ _02376_ _02380_ _02375_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__or4b_1
XANTENNA__10131__B1 _04455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06625_ genblk1\[3\].osc.clkdiv_C.cnt\[3\] _01528_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__and2_1
X_09413_ _03968_ _03975_ _03976_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06886__B1 _01739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11760__A _02203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09344_ genblk2\[0\].wave_shpr.div.acc\[17\] _03921_ _03803_ VGND VGND VPWR VPWR
+ _03922_ sky130_fd_sc_hd__mux2_1
X_06556_ _01451_ _01470_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12890__RESET_B net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09275_ _03804_ _03868_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06487_ genblk1\[2\].osc.clkdiv_C.cnt\[12\] _01411_ _01412_ _01183_ VGND VGND VPWR
+ VPWR _01413_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07669__B _01440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08226_ _02932_ _02842_ genblk2\[4\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR
+ _02933_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08157_ genblk1\[3\].osc.clkdiv_C.cnt\[14\] _01361_ _02851_ _02863_ VGND VGND VPWR
+ VPWR _02864_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07108_ genblk1\[8\].osc.clkdiv_C.cnt\[14\] _01910_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__and2_1
X_08088_ genblk2\[5\].wave_shpr.div.fin_quo\[6\] _02794_ VGND VGND VPWR VPWR _02795_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07039_ genblk1\[8\].osc.clkdiv_C.cnt\[5\] _01487_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10050_ net1188 _01248_ _04238_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10050__S _04238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13740_ clknet_leaf_46_clk _01051_ net121 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10952_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__and2_1
X_13671_ clknet_leaf_40_clk _00984_ net118 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10883_ _05025_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12622_ clknet_leaf_17_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[7\] net83 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12553_ clknet_leaf_55_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[10\] net176 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08094__A2 _01359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11504_ net404 _05442_ _05446_ net676 VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12484_ clknet_leaf_107_clk _00046_ net151 VGND VGND VPWR VPWR sig_norm.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09043__A1 _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11435_ genblk2\[8\].wave_shpr.div.acc\[21\] _05410_ VGND VGND VPWR VPWR _05411_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11366_ genblk2\[7\].wave_shpr.div.acc\[25\] _05346_ VGND VGND VPWR VPWR _05348_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13766__RESET_B net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10317_ _04626_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__clkbuf_1
X_13105_ clknet_leaf_12_clk _00430_ net52 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11297_ net893 _05296_ _05222_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__mux2_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ clknet_leaf_123_clk _00363_ net76 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10248_ _00010_ _04560_ net1148 VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10179_ _04399_ _04368_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__or2b_1
XANTENNA__06580__A2 _01344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10664__B2 net308 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06410_ _01178_ _01176_ freq_div.state\[0\] VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__mux2_2
XFILLER_0_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07390_ _02139_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__inv_2
XANTENNA__09806__B1 _04252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09050__A _03708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06341_ genblk1\[0\].osc.clkdiv_C.cnt\[12\] _01290_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06393__B _01226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09060_ _03720_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06272_ _01229_ _01230_ _01233_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__a21o_2
XFILLER_0_4_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08011_ genblk1\[6\].osc.clkdiv_C.cnt\[5\] _01367_ _01747_ genblk1\[6\].osc.clkdiv_C.cnt\[4\]
+ _02717_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold602 genblk2\[3\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__S _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold613 PWM.counter\[2\] VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold624 genblk2\[4\].wave_shpr.div.acc\[4\] VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold635 _00749_ VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 genblk2\[8\].wave_shpr.div.b1\[0\] VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 genblk2\[11\].wave_shpr.div.acc\[12\] VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold668 genblk2\[9\].wave_shpr.div.acc\[4\] VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 genblk2\[11\].wave_shpr.div.acc\[15\] VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ _03690_ _04358_ _04359_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__nor3_1
X_08913_ sig_norm.acc\[5\] _03611_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__or2_1
X_09893_ _04192_ _04309_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__xnor2_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _03540_ _03550_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__nand2_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08775_ _03465_ _03480_ _03481_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__nor3_2
XFILLER_0_79_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ _01342_ _01241_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__nor2_4
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07657_ net136 VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06608_ genblk1\[3\].osc.clkdiv_C.cnt\[9\] _01210_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__xnor2_1
X_07588_ _02284_ _02283_ _02293_ _02294_ _02285_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__o311a_1
XFILLER_0_137_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09327_ genblk2\[0\].wave_shpr.div.acc\[13\] _03908_ _03889_ VGND VGND VPWR VPWR
+ _03909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06539_ genblk1\[2\].osc.clkdiv_C.cnt\[4\] _01456_ genblk1\[2\].osc.clkdiv_C.cnt\[5\]
+ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08076__A2 _01678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09258_ net265 _03845_ _03847_ net636 _03858_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08209_ _02910_ _02914_ _02915_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__a21oi_1
X_09189_ _03701_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11206__B1_N _03717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11220_ net331 _05246_ _05250_ net693 VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__a22o_1
XANTENNA__07036__B1 _01578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11151_ genblk2\[7\].wave_shpr.div.b1\[15\] genblk2\[7\].wave_shpr.div.acc\[15\]
+ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__and2b_1
X_10102_ net525 _04457_ _04454_ net631 _04460_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11082_ genblk2\[6\].wave_shpr.div.acc\[23\] _05020_ _05149_ VGND VGND VPWR VPWR
+ _05150_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10033_ genblk2\[3\].wave_shpr.div.fin_quo\[3\] genblk2\[3\].wave_shpr.div.quo\[2\]
+ _04422_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11984_ genblk2\[11\].wave_shpr.div.b1\[1\] _03813_ _05433_ VGND VGND VPWR VPWR _05797_
+ sky130_fd_sc_hd__mux2_1
X_13723_ clknet_leaf_96_clk net431 net160 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10935_ _02152_ genblk2\[6\].wave_shpr.div.busy _02186_ VGND VGND VPWR VPWR _05053_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_105_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13654_ clknet_leaf_41_clk _00967_ net116 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10866_ genblk2\[6\].wave_shpr.div.b1\[14\] genblk2\[6\].wave_shpr.div.acc\[14\]
+ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__and2b_1
XANTENNA__06494__A _01242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12605_ clknet_leaf_22_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[8\] net94 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_4
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13585_ clknet_leaf_76_clk _00900_ net207 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10797_ genblk2\[5\].wave_shpr.div.acc\[23\] _04818_ VGND VGND VPWR VPWR _04949_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12536_ clknet_leaf_44_clk _00088_ net123 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07102__B genblk1\[8\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12467_ clknet_leaf_33_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[1\] net99 VGND VGND
+ VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.cnt\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11418_ genblk2\[8\].wave_shpr.div.b1\[10\] genblk2\[8\].wave_shpr.div.acc\[10\]
+ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__and2b_1
X_12398_ genblk2\[11\].wave_shpr.div.acc\[12\] _06070_ _06055_ VGND VGND VPWR VPWR
+ _06071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11349_ genblk2\[7\].wave_shpr.div.acc\[20\] _05334_ VGND VGND VPWR VPWR _05336_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07042__A3 _01855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06250__B2 genblk1\[0\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13019_ clknet_leaf_123_clk _00346_ net76 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_06890_ genblk1\[6\].osc.clkdiv_C.cnt\[12\] _01519_ _01739_ genblk1\[6\].osc.clkdiv_C.cnt\[8\]
+ _01743_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__a221o_1
XANTENNA__06669__A _01349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08560_ genblk2\[8\].wave_shpr.div.fin_quo\[2\] _02362_ _02636_ VGND VGND VPWR VPWR
+ _03267_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07511_ _02230_ PWM.final_sample_in\[5\] VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__and2_1
XANTENNA__10637__A1 _04223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08491_ _03066_ _03070_ VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06305__A2 _01227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07442_ _02178_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07373_ genblk1\[11\].osc.clkdiv_C.cnt\[10\] _02123_ VGND VGND VPWR VPWR _02127_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08058__A2 _01172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09112_ genblk2\[0\].wave_shpr.div.acc\[3\] genblk2\[0\].wave_shpr.div.b1\[3\] VGND
+ VGND VPWR VPWR _03760_ sky130_fd_sc_hd__or2b_1
XANTENNA__10357__C _01367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06324_ _01269_ _01279_ _01280_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_72_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09043_ genblk2\[0\].wave_shpr.div.b1\[2\] _02002_ _03708_ VGND VGND VPWR VPWR _03710_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06255_ genblk1\[0\].osc.clkdiv_C.cnt\[0\] _01211_ _01215_ genblk1\[0\].osc.clkdiv_C.cnt\[4\]
+ _01216_ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__a221o_1
XANTENNA__07947__B _01574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold410 genblk2\[7\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09558__A2 _04042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06186_ _01155_ _01150_ _01156_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__a21oi_4
Xhold421 genblk2\[2\].wave_shpr.div.quo\[22\] VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold432 _00867_ VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07569__A1 genblk1\[9\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold443 genblk2\[7\].wave_shpr.div.quo\[4\] VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold454 genblk2\[4\].wave_shpr.div.quo\[10\] VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold465 _00953_ VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold476 genblk2\[4\].wave_shpr.div.acc\[20\] VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 genblk2\[10\].wave_shpr.div.acc\[20\] VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06241__A1 _01201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold498 genblk2\[2\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09945_ _04346_ _04212_ genblk2\[2\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR
+ _04348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _04184_ _04296_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__xnor2_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 genblk2\[9\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net1328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06579__A _01172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 sig_norm.quo\[4\] VGND VGND VPWR VPWR net1339 sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ genblk2\[2\].wave_shpr.div.fin_quo\[0\] _02592_ _02468_ genblk2\[2\].wave_shpr.div.fin_quo\[1\]
+ _03114_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__a221o_1
XANTENNA__07741__A1 genblk1\[1\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07741__B2 genblk1\[1\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _03258_ _03452_ _03464_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__and3_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10628__A1 _01189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _02415_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__buf_2
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _03366_ _03376_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _04786_ _04891_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__xnor2_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07203__A genblk1\[9\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10651_ _02183_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10582_ genblk2\[5\].wave_shpr.div.b1\[15\] genblk2\[5\].wave_shpr.div.acc\[15\]
+ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__and2b_1
X_13370_ clknet_leaf_116_clk _00689_ net140 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12321_ genblk2\[11\].wave_shpr.div.quo\[14\] _06014_ _06015_ net342 _06018_ VGND
+ VGND VPWR VPWR _01047_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12252_ _05986_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11203_ _03726_ _01869_ _05242_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12183_ genblk2\[10\].wave_shpr.div.i\[3\] _02207_ _05920_ VGND VGND VPWR VPWR _05923_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_102_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_61_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11134_ _05175_ _05192_ _05193_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__a21o_1
XANTENNA__12305__A1 net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11065_ genblk2\[6\].wave_shpr.div.acc\[25\] genblk2\[6\].wave_shpr.div.acc\[24\]
+ genblk2\[6\].wave_shpr.div.acc\[26\] _05021_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__nor4_1
X_10016_ _04362_ _04410_ _04411_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__o21bai_1
XANTENNA_clkbuf_leaf_76_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12069__B1 _05815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11967_ _05788_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10095__A2 _04452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13706_ clknet_leaf_37_clk _01017_ net114 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10918_ net1253 net34 _05042_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11898_ genblk2\[0\].wave_shpr.div.i\[1\] genblk2\[0\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _05724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_134_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13637_ clknet_leaf_93_clk _00950_ net159 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10849_ _04978_ _04991_ _04992_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09739__S _00009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13568_ clknet_leaf_55_clk _00883_ net176 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07799__A1 genblk1\[0\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12519_ clknet_leaf_104_clk PWM.next_counter\[3\] net157 VGND VGND VPWR VPWR PWM.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13499_ clknet_leaf_86_clk _00816_ net179 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout208 net209 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_4
X_07991_ _02604_ _02645_ _02648_ _02696_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__a22o_1
XANTENNA__07971__A1 _01201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_09730_ genblk2\[2\].wave_shpr.div.acc\[19\] _04209_ VGND VGND VPWR VPWR _04210_
+ sky130_fd_sc_hd__or2_1
X_06942_ genblk1\[6\].osc.clkdiv_C.cnt\[13\] genblk1\[6\].osc.clkdiv_C.cnt\[12\] _01779_
+ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__and3_1
X_09661_ net1107 _04048_ _04045_ _04146_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__a22o_1
X_06873_ genblk1\[6\].osc.clkdiv_C.cnt\[10\] _01726_ genblk1\[6\].osc.clkdiv_C.cnt\[14\]
+ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__o21bai_1
X_08612_ genblk2\[5\].wave_shpr.div.fin_quo\[2\] _02521_ _02791_ VGND VGND VPWR VPWR
+ _03319_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12663__RESET_B net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09592_ genblk2\[1\].wave_shpr.div.acc\[7\] _04094_ _04095_ VGND VGND VPWR VPWR _04096_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08543_ _02225_ _02682_ _03249_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__a21o_1
XANTENNA__10649__A _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08474_ genblk2\[5\].wave_shpr.div.fin_quo\[4\] _02308_ _02791_ VGND VGND VPWR VPWR
+ _03181_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07425_ _02165_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07356_ genblk1\[11\].osc.clkdiv_C.cnt\[6\] _02108_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06307_ _01268_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__clkbuf_4
X_07287_ genblk1\[10\].osc.clkdiv_C.cnt\[13\] _02053_ _02055_ VGND VGND VPWR VPWR
+ genblk1\[10\].osc.clkdiv_C.next_cnt\[13\] sky130_fd_sc_hd__o21a_1
XFILLER_0_33_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09026_ genblk2\[9\].wave_shpr.div.i\[1\] genblk2\[9\].wave_shpr.div.i\[0\] genblk2\[9\].wave_shpr.div.i\[2\]
+ genblk2\[9\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__a31o_1
X_06238_ _01181_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__buf_6
XFILLER_0_32_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06169_ _01129_ _01140_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__nor2_1
Xhold240 _00305_ VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 genblk2\[8\].wave_shpr.div.quo\[10\] VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 genblk2\[2\].wave_shpr.div.quo\[14\] VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _00399_ VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold284 genblk2\[8\].wave_shpr.div.quo\[16\] VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold295 genblk2\[9\].wave_shpr.div.quo\[18\] VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__dlygate4sd3_1
X_09928_ _04208_ net22 genblk2\[2\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR _04337_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__12299__B1 _06010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout74_A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07562__A2_N _01799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09859_ _04176_ _04283_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__xnor2_1
X_12870_ clknet_leaf_134_clk _00201_ net59 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ net984 _05652_ _05653_ _05667_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__a22o_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ genblk2\[9\].wave_shpr.div.quo\[7\] _05623_ _05624_ net267 VGND VGND VPWR
+ VPWR _00872_ sky130_fd_sc_hd__a22o_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ genblk2\[5\].wave_shpr.div.acc_next\[0\] _04856_ VGND VGND VPWR VPWR _04879_
+ sky130_fd_sc_hd__or2b_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ genblk2\[9\].wave_shpr.div.b1\[0\] _05573_ _05574_ VGND VGND VPWR VPWR _05575_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13422_ clknet_leaf_92_clk _00741_ net149 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10634_ _01742_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13353_ clknet_leaf_4_clk _00674_ net45 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10565_ _04774_ _04791_ _04792_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12304_ net731 _06009_ _06010_ net767 VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13284_ clknet_leaf_117_clk _00605_ net137 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_10496_ net1074 _04715_ _04722_ _04737_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12235_ _05926_ _05972_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__and2b_1
X_12166_ _05816_ _05910_ _05911_ _05818_ net536 VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__a32o_1
X_11117_ genblk2\[7\].wave_shpr.div.b1\[4\] genblk2\[7\].wave_shpr.div.acc\[4\] VGND
+ VGND VPWR VPWR _05177_ sky130_fd_sc_hd__or2b_1
X_12097_ genblk2\[10\].wave_shpr.div.b1\[6\] genblk2\[10\].wave_shpr.div.acc\[6\]
+ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__xor2_1
XANTENNA__12014__A _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07108__A genblk1\[8\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11048_ net921 _05119_ _05093_ _05125_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__a22o_1
Xinput8 pb[2] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_127_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12999_ clknet_leaf_132_clk _00328_ net60 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11265__A1 _03819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09469__S _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07210_ _01359_ _01224_ _01241_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08190_ _02697_ _02747_ _02896_ VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_859 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07141_ _01935_ _01939_ _01940_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07072_ genblk1\[8\].osc.clkdiv_C.cnt\[1\] genblk1\[8\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01889_ sky130_fd_sc_hd__nand2_2
XFILLER_0_140_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08105__C _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12844__RESET_B net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10143__S _04420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07974_ _02676_ _02679_ _02680_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__o21ai_2
X_09713_ genblk2\[2\].wave_shpr.div.b1\[10\] genblk2\[2\].wave_shpr.div.acc\[10\]
+ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__and2b_1
X_06925_ genblk1\[6\].osc.clkdiv_C.cnt\[7\] _01770_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09644_ net874 _04109_ _04113_ _04135_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06856_ _01693_ _01715_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__nor2_1
XANTENNA__10700__B1 _04856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09575_ genblk2\[1\].wave_shpr.div.acc\[3\] _04082_ _04011_ VGND VGND VPWR VPWR _04083_
+ sky130_fd_sc_hd__mux2_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06787_ genblk1\[5\].osc.clkdiv_C.cnt\[10\] _01658_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__xor2_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06576__B _01302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _03227_ _03229_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08457_ _02648_ _03162_ _03158_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_147_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13632__RESET_B net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07408_ _02152_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__buf_6
XFILLER_0_80_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08388_ _03090_ _03092_ _03094_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07339_ _02100_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07200__B genblk1\[9\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10350_ _04642_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06986__A2 _01227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09009_ _03684_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__clkbuf_1
X_10281_ _04577_ _04591_ _04592_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12020_ _05815_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__buf_4
X_12922_ clknet_leaf_35_clk _00253_ net105 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12853_ clknet_leaf_119_clk _00184_ net139 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _05576_ _05654_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__xnor2_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ clknet_leaf_40_clk _00117_ net123 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08982__A _01097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11735_ _05620_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__clkbuf_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08663__A2 _02521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09289__S _03804_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11666_ genblk2\[9\].wave_shpr.div.acc\[13\] genblk2\[9\].wave_shpr.div.b1\[13\]
+ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__or2b_1
X_13405_ clknet_leaf_90_clk _00724_ net143 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10617_ _03701_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11597_ _05395_ _05508_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06426__A1 _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13336_ clknet_leaf_6_clk _00657_ net48 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06426__B2 genblk1\[1\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10548_ genblk2\[5\].wave_shpr.div.b1\[4\] genblk2\[5\].wave_shpr.div.acc\[4\] VGND
+ VGND VPWR VPWR _04776_ sky130_fd_sc_hd__or2b_1
XFILLER_0_122_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13267_ clknet_leaf_1_clk _00590_ net38 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10479_ genblk2\[4\].wave_shpr.div.acc\[13\] _04724_ _04704_ VGND VGND VPWR VPWR
+ _04725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12218_ _05935_ _05954_ _05955_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__a21o_1
X_13198_ clknet_leaf_114_clk _00521_ net134 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12149_ _05782_ _05899_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10930__B1 _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09752__S _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06710_ _01599_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__buf_2
XFILLER_0_79_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11486__A1 _03831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07690_ _02003_ _01991_ _02393_ _02396_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_79_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06641_ genblk1\[3\].osc.clkdiv_C.cnt\[9\] _01538_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__and2_1
XANTENNA__06396__B _01262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09360_ genblk2\[0\].wave_shpr.div.acc\[22\] _03931_ VGND VGND VPWR VPWR _03933_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06572_ genblk1\[2\].osc.clkdiv_C.cnt\[16\] _01478_ _01481_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[16\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08311_ _02366_ _03017_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09291_ _03773_ _03758_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__or2b_1
XANTENNA__09199__S _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08242_ genblk2\[7\].wave_shpr.div.fin_quo\[6\] _02309_ VGND VGND VPWR VPWR _02949_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07862__B1 _02361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08173_ _01486_ _01858_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07124_ _01336_ _01355_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06968__A2 _01801_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07055_ genblk1\[8\].osc.clkdiv_C.cnt\[8\] _01430_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07917__A1 genblk1\[8\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06601__A2_N _01507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07957_ genblk1\[7\].osc.clkdiv_C.cnt\[8\] _01920_ _01947_ genblk1\[7\].osc.clkdiv_C.cnt\[7\]
+ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__a22o_1
XANTENNA__11493__A _02152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06908_ net837 _01761_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11477__A1 _03704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07888_ _02513_ genblk2\[0\].wave_shpr.div.fin_quo\[5\] _02510_ VGND VGND VPWR VPWR
+ _02595_ sky130_fd_sc_hd__or3b_1
Xmax_cap26 _03602_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
XANTENNA__07145__A2 _01514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_cap37 _01320_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_4
X_09627_ net774 _04109_ _04113_ _04122_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__a22o_1
X_06839_ genblk1\[5\].osc.clkdiv_C.cnt\[6\] _01703_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__and2_1
X_09558_ net588 _04042_ _04046_ genblk2\[1\].wave_shpr.div.quo\[24\] _04070_ VGND
+ VGND VPWR VPWR _00232_ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08509_ _03208_ _03215_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09489_ _01420_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11520_ net312 _05454_ _05449_ net482 _05456_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11451_ _05422_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10048__S _04238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10402_ net255 _04661_ _04663_ net531 _04669_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11382_ genblk2\[8\].wave_shpr.div.acc\[17\] genblk2\[8\].wave_shpr.div.b1\[17\]
+ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13121_ clknet_leaf_136_clk _00446_ net43 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10333_ _03714_ net692 _01262_ _03705_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__o22a_1
XANTENNA__12263__S _05802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13052_ clknet_leaf_113_clk net780 net131 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10264_ genblk2\[4\].wave_shpr.div.acc\[6\] genblk2\[4\].wave_shpr.div.b1\[6\] VGND
+ VGND VPWR VPWR _04576_ sky130_fd_sc_hd__or2b_1
XANTENNA__12762__SET_B net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12003_ _05806_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__clkbuf_1
X_10195_ genblk2\[3\].wave_shpr.div.acc\[13\] _04524_ _04507_ VGND VGND VPWR VPWR
+ _04525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11468__A1 _01811_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12905_ clknet_leaf_37_clk _00236_ net104 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10140__A1 _04454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12836_ clknet_leaf_64_clk _00169_ net196 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07105__B genblk1\[8\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output18_A net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12767_ clknet_leaf_93_clk _00100_ net148 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11718_ genblk2\[9\].wave_shpr.div.acc\[22\] _05609_ VGND VGND VPWR VPWR _05610_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_126_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12698_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[11\] net172 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_127_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11649_ _05545_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__clkbuf_1
Xinput11 pb[5] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09747__S _00009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold806 genblk2\[4\].wave_shpr.div.acc\[10\] VGND VGND VPWR VPWR net1024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 genblk2\[10\].wave_shpr.div.acc\[9\] VGND VGND VPWR VPWR net1035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13319_ clknet_leaf_26_clk net621 net87 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold828 genblk2\[9\].wave_shpr.div.acc\[12\] VGND VGND VPWR VPWR net1046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold839 genblk2\[3\].wave_shpr.div.acc\[3\] VGND VGND VPWR VPWR net1057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08860_ _03507_ _03451_ _03506_ _03566_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__or4_1
X_07811_ _02517_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__buf_2
XANTENNA__08572__B2 _02362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08791_ _03484_ _03485_ _03497_ VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__nor3b_2
X_07742_ _02445_ _02446_ _02447_ _02448_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_74_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09521__B1 _04045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07673_ genblk1\[10\].osc.clkdiv_C.cnt\[0\] _02001_ _02379_ _02013_ genblk1\[10\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__a32o_1
XANTENNA__13295__RESET_B net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09412_ genblk2\[1\].wave_shpr.div.b1\[3\] genblk2\[1\].wave_shpr.div.acc\[3\] VGND
+ VGND VPWR VPWR _03976_ sky130_fd_sc_hd__and2b_1
X_06624_ _01523_ _01528_ _01529_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09343_ _03796_ _03920_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__xnor2_1
X_06555_ genblk1\[2\].osc.clkdiv_C.cnt\[11\] _01468_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09274_ _03764_ _03765_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06486_ genblk1\[2\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08225_ _02837_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__buf_2
XFILLER_0_118_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08156_ genblk1\[3\].osc.clkdiv_C.cnt\[14\] _01361_ _01576_ genblk1\[3\].osc.clkdiv_C.cnt\[15\]
+ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_31_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07063__A1 _01441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07107_ net1182 _01908_ _01911_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_141_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08087_ genblk2\[5\].wave_shpr.div.fin_quo\[5\] _02789_ _02793_ VGND VGND VPWR VPWR
+ _02794_ sky130_fd_sc_hd__or3b_1
XFILLER_0_30_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07038_ _01436_ _01855_ genblk1\[8\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _01856_
+ sky130_fd_sc_hd__a21oi_1
X_08989_ sig_norm.quo\[9\] _03672_ _01155_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__mux2_1
XANTENNA__10370__B2 _04655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10331__S _03689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09512__B1 _04047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10951_ _04268_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08866__A2 _02248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13670_ clknet_leaf_40_clk _00983_ net117 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10882_ genblk2\[6\].wave_shpr.div.fin_quo\[1\] genblk2\[6\].wave_shpr.div.quo\[0\]
+ _00017_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__mux2_1
X_12621_ clknet_leaf_17_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[6\] net80 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12552_ clknet_leaf_60_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[9\] net186 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08037__A _02364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11503_ net676 _05442_ _05446_ net751 VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12483_ clknet_leaf_108_clk _00045_ net151 VGND VGND VPWR VPWR sig_norm.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11434_ genblk2\[8\].wave_shpr.div.acc\[20\] genblk2\[8\].wave_shpr.div.acc\[18\]
+ genblk2\[8\].wave_shpr.div.acc\[19\] _05409_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__or4_1
XANTENNA__07054__A1 genblk1\[8\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_100_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_100_clk sky130_fd_sc_hd__clkbuf_16
X_11365_ net1053 _05251_ _05248_ _05347_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__a22o_1
X_13104_ clknet_leaf_13_clk _00429_ net52 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_10316_ genblk2\[4\].wave_shpr.div.fin_quo\[2\] genblk2\[4\].wave_shpr.div.quo\[1\]
+ _00013_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06801__B2 _01436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11296_ _05194_ _05295_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__xnor2_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ clknet_leaf_122_clk _00362_ net76 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10247_ _04454_ _04559_ _04561_ _04457_ net725 VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__a32o_1
X_10178_ net790 _04486_ _04490_ _04511_ VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__a22o_1
XANTENNA__12022__A _05815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09503__B1 _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10664__A2 _04853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12819_ clknet_leaf_66_clk _00152_ net196 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08609__A2 _02789_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10416__A2 _04651_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06340_ _01269_ _01289_ _01290_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_151_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12688__RESET_B net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06271_ _01232_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12169__A2 _05818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08010_ genblk1\[6\].osc.clkdiv_C.cnt\[5\] _01365_ genblk1\[6\].osc.clkdiv_C.cnt\[3\]
+ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold603 genblk2\[0\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold614 _01160_ VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold625 _00489_ VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 genblk2\[0\].wave_shpr.div.acc\[3\] VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 genblk2\[1\].wave_shpr.div.acc\[13\] VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11101__A _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold658 genblk2\[11\].wave_shpr.div.acc\[8\] VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ genblk2\[2\].wave_shpr.div.i\[3\] _02163_ _04356_ VGND VGND VPWR VPWR _04359_
+ sky130_fd_sc_hd__and3_1
Xhold669 genblk2\[2\].wave_shpr.div.acc\[6\] VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08912_ net1027 _02260_ _03613_ _03574_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09892_ _04193_ _04163_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__or2b_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12341__A2 _03942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08843_ _03529_ _03547_ _03549_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__and3_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09506__A _02170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout191_A net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10352__A1 _04643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08774_ _03258_ _03452_ _03464_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__a21oi_1
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07725_ genblk1\[1\].osc.clkdiv_C.cnt\[4\] _01305_ _01313_ genblk1\[1\].osc.clkdiv_C.cnt\[3\]
+ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__a22o_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07656_ genblk2\[11\].wave_shpr.div.fin_quo\[7\] _02362_ VGND VGND VPWR VPWR _02363_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06607_ genblk1\[3\].osc.clkdiv_C.cnt\[3\] _01513_ _01514_ genblk1\[3\].osc.clkdiv_C.cnt\[4\]
+ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12078__S _05787_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10387__A _04651_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07587_ genblk1\[9\].osc.clkdiv_C.cnt\[7\] _01234_ _01513_ genblk1\[9\].osc.clkdiv_C.cnt\[6\]
+ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09326_ _03788_ _03907_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06538_ genblk1\[2\].osc.clkdiv_C.cnt\[5\] genblk1\[2\].osc.clkdiv_C.cnt\[4\] _01456_
+ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__and3_1
XANTENNA__07808__B1 _02224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_838 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11080__A2 _05057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09257_ _03853_ genblk1\[0\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__and2_1
X_06469_ genblk1\[1\].osc.clkdiv_C.cnt\[12\] _01398_ _01400_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08208_ _02901_ _02419_ _02905_ _02909_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__and4_1
XFILLER_0_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09188_ _03714_ _03821_ _03705_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11368__A0 _05249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09025__A2 _03694_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07036__A1 genblk1\[8\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08139_ net10 _02364_ _02365_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__and3_2
XFILLER_0_121_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07587__A2 _01234_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11150_ _05167_ _05208_ _05209_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__a21o_1
X_10101_ _04269_ genblk1\[3\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__and2_1
X_11081_ _05021_ _05138_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10032_ _04425_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__clkbuf_1
X_11983_ _03732_ net1007 _05796_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13722_ clknet_leaf_97_clk _01033_ net161 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10934_ _05051_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13653_ clknet_leaf_41_clk net354 net116 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10865_ _04970_ _05007_ _05008_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06494__B _01223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12604_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[7\] net97 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13584_ clknet_leaf_75_clk _00899_ net207 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10796_ net1012 _04858_ _04922_ _04948_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__a22o_1
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12535_ clknet_leaf_45_clk _00087_ net186 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08472__B1 _02526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09297__S _03804_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12466_ clknet_leaf_33_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[0\] net101 VGND VGND
+ VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.cnt\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11417_ _05366_ _05391_ _05392_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__a21o_1
X_12397_ _05964_ _06069_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11348_ net923 _05311_ _05315_ _05335_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__a22o_1
XANTENNA__06250__A2 _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10760__A _04856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11279_ _05249_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__clkbuf_4
X_13018_ clknet_leaf_123_clk _00345_ net76 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10334__A1 _01240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06669__B _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07510_ PWM.counter\[5\] VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10098__B1 _04454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08490_ _03164_ _03169_ _03163_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__a21bo_1
X_07441_ _02175_ _02153_ genblk2\[4\].wave_shpr.div.busy VGND VGND VPWR VPWR _02178_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07372_ _02126_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[9\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__08058__A3 _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09111_ genblk2\[0\].wave_shpr.div.acc\[4\] genblk2\[0\].wave_shpr.div.b1\[4\] VGND
+ VGND VPWR VPWR _03759_ sky130_fd_sc_hd__or2b_1
XFILLER_0_44_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06323_ genblk1\[0\].osc.clkdiv_C.cnt\[4\] _01276_ genblk1\[0\].osc.clkdiv_C.cnt\[5\]
+ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10935__A _02152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12451__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09042_ _03709_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06254_ genblk1\[0\].osc.clkdiv_C.cnt\[4\] _01215_ _01193_ genblk1\[0\].osc.clkdiv_C.cnt\[9\]
+ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_143_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12011__A1 _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold400 _00814_ VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__dlygate4sd3_1
X_06185_ _01152_ _01097_ sig_norm.busy VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__and3b_1
Xhold411 sig_norm.acc\[1\] VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 genblk2\[7\].wave_shpr.div.quo\[13\] VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07569__A2 _01577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold433 genblk2\[10\].wave_shpr.div.b1\[5\] VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _00716_ VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09963__B1 _03855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold455 _00469_ VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 genblk2\[1\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 genblk1\[10\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ genblk2\[2\].wave_shpr.div.acc\[24\] _04253_ _04322_ _04347_ VGND VGND VPWR
+ VPWR _00341_ sky130_fd_sc_hd__a22o_1
Xhold488 genblk2\[7\].wave_shpr.div.acc\[22\] VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 sig_norm.acc\[9\] VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12361__S _05982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _04185_ _04167_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__or2b_1
Xhold1100 genblk2\[7\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net1318 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11522__B1 _05449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06579__B _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 genblk2\[2\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net1329 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 genblk2\[4\].wave_shpr.div.acc\[7\] VGND VGND VPWR VPWR net1340 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ _02575_ _03532_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__xor2_2
XANTENNA__07741__A2 _01337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08757_ _03461_ _03463_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__and2_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10089__B1 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _02225_ _02403_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__and2_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _03384_ _03393_ _03394_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__or3_2
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ _02333_ _02334_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__or2b_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11006__A _05054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10650_ _04852_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09309_ _03780_ _03894_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10581_ _04766_ _04807_ _04808_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12320_ _05835_ genblk1\[11\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10800__A2 _04855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12002__A1 _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12251_ genblk2\[11\].wave_shpr.div.fin_quo\[3\] net402 _00005_ VGND VGND VPWR VPWR
+ _05986_ sky130_fd_sc_hd__mux2_1
X_11202_ _03702_ net1147 VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__nor2_1
X_12182_ _00002_ _05920_ net1153 VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__a21oi_1
X_11133_ genblk2\[7\].wave_shpr.div.b1\[6\] genblk2\[7\].wave_shpr.div.acc\[6\] VGND
+ VGND VPWR VPWR _05193_ sky130_fd_sc_hd__and2b_1
XANTENNA__12305__A2 _06009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11064_ net560 _05119_ _05126_ _05137_ VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__a22o_1
XANTENNA__11513__B1 _05449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09182__A1 _01214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10015_ _04245_ genblk2\[3\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR _04411_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07732__A2 _02433_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11966_ genblk2\[10\].wave_shpr.div.fin_quo\[0\] _05787_ _00003_ VGND VGND VPWR VPWR
+ _05788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10917_ _05043_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__clkbuf_1
X_13705_ clknet_leaf_37_clk _01016_ net113 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11897_ genblk2\[0\].wave_shpr.div.i\[1\] genblk2\[0\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _05723_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13636_ clknet_leaf_68_clk _00949_ net195 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_27_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10848_ genblk2\[6\].wave_shpr.div.b1\[5\] genblk2\[6\].wave_shpr.div.acc\[5\] VGND
+ VGND VPWR VPWR _04992_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13567_ clknet_leaf_55_clk net350 net176 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10779_ genblk2\[5\].wave_shpr.div.acc\[17\] _04936_ _04907_ VGND VGND VPWR VPWR
+ _04937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10755__A _02183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07799__A2 _01349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12518_ clknet_leaf_105_clk PWM.next_counter\[2\] net155 VGND VGND VPWR VPWR PWM.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08225__A _02837_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13498_ clknet_leaf_86_clk _00815_ net178 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12449_ clknet_leaf_106_clk net766 net153 VGND VGND VPWR VPWR sig_norm.i\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09755__S _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11752__B1 _05624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07990_ _02604_ _02645_ _02648_ _02696_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__nand4_2
Xfanout209 net210 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06941_ genblk1\[6\].osc.clkdiv_C.cnt\[12\] _01779_ _01782_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__11504__B1 _05446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09660_ genblk2\[1\].wave_shpr.div.acc\[25\] _04009_ _04145_ VGND VGND VPWR VPWR
+ _04146_ sky130_fd_sc_hd__a21bo_1
X_06872_ _01441_ _01366_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__nor2_1
X_08611_ _03316_ _02223_ _03317_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__or3b_1
XANTENNA__07723__A2 _01323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09591_ _04010_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__buf_4
X_08542_ genblk2\[7\].wave_shpr.div.fin_quo\[0\] _02526_ _02308_ genblk2\[7\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11205__B1_N _03728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08473_ genblk2\[5\].wave_shpr.div.fin_quo\[3\] _03178_ _03179_ VGND VGND VPWR VPWR
+ _03180_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11283__A2 _05279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07424_ _02162_ _02153_ genblk2\[2\].wave_shpr.div.busy VGND VGND VPWR VPWR _02165_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_64_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12632__RESET_B net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07355_ _02112_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10243__B1 _04457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06306_ _01169_ _01185_ _01219_ _01267_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__o211a_2
XFILLER_0_122_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07286_ genblk1\[10\].osc.clkdiv_C.cnt\[13\] _02053_ _02027_ VGND VGND VPWR VPWR
+ _02055_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09025_ _03691_ _03694_ _03695_ _03696_ net1149 VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__a32o_1
X_06237_ genblk1\[0\].osc.clkdiv_C.cnt\[17\] _01197_ _01198_ VGND VGND VPWR VPWR _01199_
+ sky130_fd_sc_hd__a21o_1
Xhold230 genblk2\[1\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06168_ _01133_ _01137_ _01139_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__a21oi_1
Xhold241 genblk2\[5\].wave_shpr.div.quo\[23\] VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 _00806_ VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 genblk2\[9\].wave_shpr.div.quo\[11\] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12091__S _05787_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold274 genblk2\[7\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10604__S _00015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold285 genblk2\[5\].wave_shpr.div.quo\[20\] VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 genblk2\[3\].wave_shpr.div.quo\[15\] VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09927_ _04209_ net22 VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__or2_1
XANTENNA__12299__B2 _05982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09858_ genblk2\[2\].wave_shpr.div.b1\[2\] genblk2\[2\].wave_shpr.div.acc\[2\] VGND
+ VGND VPWR VPWR _04283_ sky130_fd_sc_hd__xor2_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout67_A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08809_ _03513_ _03514_ _03511_ _03515_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__a211o_1
X_09789_ net730 VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__inv_2
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ genblk2\[9\].wave_shpr.div.acc\[6\] _05666_ _05613_ VGND VGND VPWR VPWR _05667_
+ sky130_fd_sc_hd__mux2_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07214__A _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ net267 _05623_ _05624_ net712 VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__a22o_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_80_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ genblk2\[5\].wave_shpr.div.acc_next\[0\] _02183_ _04856_ net324 _04878_ VGND
+ VGND VPWR VPWR _00568_ sky130_fd_sc_hd__a221o_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11682_ genblk2\[9\].wave_shpr.div.b1\[1\] genblk2\[9\].wave_shpr.div.acc\[1\] VGND
+ VGND VPWR VPWR _05574_ sky130_fd_sc_hd__xor2_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13421_ clknet_leaf_92_clk _00740_ net147 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10633_ _04843_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13352_ clknet_leaf_4_clk _00673_ net45 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10564_ genblk2\[5\].wave_shpr.div.b1\[6\] genblk2\[5\].wave_shpr.div.acc\[6\] VGND
+ VGND VPWR VPWR _04792_ sky130_fd_sc_hd__and2b_1
XFILLER_0_140_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12303_ net767 _06009_ _06010_ net776 VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__a22o_1
XANTENNA__11982__B1 _03702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13283_ clknet_leaf_117_clk _00604_ net137 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_10495_ genblk2\[4\].wave_shpr.div.acc\[17\] _04736_ _04622_ VGND VGND VPWR VPWR
+ _04737_ sky130_fd_sc_hd__mux2_1
XANTENNA__09575__S _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12234_ _05927_ _05970_ _05971_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12165_ genblk2\[10\].wave_shpr.div.acc\[22\] _05908_ genblk2\[10\].wave_shpr.div.acc\[23\]
+ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_20_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11116_ genblk2\[7\].wave_shpr.div.acc\[5\] genblk2\[7\].wave_shpr.div.b1\[5\] VGND
+ VGND VPWR VPWR _05176_ sky130_fd_sc_hd__or2b_1
XANTENNA__07953__A2 _01732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12096_ net1241 _05844_ _05850_ _05859_ VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11047_ genblk2\[6\].wave_shpr.div.acc\[13\] _05124_ _05105_ VGND VGND VPWR VPWR
+ _05125_ sky130_fd_sc_hd__mux2_1
Xinput9 pb[3] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12998_ clknet_leaf_131_clk _00327_ net64 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07124__A _01336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08666__B1 _02316_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11949_ _05736_ _05769_ _05770_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13619_ clknet_leaf_68_clk _00932_ net211 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07140_ genblk1\[9\].osc.clkdiv_C.cnt\[6\] _01334_ _01328_ genblk1\[9\].osc.clkdiv_C.cnt\[13\]
+ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_109_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07071_ genblk1\[8\].osc.clkdiv_C.cnt\[1\] genblk1\[8\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01888_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07973_ genblk1\[7\].osc.clkdiv_C.cnt\[16\] genblk1\[7\].osc.clkdiv_C.cnt\[17\] VGND
+ VGND VPWR VPWR _02680_ sky130_fd_sc_hd__nor2_1
X_09712_ _04164_ _04190_ _04191_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__a21o_1
X_06924_ _01761_ _01770_ _01771_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
X_09643_ _04133_ _04134_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__nand2_1
X_06855_ genblk1\[5\].osc.clkdiv_C.cnt\[12\] _01714_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__and2_1
X_09574_ _03975_ _04081_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06786_ _01489_ net37 VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__nand2_2
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _02310_ _03231_ _02314_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__o21a_1
XANTENNA__07034__A genblk1\[8\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_62_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08121__A2 _01439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08456_ _02946_ _03158_ _03162_ VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__or3b_2
XFILLER_0_65_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07407_ genblk2\[0\].wave_shpr.div.start VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__inv_6
XFILLER_0_46_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08387_ genblk1\[2\].osc.clkdiv_C.cnt\[6\] _01433_ _03093_ VGND VGND VPWR VPWR _03094_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10395__A _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06592__B _01437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07338_ _02092_ _02098_ _02099_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07269_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _02041_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09008_ net1132 sig_norm.quo\[5\] _01154_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__mux2_1
XANTENNA__07132__A1_N genblk1\[9\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10280_ genblk2\[4\].wave_shpr.div.b1\[5\] genblk2\[4\].wave_shpr.div.acc\[5\] VGND
+ VGND VPWR VPWR _04592_ sky130_fd_sc_hd__and2b_1
XFILLER_0_103_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10334__S _04440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07209__A _01556_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_133_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12921_ clknet_leaf_35_clk _00252_ net105 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ clknet_leaf_118_clk _00183_ net138 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold915_A genblk1\[0\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06371__B2 genblk1\[1\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _05577_ _05571_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__or2b_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ clknet_leaf_40_clk _00116_ net117 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11734_ genblk2\[9\].wave_shpr.div.fin_quo\[6\] genblk2\[9\].wave_shpr.div.quo\[5\]
+ _00023_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__mux2_1
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11665_ genblk2\[9\].wave_shpr.div.acc\[14\] genblk2\[9\].wave_shpr.div.b1\[14\]
+ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__or2b_1
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10616_ _04833_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__clkbuf_1
X_13404_ clknet_leaf_90_clk net371 net143 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11596_ _05396_ _05364_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__or2b_1
XFILLER_0_51_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13335_ clknet_leaf_6_clk _00656_ net48 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10547_ genblk2\[5\].wave_shpr.div.acc\[5\] genblk2\[5\].wave_shpr.div.b1\[5\] VGND
+ VGND VPWR VPWR _04775_ sky130_fd_sc_hd__or2b_1
XFILLER_0_40_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13266_ clknet_leaf_0_clk _00589_ net38 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10478_ _04607_ _04723_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__xnor2_1
X_12217_ genblk2\[11\].wave_shpr.div.b1\[7\] genblk2\[11\].wave_shpr.div.acc\[7\]
+ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__and2b_1
X_13197_ clknet_leaf_113_clk _00520_ net134 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11183__A1 _04242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12148_ genblk2\[10\].wave_shpr.div.acc\[25\] genblk2\[10\].wave_shpr.div.acc\[26\]
+ _05785_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__nor3_2
XANTENNA__10930__A1 _03726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12079_ net989 _05844_ _05817_ _05846_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__a22o_1
XANTENNA__07139__B1 _01196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06677__B _01565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10694__B1 _04856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06640_ _01523_ _01538_ _01539_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_78_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08639__B1 _02526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06571_ _01451_ _01480_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_44_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_16
X_08310_ _03014_ _03015_ _03016_ _02360_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__o211a_1
X_09290_ net823 _03870_ _03877_ _03880_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07311__B1 _01262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08241_ _02683_ _02682_ _02689_ _02527_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__o31ai_1
XANTENNA__07862__A1 _02525_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08172_ genblk1\[3\].osc.clkdiv_C.cnt\[13\] _01498_ _02867_ VGND VGND VPWR VPWR _02879_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__07301__B _01595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07123_ _01432_ _01344_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__nand2_4
XFILLER_0_132_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07614__A1 _01171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07054_ genblk1\[8\].osc.clkdiv_C.cnt\[15\] _01436_ _01864_ _01868_ _01871_ VGND
+ VGND VPWR VPWR _01872_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11758__B genblk1\[9\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07917__A2 _01858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07956_ genblk1\[7\].osc.clkdiv_C.cnt\[3\] _02656_ _02659_ _02660_ _02662_ VGND VGND
+ VPWR VPWR _02663_ sky130_fd_sc_hd__a221o_1
X_06907_ net28 VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__clkbuf_4
X_07887_ _02469_ _02593_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06587__B _01494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09626_ genblk2\[1\].wave_shpr.div.acc\[15\] _04121_ _04095_ VGND VGND VPWR VPWR
+ _04122_ sky130_fd_sc_hd__mux2_1
X_06838_ _01693_ _01703_ _01704_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_97_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09557_ _04069_ genblk1\[1\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__and2_1
X_06769_ _01644_ _01642_ _01645_ _01600_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_35_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_16
X_08508_ _03210_ _03214_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__xnor2_1
X_09488_ _04033_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07302__B1 _02064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09842__A2 _04247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08439_ _02404_ _02407_ genblk2\[10\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR
+ _03146_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_93_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11450_ genblk2\[8\].wave_shpr.div.fin_quo\[4\] net1321 _00021_ VGND VGND VPWR VPWR
+ _05422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10401_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06408__A2 _01323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11381_ net328 _05356_ _05357_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13120_ clknet_leaf_136_clk _00445_ net43 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10332_ _03717_ _04634_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13051_ clknet_leaf_113_clk net738 net128 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10064__S _04440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10263_ genblk2\[4\].wave_shpr.div.acc\[7\] genblk2\[4\].wave_shpr.div.b1\[7\] VGND
+ VGND VPWR VPWR _04575_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08042__B _01359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12002_ net1204 _02002_ _05802_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__mux2_1
X_10194_ _04404_ _04523_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12904_ clknet_leaf_37_clk _00235_ net104 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ clknet_leaf_64_clk net689 net196 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_26_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ clknet_leaf_91_clk _00099_ net146 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11717_ genblk2\[9\].wave_shpr.div.acc\[21\] genblk2\[9\].wave_shpr.div.acc\[20\]
+ genblk2\[9\].wave_shpr.div.acc\[19\] _05608_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__or4_1
X_12697_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[10\] net172 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_127_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11648_ _05444_ _05441_ genblk2\[8\].wave_shpr.div.i\[0\] VGND VGND VPWR VPWR _05545_
+ sky130_fd_sc_hd__mux2_1
Xinput12 pb[6] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11579_ _05388_ _05368_ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold807 genblk2\[2\].wave_shpr.div.b1\[16\] VGND VGND VPWR VPWR net1025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09329__A _03838_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold818 genblk2\[2\].wave_shpr.div.acc\[15\] VGND VGND VPWR VPWR net1036 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ clknet_leaf_25_clk net624 net86 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold829 genblk2\[2\].wave_shpr.div.b1\[2\] VGND VGND VPWR VPWR net1047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13249_ clknet_leaf_2_clk _00572_ net52 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07810_ net1 net150 _02312_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__and3_1
XANTENNA__07791__B _01263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08790_ _03489_ _03496_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__xor2_1
XANTENNA__06688__A _01577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07780__B1 _01215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07741_ genblk1\[1\].osc.clkdiv_C.cnt\[11\] _01337_ _01312_ genblk1\[1\].osc.clkdiv_C.cnt\[10\]
+ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__o22a_1
XANTENNA__10667__B1 _04855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07672_ _01308_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10131__A2 _04451_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09411_ _03969_ _03973_ _03974_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__a21o_1
X_06623_ genblk1\[3\].osc.clkdiv_C.cnt\[1\] genblk1\[3\].osc.clkdiv_C.cnt\[0\] genblk1\[3\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06886__A2 _01738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_17_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_16
X_09342_ _03797_ _03746_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__or2b_1
X_06554_ net1159 _01466_ _01469_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[10\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09285__B1 _03840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09273_ genblk2\[0\].wave_shpr.div.acc\[1\] _03803_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__or2_1
X_06485_ _01241_ _01337_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__or2_2
XFILLER_0_117_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08224_ _02527_ _02928_ _02929_ _02930_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__a31o_1
XANTENNA__13264__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08155_ genblk1\[3\].osc.clkdiv_C.cnt\[7\] _01483_ _01494_ genblk1\[3\].osc.clkdiv_C.cnt\[6\]
+ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__o22a_1
X_07106_ _01886_ _01910_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08086_ genblk2\[5\].wave_shpr.div.fin_quo\[4\] _02792_ VGND VGND VPWR VPWR _02793_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07037_ _01230_ _01564_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__nand2_4
X_08988_ _03670_ _03671_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__xnor2_1
X_07939_ _02217_ _02553_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__nor2_1
XANTENNA__10658__B1 _04857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10950_ net477 _05057_ _05055_ net515 _05058_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__a221o_1
X_09609_ genblk2\[1\].wave_shpr.div.acc\[12\] _04076_ _04080_ _04108_ VGND VGND VPWR
+ VPWR _00245_ sky130_fd_sc_hd__a22o_1
X_10881_ _05024_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12620_ clknet_leaf_17_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[5\] net83 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__09276__B1 _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12551_ clknet_leaf_60_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[8\] net187 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__10059__S _04238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11502_ net751 _05442_ _05446_ net795 VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12482_ clknet_leaf_108_clk _00044_ net151 VGND VGND VPWR VPWR sig_norm.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11433_ _05358_ _05407_ _05408_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11364_ _05345_ _05342_ _05346_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11398__B genblk2\[8\].wave_shpr.div.b1\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07054__A2 _01436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10315_ _04625_ VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__clkbuf_1
X_13103_ clknet_leaf_12_clk _00428_ net51 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06262__B1 _01223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11295_ _05195_ _05174_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__or2b_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09583__S _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13034_ clknet_leaf_127_clk _00361_ net66 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10246_ _04560_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10177_ genblk2\[3\].wave_shpr.div.acc\[9\] _04510_ _04507_ VGND VGND VPWR VPWR _04511_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06301__A _01238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09503__A1 _03714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12818_ clknet_leaf_67_clk _00151_ net193 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_57_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09806__A2 _04248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ clknet_leaf_46_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[8\] net119 VGND VGND
+ VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_151_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09758__S _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06270_ freq_div.state\[0\] freq_div.state\[1\] VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold604 genblk2\[7\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 genblk2\[8\].wave_shpr.div.acc\[13\] VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 genblk2\[10\].wave_shpr.div.acc\[11\] VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold637 genblk2\[5\].wave_shpr.div.i\[4\] VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 genblk2\[0\].wave_shpr.div.acc\[6\] VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ _00008_ _04356_ net1123 VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__a21oi_1
Xhold659 genblk2\[7\].wave_shpr.div.acc\[4\] VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_122_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08911_ _03611_ _03612_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__nand2_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09891_ net952 _04282_ _04289_ _04308_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__a22o_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08842_ _03545_ _03548_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__and2b_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _03474_ _03479_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout184_A net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07724_ genblk1\[1\].osc.clkdiv_C.cnt\[2\] _01323_ _01313_ genblk1\[1\].osc.clkdiv_C.cnt\[3\]
+ VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__o22a_1
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07505__B1 _02225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09522__A _03853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07655_ _02361_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10668__A _04672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06606_ _01234_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07586_ _02278_ _02279_ _02281_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__a21o_1
X_09325_ _03789_ _03750_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__or2b_1
X_06537_ _01452_ _01458_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09256_ genblk2\[0\].wave_shpr.div.quo\[20\] _03845_ _03847_ net298 _03857_ VGND
+ VGND VPWR VPWR _00143_ sky130_fd_sc_hd__a221o_1
X_06468_ _01373_ _01399_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__nor2_1
XANTENNA__06881__A _01189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08207_ _02310_ _02913_ _02314_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__o21a_1
XFILLER_0_106_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09187_ net1173 VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__inv_2
X_06399_ _01173_ _01175_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__or2_1
XANTENNA__11368__A1 _05245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08138_ genblk2\[4\].wave_shpr.div.fin_quo\[7\] _02309_ _02844_ _02527_ VGND VGND
+ VPWR VPWR _02845_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08069_ genblk1\[5\].osc.clkdiv_C.cnt\[2\] _01592_ _02775_ VGND VGND VPWR VPWR _02776_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10100_ net631 _04457_ _04454_ net538 _04459_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout97_A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11080_ net659 _05057_ _05126_ _05148_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__a22o_1
X_10031_ genblk2\[3\].wave_shpr.div.fin_quo\[2\] net326 _04422_ VGND VGND VPWR VPWR
+ _04425_ sky130_fd_sc_hd__mux2_1
XANTENNA__10342__S _04637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07744__B1 _01344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12096__A2 _05844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11982_ _01441_ _01320_ _03702_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__o21ai_4
X_13721_ clknet_leaf_40_clk _01032_ net118 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10933_ _02188_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13652_ clknet_leaf_40_clk _00965_ net116 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10864_ genblk2\[6\].wave_shpr.div.b1\[13\] genblk2\[6\].wave_shpr.div.acc\[13\]
+ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12603_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[6\] net97 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10795_ genblk2\[5\].wave_shpr.div.acc\[22\] _04817_ _04947_ VGND VGND VPWR VPWR
+ _04948_ sky130_fd_sc_hd__a21o_1
X_13583_ clknet_leaf_76_clk _00898_ net207 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12534_ clknet_leaf_45_clk _00086_ net186 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12465_ clknet_leaf_31_clk smpl_rt_clkdiv.clkDiv_inst.next_hzX net99 VGND VGND VPWR
+ VPWR genblk2\[0\].wave_shpr.div.start sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11202__A _03702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08224__A1 _02527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11416_ genblk2\[8\].wave_shpr.div.b1\[9\] genblk2\[8\].wave_shpr.div.acc\[9\] VGND
+ VGND VPWR VPWR _05392_ sky130_fd_sc_hd__and2b_1
X_12396_ _05965_ _05930_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__or2b_1
XFILLER_0_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11347_ genblk2\[7\].wave_shpr.div.acc\[19\] _05217_ _05334_ VGND VGND VPWR VPWR
+ _05335_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_120_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11278_ net992 _05279_ _05250_ _05282_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__a22o_1
X_10229_ genblk2\[3\].wave_shpr.div.acc\[23\] _04417_ VGND VGND VPWR VPWR _04549_
+ sky130_fd_sc_hd__nor2_1
X_13017_ clknet_leaf_124_clk _00344_ net76 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold1 PWM.pwm_out VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__A _01192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10098__B2 genblk2\[3\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07440_ _02177_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07371_ _02091_ _02124_ _02125_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__and3_1
X_09110_ genblk2\[0\].wave_shpr.div.acc\[5\] genblk2\[0\].wave_shpr.div.b1\[5\] VGND
+ VGND VPWR VPWR _03758_ sky130_fd_sc_hd__or2b_1
X_06322_ genblk1\[0\].osc.clkdiv_C.cnt\[5\] genblk1\[0\].osc.clkdiv_C.cnt\[4\] _01276_
+ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09041_ net1243 _03706_ _03708_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__mux2_1
X_06253_ _01213_ _01214_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__nand2_2
XFILLER_0_115_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06184_ _01094_ _01095_ _01096_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__or3_4
Xhold401 genblk2\[11\].wave_shpr.div.acc\[23\] VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 genblk2\[5\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 genblk2\[11\].wave_shpr.div.acc\[19\] VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold434 genblk2\[0\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12491__RESET_B net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold445 sig_norm.acc\[10\] VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10951__A _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold456 genblk2\[10\].wave_shpr.div.b1\[15\] VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 _00209_ VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 genblk2\[2\].wave_shpr.div.quo\[4\] VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09943_ genblk2\[2\].wave_shpr.div.acc\[23\] _04211_ _04346_ VGND VGND VPWR VPWR
+ _04347_ sky130_fd_sc_hd__a21o_1
Xhold489 genblk2\[2\].wave_shpr.div.acc\[23\] VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ net887 _04282_ _04289_ _04295_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__a22o_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 genblk2\[6\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net1319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1112 genblk2\[5\].wave_shpr.div.quo\[4\] VGND VGND VPWR VPWR net1330 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _02581_ _02580_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__or2b_1
Xhold1123 genblk2\[11\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net1341 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ _03234_ _03462_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__nor2_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06876__A _01336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09252__A _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07707_ _02316_ _02411_ _02413_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__or3_1
XANTENNA__11286__B1 _05283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08687_ _03381_ _03382_ _03298_ _03333_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__o211a_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08151__B1 _01514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ _01229_ _02081_ _02085_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07569_ genblk1\[9\].osc.clkdiv_C.cnt\[15\] _01577_ _02274_ _02275_ VGND VGND VPWR
+ VPWR _02276_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09308_ _03781_ _03754_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__or2b_1
X_10580_ genblk2\[5\].wave_shpr.div.b1\[14\] genblk2\[5\].wave_shpr.div.acc\[14\]
+ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09239_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12250_ _05985_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08206__B2 _02362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11201_ _05241_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__clkbuf_1
X_12181_ _05816_ _05919_ _05921_ _05818_ net748 VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__a32o_1
XANTENNA__07965__B1 _01675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11132_ _05176_ _05190_ _05191_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__a21o_1
Xhold990 genblk2\[9\].wave_shpr.div.b1\[5\] VGND VGND VPWR VPWR net1208 sky130_fd_sc_hd__dlygate4sd3_1
X_11063_ genblk2\[6\].wave_shpr.div.acc\[17\] _05136_ _05022_ VGND VGND VPWR VPWR
+ _05137_ sky130_fd_sc_hd__mux2_1
XANTENNA__08050__B _01355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10014_ _04363_ _04408_ _04409_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08390__B1 _02011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06786__A _01489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11965_ _05786_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__clkbuf_8
X_13704_ clknet_leaf_37_clk _01015_ net113 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10916_ net1286 _01797_ _05042_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__mux2_1
XANTENNA__10101__A _04269_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11896_ _05722_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13635_ clknet_leaf_69_clk _00948_ net212 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10847_ _04979_ _04989_ _04990_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13566_ clknet_leaf_56_clk net305 net182 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10778_ _04813_ _04935_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07410__A _02154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12517_ clknet_leaf_105_clk PWM.next_counter\[1\] net155 VGND VGND VPWR VPWR PWM.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13497_ clknet_leaf_86_clk net618 net178 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12448_ clknet_leaf_105_clk _00027_ net153 VGND VGND VPWR VPWR sig_norm.i\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12379_ net876 _06039_ _06040_ _06056_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06940_ net28 _01781_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__nor2_1
XANTENNA__07971__A3 _01362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06871_ net493 _01724_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__08381__B1 _02336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08610_ _03314_ _03315_ _02789_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__or3_1
X_09590_ _03983_ _04093_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07222__A2_N _02001_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08541_ genblk2\[8\].wave_shpr.div.fin_quo\[0\] _02526_ _02308_ genblk2\[8\].wave_shpr.div.fin_quo\[1\]
+ _02636_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08472_ genblk2\[5\].wave_shpr.div.fin_quo\[3\] _03178_ _02526_ VGND VGND VPWR VPWR
+ _03179_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07423_ _02164_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout147_A net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07354_ genblk1\[11\].osc.clkdiv_C.cnt\[6\] _02108_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10243__A1 _04454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06305_ genblk1\[0\].osc.clkdiv_C.cnt\[3\] _01227_ _01236_ _01266_ VGND VGND VPWR
+ VPWR _01267_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07285_ net1119 _02052_ _02054_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09024_ _02203_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06236_ _01174_ genblk1\[0\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11777__A _04676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold220 genblk2\[11\].wave_shpr.div.quo\[22\] VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__dlygate4sd3_1
X_06167_ _01129_ _01138_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__or2_1
Xhold231 genblk2\[2\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 genblk2\[1\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 genblk2\[5\].wave_shpr.div.quo\[22\] VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 genblk2\[8\].wave_shpr.div.quo\[12\] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold275 genblk1\[5\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 genblk2\[11\].wave_shpr.div.quo\[21\] VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 genblk2\[6\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__dlygate4sd3_1
X_09926_ genblk2\[2\].wave_shpr.div.acc\[25\] genblk2\[2\].wave_shpr.div.acc\[24\]
+ genblk2\[2\].wave_shpr.div.acc\[26\] _04212_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__nor4_1
XANTENNA__12299__A2 _06009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _04247_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__clkbuf_4
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _03217_ _03510_ _03442_ _03443_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__o211a_1
X_09788_ _04244_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12401__A _03941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11259__B1 _05249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _03443_ _03444_ _03428_ _03420_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__a211oi_2
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08124__B1 _01304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ genblk2\[9\].wave_shpr.div.quo\[5\] _05623_ _05624_ net586 VGND VGND VPWR
+ VPWR _00870_ sky130_fd_sc_hd__a22o_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10701_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__and2_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ genblk2\[9\].wave_shpr.div.acc\[0\] VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13420_ clknet_leaf_91_clk _00739_ net147 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10632_ genblk2\[6\].wave_shpr.div.b1\[9\] _01923_ _04834_ VGND VGND VPWR VPWR _04843_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10563_ _04775_ _04789_ _04790_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__a21o_1
X_13351_ clknet_leaf_5_clk _00672_ net47 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11982__A1 _01441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12302_ genblk2\[11\].wave_shpr.div.quo\[3\] _06009_ _06010_ net402 VGND VGND VPWR
+ VPWR _01036_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10494_ _04615_ _04735_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__xnor2_1
X_13282_ clknet_leaf_117_clk _00603_ net137 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_122_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12233_ genblk2\[11\].wave_shpr.div.b1\[15\] genblk2\[11\].wave_shpr.div.acc\[15\]
+ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12164_ genblk2\[10\].wave_shpr.div.acc\[22\] _05908_ genblk2\[10\].wave_shpr.div.acc\[23\]
+ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__or3b_1
X_11115_ genblk2\[7\].wave_shpr.div.acc\[6\] genblk2\[7\].wave_shpr.div.b1\[6\] VGND
+ VGND VPWR VPWR _05175_ sky130_fd_sc_hd__or2b_1
XANTENNA__13548__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12095_ genblk2\[10\].wave_shpr.div.acc\[5\] _05858_ _05787_ VGND VGND VPWR VPWR
+ _05859_ sky130_fd_sc_hd__mux2_1
X_11046_ _05007_ _05123_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11498__B1 _05446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07405__A _02147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12997_ clknet_leaf_132_clk _00326_ net60 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07124__B _01355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11948_ genblk2\[10\].wave_shpr.div.b1\[12\] genblk2\[10\].wave_shpr.div.acc\[12\]
+ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__and2b_1
X_11879_ net556 _05684_ _05685_ _05711_ VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13618_ clknet_leaf_84_clk _00931_ net204 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08236__A net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13549_ clknet_leaf_110_clk _00864_ net152 VGND VGND VPWR VPWR sig_norm.b1\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07070_ net1092 _01887_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09067__A _02155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06601__B1 _01508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07972_ _02672_ _02673_ _02678_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__o21ai_2
X_09711_ genblk2\[2\].wave_shpr.div.b1\[9\] genblk2\[2\].wave_shpr.div.acc\[9\] VGND
+ VGND VPWR VPWR _04191_ sky130_fd_sc_hd__and2b_1
X_06923_ genblk1\[6\].osc.clkdiv_C.cnt\[6\] _01768_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__nor2_1
XANTENNA__06227__B1_N _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09642_ genblk2\[1\].wave_shpr.div.acc\[19\] _04130_ VGND VGND VPWR VPWR _04134_
+ sky130_fd_sc_hd__nand2_1
X_06854_ _01693_ _01713_ _01714_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__10700__A2 _02183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06785_ genblk1\[5\].osc.clkdiv_C.cnt\[4\] _01483_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__xnor2_1
X_09573_ _03976_ _03968_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__or2b_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _02216_ _02552_ genblk2\[9\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR
+ _03231_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07034__B _01359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09530__A _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08455_ _03159_ _03160_ _03161_ _02694_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__a211o_1
XANTENNA__10676__A _04672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07406_ _02151_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__inv_2
X_08386_ _01200_ genblk1\[2\].osc.clkdiv_C.cnt\[4\] genblk1\[2\].osc.clkdiv_C.cnt\[5\]
+ _01441_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07337_ genblk1\[11\].osc.clkdiv_C.cnt\[1\] genblk1\[11\].osc.clkdiv_C.cnt\[0\] genblk1\[11\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07268_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _02041_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07632__A2 _01262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09007_ _03683_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__clkbuf_1
X_06219_ _01174_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__buf_6
XFILLER_0_104_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10615__S _04637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07199_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01981_ _01984_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08593__B1 _02361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07209__B _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09909_ _04250_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__clkbuf_4
X_12920_ clknet_leaf_35_clk _00251_ net118 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ clknet_leaf_118_clk _00182_ net138 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06371__A2 _01311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11802_ _03693_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__clkbuf_4
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ clknet_leaf_40_clk _00115_ net117 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11733_ _05619_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__clkbuf_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11652__B1 _05448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11664_ genblk2\[9\].wave_shpr.div.acc\[15\] genblk2\[9\].wave_shpr.div.b1\[15\]
+ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__or2b_1
XFILLER_0_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13403_ clknet_leaf_92_clk _00722_ net147 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10615_ genblk2\[6\].wave_shpr.div.b1\[2\] _01684_ _04637_ VGND VGND VPWR VPWR _04833_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11595_ _05441_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__clkbuf_4
X_13334_ clknet_leaf_6_clk _00655_ net48 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10546_ genblk2\[5\].wave_shpr.div.acc\[6\] genblk2\[5\].wave_shpr.div.b1\[6\] VGND
+ VGND VPWR VPWR _04774_ sky130_fd_sc_hd__or2b_1
XFILLER_0_51_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13265_ clknet_leaf_0_clk _00588_ net38 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10477_ _04608_ _04569_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__or2b_1
XFILLER_0_20_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12216_ _05936_ _05952_ _05953_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13196_ clknet_leaf_114_clk _00519_ net134 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_103_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12147_ net590 _05876_ _05883_ _05898_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__a22o_1
XANTENNA__07119__B _01227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09615__A _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07139__A1 genblk1\[9\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12078_ genblk2\[10\].wave_shpr.div.acc\[1\] _05845_ _05787_ VGND VGND VPWR VPWR
+ _05846_ sky130_fd_sc_hd__mux2_1
X_11029_ _04999_ _05110_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07899__A1_N _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06570_ genblk1\[2\].osc.clkdiv_C.cnt\[16\] _01478_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07789__B _01263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09851__A3 _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08240_ _02682_ _02689_ _02683_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08171_ _02861_ _02862_ _02865_ _02876_ _02877_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_133_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07122_ genblk1\[9\].osc.clkdiv_C.cnt\[6\] _01334_ _01328_ genblk1\[9\].osc.clkdiv_C.cnt\[13\]
+ _01921_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__o221a_1
XANTENNA__07614__A2 _01192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07053_ genblk1\[8\].osc.clkdiv_C.cnt\[12\] _01869_ _01870_ genblk1\[8\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_3_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10382__B1 _04655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07955_ _02661_ _02653_ _02652_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__or3b_1
X_06906_ _01675_ _01727_ _01737_ _01756_ _01759_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__10134__B1 _04455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07886_ genblk2\[1\].wave_shpr.div.fin_quo\[7\] _02539_ _02591_ _02592_ VGND VGND
+ VPWR VPWR _02593_ sky130_fd_sc_hd__a22o_1
X_09625_ _03999_ _04120_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06837_ genblk1\[5\].osc.clkdiv_C.cnt\[4\] _01700_ genblk1\[5\].osc.clkdiv_C.cnt\[5\]
+ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09556_ _03707_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__clkbuf_4
X_06768_ genblk1\[4\].osc.clkdiv_C.cnt\[13\] _01641_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__or2_1
XANTENNA__06884__A _01241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08507_ _03114_ _03213_ _03122_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09487_ net1304 _04032_ _04024_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__mux2_1
X_06699_ _01320_ _01321_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__nand2_4
X_08438_ _03141_ _03144_ _02901_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09055__A1 _03704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08369_ _03052_ _03053_ _03030_ _03051_ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_150_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10400_ net531 _04661_ _04663_ genblk2\[4\].wave_shpr.div.quo\[16\] _04668_ VGND
+ VGND VPWR VPWR _00476_ sky130_fd_sc_hd__a221o_1
XANTENNA__07066__B1 _01870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11380_ net328 _05356_ _03855_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08604__A _02261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07053__A2_N _01869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10331_ _04633_ _01304_ _03689_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10345__S _04637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10262_ genblk2\[4\].wave_shpr.div.acc\[8\] genblk2\[4\].wave_shpr.div.b1\[8\] VGND
+ VGND VPWR VPWR _04574_ sky130_fd_sc_hd__or2b_1
X_13050_ clknet_leaf_113_clk net327 net128 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12001_ _05805_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__clkbuf_1
X_10193_ _04405_ _04365_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__or2b_1
XANTENNA__11190__B1_N _04241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12903_ clknet_leaf_37_clk net753 net104 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12834_ clknet_leaf_64_clk _00167_ net196 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06794__A _01440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ clknet_leaf_93_clk _00098_ net146 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ genblk2\[9\].wave_shpr.div.acc\[18\] _05607_ VGND VGND VPWR VPWR _05608_
+ sky130_fd_sc_hd__or2_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12696_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[9\] net172 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_154_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11647_ net615 _05448_ _05445_ _05544_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__a22o_1
Xinput13 pb[7] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11578_ net950 _05447_ _05484_ _05494_ VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06960__C _01514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13317_ clknet_leaf_24_clk net345 net88 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold808 genblk2\[9\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold819 genblk2\[5\].wave_shpr.div.acc\[7\] VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ _04655_ _04757_ _04759_ _04657_ net734 VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__a32o_1
XANTENNA__08233__B _02885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13248_ clknet_leaf_13_clk net911 net52 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08557__B1 genblk2\[8\].wave_shpr.div.fin_quo\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13179_ clknet_leaf_131_clk _00504_ net65 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08021__A2 _01577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06969__A _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07740_ genblk1\[1\].osc.clkdiv_C.cnt\[9\] _01334_ _01356_ genblk1\[1\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_74_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09521__A2 _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07671_ _01308_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__and2_1
X_09410_ genblk2\[1\].wave_shpr.div.b1\[2\] genblk2\[1\].wave_shpr.div.acc\[2\] VGND
+ VGND VPWR VPWR _03974_ sky130_fd_sc_hd__and2b_1
X_06622_ genblk1\[3\].osc.clkdiv_C.cnt\[2\] genblk1\[3\].osc.clkdiv_C.cnt\[1\] genblk1\[3\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__and3_1
X_09341_ net786 _03903_ _03910_ _03919_ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__a22o_1
X_06553_ _01451_ _01468_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_89_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06484_ genblk1\[2\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09272_ _03865_ _03866_ net1066 _03836_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_23_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_132_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08223_ genblk2\[5\].wave_shpr.div.fin_quo\[6\] _02308_ _02791_ VGND VGND VPWR VPWR
+ _02930_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09037__A1 _03704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10954__A _04676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07048__B1 _01336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12041__B1 _05816_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08154_ _02858_ _02859_ _02860_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07105_ genblk1\[8\].osc.clkdiv_C.cnt\[13\] genblk1\[8\].osc.clkdiv_C.cnt\[12\] _01906_
+ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08085_ genblk2\[5\].wave_shpr.div.fin_quo\[0\] genblk2\[5\].wave_shpr.div.fin_quo\[1\]
+ genblk2\[5\].wave_shpr.div.fin_quo\[2\] genblk2\[5\].wave_shpr.div.fin_quo\[3\]
+ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__or4_1
XANTENNA__09239__B genblk1\[0\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07036_ genblk1\[8\].osc.clkdiv_C.cnt\[16\] _01853_ _01578_ VGND VGND VPWR VPWR _01854_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09255__A _03853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08987_ _03134_ _03135_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__nor2_1
XANTENNA__06598__B _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
X_07938_ genblk2\[8\].wave_shpr.div.fin_quo\[7\] _02539_ _02636_ _02644_ VGND VGND
+ VPWR VPWR _02645_ sky130_fd_sc_hd__a211o_1
XANTENNA__09512__A2 _04043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07869_ genblk2\[0\].wave_shpr.div.fin_quo\[0\] _02524_ _02307_ genblk2\[0\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__a22o_1
XANTENNA__11724__S _00023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09608_ net366 _04107_ _04095_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__mux2_1
X_10880_ genblk2\[6\].wave_shpr.div.fin_quo\[0\] _05023_ _00017_ VGND VGND VPWR VPWR
+ _05024_ sky130_fd_sc_hd__mux2_1
XANTENNA__07503__A _02223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09539_ net462 _04052_ _04053_ genblk2\[1\].wave_shpr.div.quo\[15\] _04060_ VGND
+ VGND VPWR VPWR _00223_ sky130_fd_sc_hd__a221o_1
XANTENNA__08079__A2 _01355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09276__A1 _03839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12550_ clknet_leaf_60_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[7\] net186 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11501_ genblk2\[8\].wave_shpr.div.quo\[4\] _05442_ _05446_ net346 VGND VGND VPWR
+ VPWR _00799_ sky130_fd_sc_hd__a22o_1
X_12481_ clknet_leaf_108_clk net1028 net151 VGND VGND VPWR VPWR sig_norm.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11432_ genblk2\[8\].wave_shpr.div.b1\[17\] genblk2\[8\].wave_shpr.div.acc\[17\]
+ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10075__S _04440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11363_ genblk2\[7\].wave_shpr.div.acc\[24\] _05273_ _05342_ VGND VGND VPWR VPWR
+ _05346_ sky130_fd_sc_hd__or3b_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09864__S _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13102_ clknet_leaf_118_clk _00013_ net139 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
X_10314_ genblk2\[4\].wave_shpr.div.fin_quo\[1\] net1309 _00013_ VGND VGND VPWR VPWR
+ _04625_ sky130_fd_sc_hd__mux2_1
X_11294_ net893 _05279_ _05283_ _05294_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ clknet_leaf_123_clk _00360_ net79 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10245_ genblk2\[3\].wave_shpr.div.i\[1\] genblk2\[3\].wave_shpr.div.i\[0\] genblk2\[3\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__and3_1
XANTENNA__08003__A2 _01666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10176_ _04396_ _04509_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07762__A1 _02458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10104__A _04455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout190 net198 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06301__B _01262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12817_ clknet_leaf_59_clk _00150_ net193 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ clknet_leaf_50_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[7\] net111 VGND VGND
+ VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12679_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[10\] net82 VGND VGND
+ VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12023__B1 _05817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold605 genblk2\[0\].wave_shpr.div.acc\[5\] VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold616 genblk2\[5\].wave_shpr.div.b1\[16\] VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 genblk2\[2\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 _04964_ VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold649 genblk2\[6\].wave_shpr.div.acc\[8\] VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__dlygate4sd3_1
X_08910_ _03586_ net26 sig_norm.acc\[4\] VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11809__S _05613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ genblk2\[2\].wave_shpr.div.acc\[9\] _04307_ _04301_ VGND VGND VPWR VPWR _04308_
+ sky130_fd_sc_hd__mux2_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08841_ _03542_ _03544_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__or2_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _03477_ _03478_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__xnor2_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12626__RESET_B net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07307__B _01223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07723_ genblk1\[1\].osc.clkdiv_C.cnt\[2\] _01323_ _02429_ genblk1\[1\].osc.clkdiv_C.cnt\[1\]
+ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07654_ _02307_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06605_ _01512_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__clkbuf_4
X_07585_ genblk1\[9\].osc.clkdiv_C.cnt\[3\] _01311_ _02290_ _02291_ VGND VGND VPWR
+ VPWR _02292_ sky130_fd_sc_hd__a22o_1
X_09324_ net920 _03903_ _03877_ _03906_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06536_ genblk1\[2\].osc.clkdiv_C.cnt\[4\] _01456_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09255_ _03853_ genblk1\[0\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__and2_1
XANTENNA__10684__A _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06467_ genblk1\[1\].osc.clkdiv_C.cnt\[12\] _01398_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__and2_1
XANTENNA__06881__B _01678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08206_ _02911_ _02912_ genblk2\[9\].wave_shpr.div.fin_quo\[6\] _02362_ VGND VGND
+ VPWR VPWR _02913_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09186_ _03704_ net651 _03820_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__a21o_1
X_06398_ _01188_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08137_ genblk2\[4\].wave_shpr.div.fin_quo\[6\] _02843_ VGND VGND VPWR VPWR _02844_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08068_ _01196_ _01254_ genblk1\[5\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR _02775_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07019_ _01822_ _01842_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__nor2_1
X_10030_ _04424_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07744__A1 genblk1\[1\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11540__A2 _05441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07744__B2 genblk1\[1\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11981_ _05795_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__clkbuf_1
X_13720_ clknet_leaf_39_clk _01031_ net115 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10932_ _05050_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13651_ clknet_leaf_41_clk _00964_ net116 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10863_ _04971_ _05005_ _05006_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12602_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[5\] net95 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13582_ clknet_leaf_76_clk _00897_ net207 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10794_ _04818_ _04819_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__and2b_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12533_ clknet_leaf_61_clk _00085_ net186 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06791__B _01578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12464_ clknet_leaf_103_clk _00037_ net156 VGND VGND VPWR VPWR PWM.final_sample_in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11415_ _05367_ _05389_ _05390_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__a21o_1
X_12395_ net875 _06039_ _06040_ _06068_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11346_ genblk2\[7\].wave_shpr.div.acc\[19\] _05331_ VGND VGND VPWR VPWR _05334_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_120_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11277_ genblk2\[7\].wave_shpr.div.acc\[2\] _05281_ _05222_ VGND VGND VPWR VPWR _05282_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12314__A _03942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09185__B1 _03819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13016_ clknet_leaf_121_clk _00011_ net77 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07408__A _02152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10228_ net1000 _04457_ _04522_ _04548_ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10159_ _04496_ _04388_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__xnor2_1
Xhold2 genblk2\[10\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10098__A2 _04457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07143__A genblk1\[9\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07370_ genblk1\[11\].osc.clkdiv_C.cnt\[9\] _02119_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__or2_1
X_06321_ net1133 _01276_ _01278_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06252_ _01187_ _01188_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__nand2b_4
X_09040_ _03707_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__buf_8
XFILLER_0_60_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06183_ _01099_ _01150_ _01154_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold402 genblk2\[6\].wave_shpr.div.quo\[13\] VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold413 genblk2\[3\].wave_shpr.div.quo\[10\] VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold424 PWM.counter\[1\] VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 genblk2\[0\].wave_shpr.div.acc\[23\] VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold446 genblk2\[1\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 genblk2\[4\].wave_shpr.div.quo\[12\] VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 genblk2\[9\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ _04212_ _04335_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__nor2_1
Xhold479 _00296_ VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ genblk2\[2\].wave_shpr.div.acc\[5\] _04294_ _04214_ VGND VGND VPWR VPWR _04295_
+ sky130_fd_sc_hd__mux2_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _03482_ _03529_ _03530_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__or3_1
Xhold1102 genblk2\[6\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net1320 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 genblk2\[8\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net1331 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07037__B _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1124 genblk2\[5\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net1342 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ _03232_ _03233_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__nor2_1
XANTENNA__06876__B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10089__A2 _04452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07706_ genblk2\[10\].wave_shpr.div.fin_quo\[4\] genblk2\[10\].wave_shpr.div.fin_quo\[5\]
+ _02404_ _02409_ _02412_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__o41a_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _03386_ _03392_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _02338_ _02340_ _02341_ _02342_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07568_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01349_ _01246_ genblk1\[9\].osc.clkdiv_C.cnt\[13\]
+ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09307_ net956 _03870_ _03877_ _03893_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06519_ genblk1\[2\].osc.clkdiv_C.cnt\[7\] _01433_ _01418_ genblk1\[2\].osc.clkdiv_C.cnt\[4\]
+ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_119_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10618__S _04834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07499_ net18 net17 VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__or2b_1
XFILLER_0_63_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09238_ _03838_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__buf_2
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09169_ genblk2\[0\].wave_shpr.div.fin_quo\[6\] net652 _00001_ VGND VGND VPWR VPWR
+ _03811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11200_ genblk2\[8\].wave_shpr.div.b1\[11\] _01565_ _05237_ VGND VGND VPWR VPWR _05241_
+ sky130_fd_sc_hd__mux2_1
X_12180_ _05920_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11131_ genblk2\[7\].wave_shpr.div.b1\[5\] genblk2\[7\].wave_shpr.div.acc\[5\] VGND
+ VGND VPWR VPWR _05191_ sky130_fd_sc_hd__and2b_1
Xhold980 _04222_ VGND VGND VPWR VPWR net1198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold991 genblk2\[9\].wave_shpr.div.acc\[0\] VGND VGND VPWR VPWR net1209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11062_ _05015_ _05135_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06132__A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11513__A2 _05448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10013_ genblk2\[3\].wave_shpr.div.b1\[15\] genblk2\[3\].wave_shpr.div.acc\[15\]
+ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06786__B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11964_ genblk2\[10\].wave_shpr.div.acc\[25\] genblk2\[10\].wave_shpr.div.acc\[26\]
+ _05785_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__or3_2
XFILLER_0_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13703_ clknet_leaf_96_clk _01014_ net161 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10915_ _03707_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11895_ _03838_ _03835_ genblk2\[0\].wave_shpr.div.i\[0\] VGND VGND VPWR VPWR _05722_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13634_ clknet_leaf_69_clk _00947_ net211 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10846_ genblk2\[6\].wave_shpr.div.b1\[4\] genblk2\[6\].wave_shpr.div.acc\[4\] VGND
+ VGND VPWR VPWR _04990_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13565_ clknet_leaf_57_clk _00880_ net182 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10777_ _04814_ _04763_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11213__A _02170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12516_ clknet_leaf_105_clk PWM.next_counter\[0\] net155 VGND VGND VPWR VPWR PWM.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07653__B1 _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13496_ clknet_leaf_86_clk net264 net178 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12447_ clknet_leaf_106_clk net940 net153 VGND VGND VPWR VPWR sig_norm.i\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12378_ genblk2\[11\].wave_shpr.div.acc\[7\] _06054_ _06055_ VGND VGND VPWR VPWR
+ _06056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11752__A2 _05623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11329_ net809 _05311_ _05315_ _05321_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08905__B1 _02248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06870_ _01725_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[16\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__10712__B1 _04857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08540_ _02647_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__inv_2
X_08471_ _03176_ _03177_ _02789_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07422_ _02147_ _02163_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07353_ _02111_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06304_ genblk1\[0\].osc.clkdiv_C.cnt\[1\] _01235_ _01253_ _01260_ _01265_ VGND VGND
+ VPWR VPWR _01266_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07284_ _02026_ _02053_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09023_ genblk2\[9\].wave_shpr.div.i\[1\] genblk2\[9\].wave_shpr.div.i\[0\] genblk2\[9\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__nand3_1
XFILLER_0_142_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06235_ _01196_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__buf_4
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold210 sig_norm.acc_next\[0\] VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09528__A _03853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06166_ _01128_ _01113_ _01117_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__and3_1
Xhold221 _01056_ VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold232 genblk2\[8\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold243 _00215_ VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10173__S _04507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold254 genblk2\[4\].wave_shpr.div.acc\[21\] VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold265 genblk2\[11\].wave_shpr.div.quo\[19\] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _00569_ VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 genblk2\[8\].wave_shpr.div.quo\[23\] VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09925_ net580 _04315_ _04322_ _04334_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__a22o_1
Xhold298 _00636_ VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ _04251_ _04279_ _04281_ _04253_ net1137 VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__a32o_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _03431_ _03438_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__nand2_1
XANTENNA__09263__A _03853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09787_ genblk2\[3\].wave_shpr.div.b1\[15\] _01365_ _04238_ VGND VGND VPWR VPWR _04244_
+ sky130_fd_sc_hd__mux2_1
X_06999_ genblk1\[7\].osc.clkdiv_C.cnt\[5\] genblk1\[7\].osc.clkdiv_C.cnt\[4\] _01827_
+ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__and3_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _03428_ _03420_ _03443_ _03444_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__o211a_2
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _03371_ _03375_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__xnor2_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11732__S _00023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ net324 _02183_ _04856_ net459 _04877_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__a221o_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ genblk2\[9\].wave_shpr.div.b1\[1\] VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10631_ _04842_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_812 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13350_ clknet_leaf_5_clk _00671_ net45 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07635__B1 _01235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07230__B _01432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10562_ genblk2\[5\].wave_shpr.div.b1\[5\] genblk2\[5\].wave_shpr.div.acc\[5\] VGND
+ VGND VPWR VPWR _04790_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12301_ net402 _06009_ _06010_ net769 VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13281_ clknet_leaf_122_clk _00602_ net79 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10493_ _04616_ _04565_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__or2b_1
XFILLER_0_32_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09388__B1 _03819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12232_ _05928_ _05968_ _05969_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__a21o_1
X_12163_ net906 _05818_ _05883_ _05909_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__a22o_1
XANTENNA__10942__B1 _05056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11114_ genblk2\[7\].wave_shpr.div.acc\[7\] genblk2\[7\].wave_shpr.div.b1\[7\] VGND
+ VGND VPWR VPWR _05174_ sky130_fd_sc_hd__or2b_1
X_12094_ _05857_ _05755_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__xnor2_1
X_11045_ _05008_ _04970_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09173__A _01342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13517__RESET_B net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12996_ clknet_leaf_132_clk _00325_ net60 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08115__A1 _01172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11947_ _05737_ _05767_ _05768_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13170__RESET_B net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11878_ _05709_ _05710_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__nand2_1
X_13617_ clknet_leaf_94_clk _00930_ net160 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10829_ genblk2\[6\].wave_shpr.div.acc\[10\] genblk2\[6\].wave_shpr.div.b1\[10\]
+ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__or2b_1
XFILLER_0_43_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13548_ clknet_leaf_110_clk _00863_ net152 VGND VGND VPWR VPWR sig_norm.b1\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13479_ clknet_leaf_99_clk net744 net168 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07971_ _01201_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01362_ _02677_ VGND VGND VPWR
+ VPWR _02678_ sky130_fd_sc_hd__o31a_1
X_09710_ _04165_ _04188_ _04189_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__a21o_1
X_06922_ genblk1\[6\].osc.clkdiv_C.cnt\[6\] _01768_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__and2_1
XANTENNA__10721__S _04821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09551__B1 _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09083__A _02170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09641_ genblk2\[1\].wave_shpr.div.acc\[19\] _04130_ VGND VGND VPWR VPWR _04133_
+ sky130_fd_sc_hd__or2_1
X_06853_ genblk1\[5\].osc.clkdiv_C.cnt\[11\] genblk1\[5\].osc.clkdiv_C.cnt\[10\] _01710_
+ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__and3_1
X_09572_ _04046_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__clkbuf_4
X_06784_ _01436_ _01304_ genblk1\[5\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _01656_
+ sky130_fd_sc_hd__a21oi_1
X_08523_ _03227_ _03229_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__and2b_1
XANTENNA__09811__A _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08454_ _02216_ _02553_ genblk2\[7\].wave_shpr.div.fin_quo\[4\] VGND VGND VPWR VPWR
+ _03161_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07405_ _02147_ _02150_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10168__S _04420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08385_ genblk1\[2\].osc.clkdiv_C.cnt\[4\] _01439_ _01418_ genblk1\[2\].osc.clkdiv_C.cnt\[3\]
+ _03091_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07617__B1 _02064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07336_ _02097_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12893__RESET_B net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07267_ _02027_ _02041_ _02042_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_103_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09006_ net1168 net1170 _01154_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__mux2_1
X_06218_ _01174_ _01177_ _01179_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__a21o_2
XFILLER_0_104_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07198_ _01952_ _01983_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06149_ _01119_ _01120_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09790__B1 _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09908_ net1002 _04315_ _04289_ _04321_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout72_A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09839_ _04269_ genblk1\[2\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__and2_1
X_12850_ clknet_leaf_118_clk _00181_ net138 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _02203_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ clknet_leaf_40_clk _00114_ net115 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11732_ genblk2\[9\].wave_shpr.div.fin_quo\[5\] net1317 _00023_ VGND VGND VPWR VPWR
+ _05619_ sky130_fd_sc_hd__mux2_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11652__A1 _05449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07320__A2 _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _05439_ genblk2\[9\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR _05555_
+ sky130_fd_sc_hd__nor2_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13402_ clknet_leaf_90_clk net303 net147 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10614_ _04832_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11594_ net917 _05447_ _05484_ _05506_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__a22o_1
X_13333_ clknet_leaf_9_clk _00654_ net54 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10545_ genblk2\[5\].wave_shpr.div.acc\[7\] genblk2\[5\].wave_shpr.div.b1\[7\] VGND
+ VGND VPWR VPWR _04773_ sky130_fd_sc_hd__or2b_1
XFILLER_0_52_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_130_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_130_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_107_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13264_ clknet_leaf_1_clk _00587_ net38 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10476_ _04654_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12215_ genblk2\[11\].wave_shpr.div.b1\[6\] genblk2\[11\].wave_shpr.div.acc\[6\]
+ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13195_ clknet_leaf_128_clk _00518_ net132 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10107__A _04269_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12146_ genblk2\[10\].wave_shpr.div.acc\[17\] _05897_ _05786_ VGND VGND VPWR VPWR
+ _05898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13769__RESET_B net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07236__A2_N _02001_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12077_ _05746_ _05747_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__xor2_1
XANTENNA__07139__A2 _01246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11028_ _05000_ _04974_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10694__A2 _02183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12979_ clknet_leaf_124_clk _00308_ net72 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06974__B _01675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08170_ genblk1\[3\].osc.clkdiv_C.cnt\[10\] _01508_ _01507_ genblk1\[3\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__a22o_1
X_07121_ genblk1\[9\].osc.clkdiv_C.cnt\[2\] _01920_ _01855_ genblk1\[9\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__o22a_1
XFILLER_0_132_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10716__S _04821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_121_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_121_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__07614__A3 _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07052_ _01441_ _01226_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__nor2_4
XANTENNA__09078__A _03702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07954_ genblk1\[7\].osc.clkdiv_C.cnt\[4\] _01805_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__and2_1
X_06905_ genblk1\[6\].osc.clkdiv_C.cnt\[3\] _01758_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__xor2_1
X_07885_ _02526_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09624_ _04000_ _03956_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__or2b_1
X_06836_ genblk1\[5\].osc.clkdiv_C.cnt\[5\] genblk1\[5\].osc.clkdiv_C.cnt\[4\] _01700_
+ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__and3_1
XANTENNA__07045__B _01430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_cap29 _01372_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlymetal6s2s_1
X_09555_ net632 _04042_ _04046_ genblk2\[1\].wave_shpr.div.quo\[23\] _04068_ VGND
+ VGND VPWR VPWR _00231_ sky130_fd_sc_hd__a221o_1
X_06767_ genblk1\[4\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__inv_2
XANTENNA__11282__S _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08506_ _03211_ _03212_ genblk2\[2\].wave_shpr.div.fin_quo\[6\] _02468_ VGND VGND
+ VPWR VPWR _03213_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09486_ _01431_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__inv_2
X_06698_ genblk1\[4\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07302__A2 _01256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08437_ _02525_ _03142_ _03143_ _02361_ genblk2\[11\].wave_shpr.div.fin_quo\[3\]
+ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08368_ _03071_ _03074_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07066__A1 genblk1\[8\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07319_ _02080_ _01242_ _01423_ _02081_ _02082_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10626__S _04834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07066__B2 genblk1\[8\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_112_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_112_clk sky130_fd_sc_hd__clkbuf_16
X_08299_ _02897_ _02925_ _02926_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10330_ genblk2\[5\].wave_shpr.div.b1\[1\] VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06405__A _01172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10261_ genblk2\[4\].wave_shpr.div.acc\[9\] genblk2\[4\].wave_shpr.div.b1\[9\] VGND
+ VGND VPWR VPWR _04573_ sky130_fd_sc_hd__or2b_1
XANTENNA_hold586_A genblk2\[0\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12000_ net1217 _03706_ _05802_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__mux2_1
X_10192_ _04455_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__06585__A1_N _01490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09515__B1 _04047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11484__A2_N _01490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12902_ clknet_leaf_30_clk _00233_ net104 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12833_ clknet_leaf_64_clk _00166_ net196 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06794__B _01171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ clknet_leaf_92_clk _00097_ net148 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11715_ _05554_ _05605_ _05606_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__a21o_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[8\] net172 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_4
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11646_ genblk2\[8\].wave_shpr.div.acc\[25\] _05414_ _05543_ VGND VGND VPWR VPWR
+ _05544_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_37_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput14 pb[8] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07057__A1 genblk1\[8\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08254__B1 _02261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_103_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_103_clk sky130_fd_sc_hd__clkbuf_16
X_11577_ genblk2\[8\].wave_shpr.div.acc\[6\] _05492_ _05493_ VGND VGND VPWR VPWR _05494_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13316_ clknet_leaf_9_clk _00637_ net50 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10528_ _04758_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__inv_2
Xhold809 sig_norm.acc\[5\] VGND VGND VPWR VPWR net1027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13247_ clknet_leaf_2_clk _00570_ net52 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08006__B1 _01738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10459_ _04600_ _04573_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08557__A1 genblk2\[8\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13178_ clknet_leaf_131_clk _00503_ net65 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12129_ _05771_ _05884_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12105__A2 _05844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07146__A _01336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10667__A2 _04858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07670_ _02375_ _02376_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__or2_1
X_06621_ _01527_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09340_ genblk2\[0\].wave_shpr.div.acc\[16\] _03918_ _03889_ VGND VGND VPWR VPWR
+ _03919_ sky130_fd_sc_hd__mux2_1
X_06552_ genblk1\[2\].osc.clkdiv_C.cnt\[10\] genblk1\[2\].osc.clkdiv_C.cnt\[9\] _01464_
+ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09271_ genblk2\[0\].wave_shpr.div.b1\[0\] genblk2\[0\].wave_shpr.div.acc\[0\] _03804_
+ _03863_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__a31o_1
X_06483_ genblk1\[1\].osc.clkdiv_C.cnt\[17\] _01407_ _01409_ _01374_ VGND VGND VPWR
+ VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[17\] sky130_fd_sc_hd__o211a_1
XFILLER_0_117_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08222_ _02789_ _02793_ genblk2\[5\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR
+ _02929_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07048__A1 _01174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08153_ genblk1\[3\].osc.clkdiv_C.cnt\[5\] _01500_ _01494_ genblk1\[3\].osc.clkdiv_C.cnt\[6\]
+ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout122_A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07104_ genblk1\[8\].osc.clkdiv_C.cnt\[12\] _01906_ _01909_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08084_ _02790_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07035_ genblk1\[8\].osc.clkdiv_C.cnt\[10\] _01852_ _01248_ VGND VGND VPWR VPWR _01853_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09536__A _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11785__B genblk1\[9\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10355__A1 _04645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11277__S _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10181__S _04507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08986_ _03225_ _03570_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__nor2_1
XANTENNA__07056__A genblk1\[8\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07937_ _02642_ _02643_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__and2b_1
XANTENNA__10658__A2 _04853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07868_ _02509_ _02572_ _02574_ _02517_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09607_ _03991_ _04106_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__xnor2_1
X_06819_ _01665_ _01668_ _01673_ _01690_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__or4b_1
X_07799_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] _01349_ _01577_ genblk1\[0\].osc.clkdiv_C.cnt\[16\]
+ _02505_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09538_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08484__B1 _02885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09469_ genblk2\[2\].wave_shpr.div.b1\[3\] _01231_ _03822_ VGND VGND VPWR VPWR _04022_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11083__A2 _05057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11500_ net346 _05442_ _05446_ net709 VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12480_ clknet_leaf_108_clk _00042_ net152 VGND VGND VPWR VPWR sig_norm.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11431_ _05359_ _05405_ _05406_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10043__B1 _03733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08787__B2 _02468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11362_ genblk2\[7\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__inv_2
XANTENNA__06135__A net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10594__A1 _04821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13101_ clknet_leaf_122_clk _00012_ net78 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
X_10313_ _04624_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07898__A1_N genblk1\[8\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06262__A2 _01221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11293_ genblk2\[7\].wave_shpr.div.acc\[6\] _05293_ _05222_ VGND VGND VPWR VPWR _05294_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13032_ clknet_leaf_121_clk _00359_ net78 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10244_ genblk2\[3\].wave_shpr.div.i\[1\] genblk2\[3\].wave_shpr.div.i\[0\] genblk2\[3\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10175_ _04397_ _04369_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__or2b_1
XANTENNA__07762__A2 _02459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout180 net185 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__buf_2
XANTENNA__06970__B1 _01801_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout191 net198 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12816_ clknet_leaf_58_clk _00149_ net192 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ clknet_leaf_49_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[6\] net108 VGND VGND
+ VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12678_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[9\] net142 VGND VGND
+ VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_37_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08227__B1 _02316_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11629_ _05471_ _05532_ net690 _05442_ VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold606 _00154_ VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 genblk2\[5\].wave_shpr.div.acc\[15\] VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold628 genblk2\[8\].wave_shpr.div.acc\[14\] VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 genblk2\[2\].wave_shpr.div.acc\[12\] VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _03464_ _03526_ _03528_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__o21ai_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07202__A1 genblk1\[9\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _03304_ _03306_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__xnor2_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07307__C _01678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07722_ _01330_ _01262_ _01591_ _01172_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__o211ai_1
XANTENNA_clkbuf_4_7_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09091__A _01201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07653_ _02349_ _02351_ _02221_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__a21o_1
XANTENNA__12666__RESET_B net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07910__C1 _01238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06604_ _01171_ _01192_ _01208_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07584_ genblk1\[9\].osc.clkdiv_C.cnt\[2\] _01234_ _01310_ genblk1\[9\].osc.clkdiv_C.cnt\[3\]
+ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__o22a_1
XFILLER_0_149_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09323_ genblk2\[0\].wave_shpr.div.acc\[12\] _03905_ _03889_ VGND VGND VPWR VPWR
+ _03906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06535_ _01452_ _01456_ _01457_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09254_ net298 _03845_ _03847_ net466 _03856_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06466_ _01373_ _01397_ _01398_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_29_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08205_ genblk2\[9\].wave_shpr.div.fin_quo\[5\] _02303_ _02265_ _02316_ VGND VGND
+ VPWR VPWR _02912_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09185_ _01430_ _01344_ _03819_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_141_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06397_ genblk1\[1\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08136_ _02842_ genblk2\[4\].wave_shpr.div.fin_quo\[5\] _02837_ VGND VGND VPWR VPWR
+ _02843_ sky130_fd_sc_hd__or3b_1
XFILLER_0_43_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06244__A2 _01190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08067_ _01660_ _02773_ genblk1\[5\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _02774_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10904__S _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07018_ genblk1\[7\].osc.clkdiv_C.cnt\[12\] _01841_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10328__A1 _01735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09194__A1 _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07744__A2 _02425_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08969_ _03565_ _03567_ _03508_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__o21a_1
X_11980_ genblk2\[10\].wave_shpr.div.fin_quo\[7\] genblk2\[10\].wave_shpr.div.quo\[6\]
+ _00003_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06891__A2_N _01666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10931_ _02171_ net1234 VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13650_ clknet_leaf_38_clk _00963_ net116 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10862_ genblk2\[6\].wave_shpr.div.b1\[12\] genblk2\[6\].wave_shpr.div.acc\[12\]
+ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[4\] net97 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13581_ clknet_leaf_76_clk _00896_ net207 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10793_ net654 _04918_ _04922_ _04946_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12532_ clknet_leaf_61_clk _00084_ net186 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12463_ clknet_leaf_103_clk _00036_ net156 VGND VGND VPWR VPWR PWM.final_sample_in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11414_ genblk2\[8\].wave_shpr.div.b1\[8\] genblk2\[8\].wave_shpr.div.acc\[8\] VGND
+ VGND VPWR VPWR _05390_ sky130_fd_sc_hd__and2b_1
X_12394_ genblk2\[11\].wave_shpr.div.acc\[11\] _06067_ _06055_ VGND VGND VPWR VPWR
+ _06068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11345_ net1048 _05311_ _05315_ _05333_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11276_ _05185_ _05280_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__xnor2_1
X_13015_ clknet_leaf_12_clk _00010_ net52 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09185__A1 _01430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10227_ genblk2\[3\].wave_shpr.div.acc\[22\] _04416_ _04547_ VGND VGND VPWR VPWR
+ _04548_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07735__A2 _02433_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10158_ _04389_ _04373_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__or2b_1
XANTENNA_clkbuf_leaf_131_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3 _00951_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10089_ genblk2\[3\].wave_shpr.div.quo\[2\] _04452_ _04456_ net326 VGND VGND VPWR
+ VPWR _00377_ sky130_fd_sc_hd__a22o_1
XANTENNA__12330__A _03689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08145__C1 _01362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07143__B _01514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08954__S _02248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08448__B1 genblk2\[8\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06320_ genblk1\[0\].osc.clkdiv_C.cnt\[4\] _01276_ _01270_ VGND VGND VPWR VPWR _01278_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06251_ _01174_ _01187_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__nand2_2
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_60_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09785__S _04238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06182_ _01153_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11755__B1 _03694_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold403 _00640_ VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold414 genblk2\[1\].wave_shpr.div.quo\[24\] VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10724__S _04821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold425 genblk2\[4\].wave_shpr.div.acc_next\[0\] VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 genblk2\[5\].wave_shpr.div.acc\[22\] VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold447 genblk2\[4\].wave_shpr.div.quo\[22\] VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 genblk2\[8\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09086__A modein.delay_octave_down_in\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09941_ net707 _04253_ _04322_ _04345_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__a22o_1
Xhold469 _00868_ VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09176__A1 _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07318__B _01262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _04293_ _04182_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10025__A _02170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _03465_ _03481_ _03480_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__o21a_1
Xhold1103 genblk2\[8\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net1321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 genblk2\[11\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net1332 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 genblk2\[2\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net1343 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ _03454_ _03460_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__xnor2_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ genblk2\[10\].wave_shpr.div.fin_quo\[6\] VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__inv_2
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _03387_ _03391_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11286__A2 _05279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_92_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08149__B _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08151__A2 _01250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _02337_ _02341_ _02342_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__or3b_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07567_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01936_ _01349_ VGND VGND VPWR VPWR _02274_
+ sky130_fd_sc_hd__o21a_1
X_09306_ genblk2\[0\].wave_shpr.div.acc\[8\] _03892_ _03889_ VGND VGND VPWR VPWR _03893_
+ sky130_fd_sc_hd__mux2_1
X_06518_ genblk1\[2\].osc.clkdiv_C.cnt\[9\] _01442_ _01439_ genblk1\[2\].osc.clkdiv_C.cnt\[5\]
+ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_8_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07498_ _02218_ _02219_ VGND VGND VPWR VPWR FSM.next_mode\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_118_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09237_ net584 _03845_ _03839_ net599 _03846_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06449_ genblk1\[1\].osc.clkdiv_C.cnt\[6\] _01385_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09168_ _03810_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11746__B1 _05624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08119_ _02822_ _02823_ _02824_ _02825_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__o31a_1
XFILLER_0_32_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09099_ genblk2\[0\].wave_shpr.div.acc\[16\] genblk2\[0\].wave_shpr.div.b1\[16\]
+ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__or2b_1
XFILLER_0_102_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07965__A2 _01577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11130_ _05179_ _05189_ _05177_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold970 genblk2\[4\].wave_shpr.div.b1\[4\] VGND VGND VPWR VPWR net1188 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06413__A genblk1\[1\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold981 genblk2\[10\].wave_shpr.div.b1\[12\] VGND VGND VPWR VPWR net1199 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ _05016_ _04966_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__or2b_1
Xhold992 _00891_ VGND VGND VPWR VPWR net1210 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06132__B net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10012_ _04364_ _04406_ _04407_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__a21o_1
XANTENNA__08390__A2 _01442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11963_ genblk2\[10\].wave_shpr.div.acc\[24\] _05784_ VGND VGND VPWR VPWR _05785_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_83_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_16
X_13702_ clknet_leaf_97_clk _01013_ net167 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10914_ _05041_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06153__A1 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11894_ net348 _03696_ _03694_ _05721_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__a22o_1
X_13633_ clknet_leaf_69_clk _00946_ net213 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10845_ _04980_ _04987_ _04988_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10776_ net828 _04918_ _04922_ _04934_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13564_ clknet_leaf_57_clk _00879_ net182 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12515_ clknet_leaf_106_clk _00024_ net154 VGND VGND VPWR VPWR sig_norm.busy sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13495_ clknet_leaf_88_clk _00812_ net178 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12446_ clknet_leaf_99_clk net219 net168 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12377_ _05981_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07956__A2 _02656_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11328_ genblk2\[7\].wave_shpr.div.acc\[14\] _05320_ _05300_ VGND VGND VPWR VPWR
+ _05321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11259_ genblk2\[7\].wave_shpr.div.quo\[23\] _05245_ _05249_ net487 _05269_ VGND
+ VGND VPWR VPWR _00734_ sky130_fd_sc_hd__a221o_1
XANTENNA__12940__RESET_B net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08381__A2 _01209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11268__A2 _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_74_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_16
X_08470_ genblk2\[5\].wave_shpr.div.fin_quo\[0\] genblk2\[5\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07421_ genblk2\[2\].wave_shpr.div.busy _02162_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07352_ _02092_ _02109_ _02110_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06303_ genblk1\[0\].osc.clkdiv_C.cnt\[14\] _01256_ _01258_ genblk1\[0\].osc.clkdiv_C.cnt\[5\]
+ _01264_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07283_ genblk1\[10\].osc.clkdiv_C.cnt\[12\] _02052_ VGND VGND VPWR VPWR _02053_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_73_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09022_ _03693_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__clkbuf_4
X_06234_ _01195_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09809__A _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold200 genblk2\[4\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold211 _00062_ VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__dlygate4sd3_1
X_06165_ _01134_ _01136_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold222 genblk2\[10\].wave_shpr.div.quo\[19\] VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold233 genblk2\[3\].wave_shpr.div.quo\[18\] VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 genblk2\[1\].wave_shpr.div.quo\[16\] VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _00507_ VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 genblk2\[7\].wave_shpr.div.b1\[14\] VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 genblk2\[0\].wave_shpr.div.quo\[13\] VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 genblk2\[8\].wave_shpr.div.quo\[11\] VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ genblk2\[2\].wave_shpr.div.acc\[17\] _04333_ _04213_ VGND VGND VPWR VPWR
+ _04334_ sky130_fd_sc_hd__mux2_1
Xhold299 genblk2\[1\].wave_shpr.div.quo\[9\] VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _04214_ _04280_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__nand2_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11285__S _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08806_ _03433_ _03437_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__or2b_1
XANTENNA__09263__B genblk1\[0\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09786_ _04243_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__clkbuf_1
X_06998_ _01823_ _01829_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07580__B1 genblk1\[9\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08737_ _03442_ _03441_ _03439_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11259__A2 _05245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_65_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08124__A2 _01340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _02838_ _03374_ _02846_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__o21a_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07619_ genblk1\[11\].osc.clkdiv_C.cnt\[5\] _01595_ _02323_ _02324_ _02325_ VGND
+ VGND VPWR VPWR _02326_ sky130_fd_sc_hd__o221a_1
X_08599_ net9 _02744_ _03305_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__and3_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ net1308 _02725_ _04834_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__mux2_1
XANTENNA__09085__B1 _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10561_ _04778_ _04788_ _04776_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12300_ genblk2\[11\].wave_shpr.div.quo\[1\] _06009_ _06010_ net430 VGND VGND VPWR
+ VPWR _01034_ sky130_fd_sc_hd__a22o_1
X_13280_ clknet_leaf_122_clk _00601_ net79 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_51_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10492_ net926 _04715_ _04722_ _04734_ VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12231_ genblk2\[11\].wave_shpr.div.b1\[14\] genblk2\[11\].wave_shpr.div.acc\[14\]
+ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__and2b_1
XFILLER_0_122_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11195__A1 _05236_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07938__A2 _02539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12162_ genblk2\[10\].wave_shpr.div.acc\[22\] _05908_ VGND VGND VPWR VPWR _05909_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06143__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11113_ genblk2\[7\].wave_shpr.div.acc\[8\] genblk2\[7\].wave_shpr.div.b1\[8\] VGND
+ VGND VPWR VPWR _05173_ sky130_fd_sc_hd__or2b_1
X_12093_ _05756_ _05742_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__nor2_1
XANTENNA__06610__A2 _01231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11044_ net883 _05119_ _05093_ _05122_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__a22o_1
XANTENNA__08899__B1 _01157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09560__A1 _03819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09173__B _01441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06374__B2 genblk1\[1\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12995_ clknet_leaf_131_clk _00324_ net64 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_56_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08115__A2 _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11946_ genblk2\[10\].wave_shpr.div.b1\[11\] genblk2\[10\].wave_shpr.div.acc\[11\]
+ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08520__C1 _02364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11877_ genblk2\[9\].wave_shpr.div.acc\[20\] _05707_ VGND VGND VPWR VPWR _05710_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13616_ clknet_leaf_94_clk _00929_ net160 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10828_ genblk2\[6\].wave_shpr.div.acc\[11\] genblk2\[6\].wave_shpr.div.b1\[11\]
+ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__or2b_1
XFILLER_0_82_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08236__C _02365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13547_ clknet_leaf_109_clk _00862_ net152 VGND VGND VPWR VPWR sig_norm.b1\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10759_ net981 _04918_ _04890_ _04921_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13478_ clknet_leaf_99_clk _00795_ net168 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12429_ genblk2\[11\].wave_shpr.div.acc\[20\] _06092_ VGND VGND VPWR VPWR _06094_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11186__A1 _01508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07970_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01577_ _02668_ VGND VGND VPWR VPWR _02677_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06921_ _01761_ _01768_ _01769_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
X_09640_ net983 _04109_ _04113_ _04132_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__a22o_1
X_06852_ genblk1\[5\].osc.clkdiv_C.cnt\[10\] _01710_ genblk1\[5\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09083__B _01201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09571_ net965 _04076_ _04047_ _04079_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__a22o_1
X_06783_ net851 _01654_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_16
X_08522_ _02416_ _03228_ net2 _02364_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07314__B1 genblk1\[11\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08453_ _02684_ _02681_ _02687_ _02526_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__o31a_1
XFILLER_0_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout152_A net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07404_ genblk2\[0\].wave_shpr.div.busy _02149_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__and2_1
X_08384_ _01437_ genblk1\[2\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07335_ genblk1\[11\].osc.clkdiv_C.cnt\[2\] genblk1\[11\].osc.clkdiv_C.cnt\[1\] genblk1\[11\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07266_ genblk1\[10\].osc.clkdiv_C.cnt\[6\] _02039_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__nor2_1
X_09005_ net1151 VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06217_ _01178_ _01176_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__nor2_4
XFILLER_0_103_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07197_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01981_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06148_ _01118_ _01108_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__and2b_1
XANTENNA__10924__A1 _02374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08593__A2 _02526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09790__A1 _03714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09907_ genblk2\[2\].wave_shpr.div.acc\[13\] _04320_ _04301_ VGND VGND VPWR VPWR
+ _04321_ sky130_fd_sc_hd__mux2_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09838_ net261 _04257_ _04259_ net656 _04270_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__a221o_1
XANTENNA__06356__A1 genblk1\[0\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout65_A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09769_ _04234_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_38_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ net1022 _05623_ _05624_ _05651_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__a22o_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ clknet_leaf_40_clk _00113_ net116 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11731_ _05618_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__clkbuf_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10359__S _04637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ genblk2\[9\].wave_shpr.div.acc\[17\] genblk2\[9\].wave_shpr.div.b1\[17\]
+ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__or2b_1
X_13401_ clknet_leaf_92_clk _00720_ net143 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10613_ genblk2\[6\].wave_shpr.div.b1\[1\] _04831_ _04637_ VGND VGND VPWR VPWR _04832_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11593_ genblk2\[8\].wave_shpr.div.acc\[10\] _05505_ _05493_ VGND VGND VPWR VPWR
+ _05506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10544_ genblk2\[5\].wave_shpr.div.acc\[8\] genblk2\[5\].wave_shpr.div.b1\[8\] VGND
+ VGND VPWR VPWR _04772_ sky130_fd_sc_hd__or2b_1
X_13332_ clknet_leaf_9_clk net284 net54 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13263_ clknet_leaf_0_clk _00586_ net38 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10475_ net901 _04715_ _04690_ _04721_ VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12214_ _05937_ _05950_ _05951_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__a21o_1
X_13194_ clknet_leaf_127_clk _00517_ net67 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09230__B1 _03839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12145_ _05779_ _05896_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09184__A _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12076_ _05812_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__clkbuf_4
X_11027_ net806 _05086_ _05093_ _05109_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06898__A2 _01367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12978_ clknet_leaf_124_clk net316 net72 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07432__A _02170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11929_ _05745_ _05749_ _05750_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07120_ _01432_ _01221_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07051_ _01336_ _01183_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__nor2_2
XFILLER_0_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12356__B1 _06010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09221__B1 _03840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09772__A1 _01256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10732__S _04821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10382__A2 _04657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09094__A _01367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07953_ genblk1\[7\].osc.clkdiv_C.cnt\[2\] _01732_ _02656_ genblk1\[7\].osc.clkdiv_C.cnt\[3\]
+ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__o22a_1
XANTENNA__08327__A2 _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06904_ _01576_ _01757_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__nand2_2
X_07884_ genblk2\[1\].wave_shpr.div.fin_quo\[6\] _02590_ VGND VGND VPWR VPWR _02591_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__10134__A2 _04451_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07535__B1 _01099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09623_ net905 _04109_ _04113_ _04119_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__a22o_1
X_06835_ net1105 _01700_ _01702_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__11563__S _05417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06766_ _01643_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[12\] sky130_fd_sc_hd__clkbuf_1
X_09554_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__and2_1
X_08505_ genblk2\[2\].wave_shpr.div.fin_quo\[5\] _03113_ _03118_ _02224_ VGND VGND
+ VPWR VPWR _03212_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09485_ _04031_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06697_ genblk1\[4\].osc.clkdiv_C.cnt\[1\] _01436_ _01304_ genblk1\[4\].osc.clkdiv_C.cnt\[7\]
+ _01586_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08436_ genblk2\[11\].wave_shpr.div.fin_quo\[2\] _02349_ _02351_ _02352_ VGND VGND
+ VPWR VPWR _03143_ sky130_fd_sc_hd__nand4_1
XFILLER_0_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08367_ _03072_ _03073_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10907__S _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07318_ genblk1\[11\].osc.clkdiv_C.cnt\[11\] _01262_ VGND VGND VPWR VPWR _02082_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07066__A2 _01578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08298_ _02969_ _03003_ _03004_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06274__B1 _01235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07249_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] genblk1\[10\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _02030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10260_ genblk2\[4\].wave_shpr.div.acc\[10\] genblk2\[4\].wave_shpr.div.b1\[10\]
+ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10191_ net1017 _04518_ _04490_ _04521_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__a22o_1
XANTENNA__10642__S _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06421__A _01336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_896 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07526__B1 _01099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12901_ clknet_leaf_30_clk net589 net102 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ clknet_leaf_64_clk _00165_ net189 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12763_ clknet_leaf_20_clk _00096_ net108 VGND VGND VPWR VPWR freq_div.state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_96_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11714_ genblk2\[9\].wave_shpr.div.b1\[17\] genblk2\[9\].wave_shpr.div.acc\[17\]
+ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__and2b_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12694_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[7\] net172 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11645_ _05414_ genblk2\[8\].wave_shpr.div.acc\[25\] genblk2\[8\].wave_shpr.div.acc\[26\]
+ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__or3b_1
XFILLER_0_140_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07057__A2 _01246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput15 pb[9] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_4
XANTENNA__08083__A _02225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11576_ _05416_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__clkbuf_4
X_13315_ clknet_leaf_9_clk net516 net48 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10527_ genblk2\[4\].wave_shpr.div.i\[1\] genblk2\[4\].wave_shpr.div.i\[0\] genblk2\[4\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__and3_1
XANTENNA__06804__A2 _01362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10458_ net928 _04683_ _04690_ _04708_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__a22o_1
X_13246_ clknet_leaf_11_clk net494 net56 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_149_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13177_ clknet_leaf_130_clk _00502_ net65 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10389_ net675 _04661_ _04655_ net602 _04662_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__a221o_1
XANTENNA__07765__B1 _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12128_ _05772_ _05735_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__or2b_1
X_12059_ _03833_ _02023_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06620_ _01524_ _01525_ _01526_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__and3_1
X_06551_ _01451_ _01466_ _01467_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_59_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09270_ genblk2\[0\].wave_shpr.div.b1\[0\] _03804_ genblk2\[0\].wave_shpr.div.acc\[0\]
+ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__a21oi_1
X_06482_ genblk1\[1\].osc.clkdiv_C.cnt\[17\] _01407_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08221_ _02793_ _02789_ genblk2\[5\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR
+ _02928_ sky130_fd_sc_hd__or3b_1
XFILLER_0_7_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_894 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08152_ genblk1\[3\].osc.clkdiv_C.cnt\[5\] _01500_ _01250_ genblk1\[3\].osc.clkdiv_C.cnt\[4\]
+ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__o22a_1
XANTENNA__07048__A2 _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10052__A1 _01870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07103_ _01887_ _01908_ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_4_3_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08083_ _02225_ _02789_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07034_ genblk1\[8\].osc.clkdiv_C.cnt\[15\] _01359_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11001__B1 _05056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08440__B _02403_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08985_ _03669_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07936_ _02637_ _02638_ _02641_ genblk2\[8\].wave_shpr.div.fin_quo\[6\] VGND VGND
+ VPWR VPWR _02643_ sky130_fd_sc_hd__a31o_1
XANTENNA__07056__B _01498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07867_ _02469_ _02573_ _02529_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__o21a_1
XANTENNA__11293__S _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06895__B _01362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09606_ _03992_ _03960_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06818_ _01669_ _01559_ _01675_ genblk1\[5\].osc.clkdiv_C.cnt\[14\] _01689_ VGND
+ VGND VPWR VPWR _01690_ sky130_fd_sc_hd__o221a_1
X_07798_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] genblk1\[0\].osc.clkdiv_C.cnt\[14\] _01209_
+ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09537_ genblk2\[1\].wave_shpr.div.quo\[15\] _04052_ _04053_ net511 _04059_ VGND
+ VGND VPWR VPWR _00222_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06749_ _01630_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09468_ _03732_ net1047 _03733_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08419_ _03001_ _03078_ _03055_ _03077_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10637__S _04834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09399_ genblk2\[1\].wave_shpr.div.acc\[8\] genblk2\[1\].wave_shpr.div.b1\[8\] VGND
+ VGND VPWR VPWR _03963_ sky130_fd_sc_hd__or2b_1
XFILLER_0_34_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11430_ _05243_ genblk2\[8\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR _05406_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_117_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06416__A _01359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10043__A1 _03732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11361_ _05220_ _05248_ _05344_ _05251_ net1029 VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10312_ genblk2\[4\].wave_shpr.div.fin_quo\[0\] _04623_ _00013_ VGND VGND VPWR VPWR
+ _04624_ sky130_fd_sc_hd__mux2_1
X_13100_ clknet_leaf_136_clk _00427_ net42 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11292_ _05192_ _05292_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__xnor2_1
X_13031_ clknet_leaf_122_clk _00358_ net79 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10243_ _04454_ _04557_ _04558_ _04457_ net1079 VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__a32o_1
X_10174_ net796 _04486_ _04490_ _04508_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__a22o_1
Xfanout170 net171 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__buf_2
Xfanout181 net185 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_4
Xfanout192 net193 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10401__A _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12815_ clknet_leaf_58_clk net579 net192 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10806__B1 _04855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12746_ clknet_leaf_49_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[5\] net108 VGND VGND
+ VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12677_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[8\] net142 VGND VGND
+ VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__12328__A _03689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11628_ genblk2\[8\].wave_shpr.div.acc\[19\] _05531_ VGND VGND VPWR VPWR _05532_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__12023__A2 _05813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11559_ genblk2\[8\].wave_shpr.div.acc\[2\] _05479_ _05417_ VGND VGND VPWR VPWR _05480_
+ sky130_fd_sc_hd__mux2_1
Xhold607 genblk2\[1\].wave_shpr.div.acc\[5\] VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07986__B1 _02527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold618 genblk2\[2\].wave_shpr.div.acc\[7\] VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold629 genblk2\[1\].wave_shpr.div.acc\[9\] VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13229_ clknet_leaf_15_clk _00552_ net56 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07157__A genblk1\[9\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _03454_ _03475_ _03476_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__o21ai_2
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11298__B1 _05283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07721_ genblk1\[1\].osc.clkdiv_C.cnt\[13\] _02425_ _02426_ _02427_ VGND VGND VPWR
+ VPWR _02428_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12002__S _05802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07652_ _02316_ _02357_ _02358_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__or3b_1
XFILLER_0_79_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06603_ _01486_ _01487_ _01492_ _01504_ _01510_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07583_ genblk1\[9\].osc.clkdiv_C.cnt\[2\] _01234_ _02287_ _02288_ _02289_ VGND VGND
+ VPWR VPWR _02290_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09322_ _03786_ _03904_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06534_ genblk1\[2\].osc.clkdiv_C.cnt\[3\] _01454_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_861 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06465_ genblk1\[1\].osc.clkdiv_C.cnt\[11\] genblk1\[1\].osc.clkdiv_C.cnt\[10\] _01394_
+ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__and3_1
X_09253_ _03855_ _01169_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__nor2_1
XANTENNA__10457__S _04704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12635__RESET_B net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08204_ _02303_ _02265_ genblk2\[9\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR
+ _02911_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09184_ _03719_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06396_ _01238_ _01262_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__nor2_4
XFILLER_0_90_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06236__A _01174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08135_ genblk2\[4\].wave_shpr.div.fin_quo\[4\] _02841_ VGND VGND VPWR VPWR _02842_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11222__B1 _05250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10981__A _05074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08066_ _01179_ _01222_ _01254_ _01171_ genblk1\[5\].osc.clkdiv_C.cnt\[0\] VGND VGND
+ VPWR VPWR _02773_ sky130_fd_sc_hd__o311a_1
X_07017_ _01822_ _01840_ _01841_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_3_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06401__B1 _01344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10920__S _05042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08968_ _03655_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__clkbuf_1
X_07919_ genblk1\[8\].osc.clkdiv_C.cnt\[7\] _01430_ _01858_ genblk1\[8\].osc.clkdiv_C.cnt\[5\]
+ _02625_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__a221o_1
X_08899_ _03574_ _03600_ _03603_ _01157_ net1069 VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__a32o_1
X_10930_ _03726_ _05049_ _03736_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07901__B1 _01328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10861_ _04972_ _05003_ _05004_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12600_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[3\] net97 VGND VGND
+ VPWR VPWR genblk1\[3\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_149_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13580_ clknet_leaf_76_clk _00895_ net207 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10792_ _04817_ _04880_ _04943_ genblk2\[5\].wave_shpr.div.acc\[21\] VGND VGND VPWR
+ VPWR _04946_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_66_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12531_ clknet_leaf_61_clk _00083_ net186 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12462_ clknet_leaf_104_clk _00035_ net155 VGND VGND VPWR VPWR PWM.final_sample_in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11413_ _05368_ _05387_ _05388_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12393_ _05962_ _06066_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11344_ _05331_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11275_ _05186_ _05181_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__or2b_1
XFILLER_0_30_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13014_ clknet_leaf_132_clk _00343_ net60 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09185__A2 _01344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10226_ _04417_ _04418_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__and2b_1
XANTENNA__07196__A1 genblk1\[9\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10157_ net963 _04486_ _04490_ _04495_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__a22o_1
Xhold4 modein.delay_in\[0\] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_2
X_10088_ net326 _04452_ _04456_ net794 VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__a22o_1
XANTENNA__11227__A _05074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07424__B _02153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12729_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[6\] net115 VGND VGND
+ VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06250_ genblk1\[0\].osc.clkdiv_C.cnt\[0\] _01211_ _01210_ genblk1\[0\].osc.clkdiv_C.cnt\[15\]
+ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11204__B1 _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06181_ sig_norm.busy _01152_ _01098_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07959__B1 _01925_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold404 genblk2\[6\].wave_shpr.div.acc\[19\] VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11755__B2 net526 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold415 _00231_ VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 _00484_ VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 genblk2\[0\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold448 _00481_ VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ genblk2\[2\].wave_shpr.div.acc\[22\] _04343_ VGND VGND VPWR VPWR _04345_
+ sky130_fd_sc_hd__xnor2_1
Xhold459 genblk2\[8\].wave_shpr.div.quo\[19\] VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _04183_ _04168_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__or2b_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _03464_ _03526_ _03528_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__or3_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 genblk2\[0\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net1322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 genblk2\[4\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net1333 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 genblk2\[5\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net1344 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ _03457_ _03459_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout182_A net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07704_ _02404_ _02405_ genblk2\[10\].wave_shpr.div.fin_quo\[6\] _02410_ VGND VGND
+ VPWR VPWR _02411_ sky130_fd_sc_hd__and4b_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _03114_ _03390_ _03122_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07635_ genblk1\[11\].osc.clkdiv_C.cnt\[9\] _01190_ _01235_ genblk1\[11\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__o22a_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07566_ _02269_ _02271_ _02272_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09041__S _03708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09305_ _03778_ _03891_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__xnor2_1
X_06517_ genblk1\[2\].osc.clkdiv_C.cnt\[5\] _01439_ _01442_ genblk1\[2\].osc.clkdiv_C.cnt\[9\]
+ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_36_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07497_ _02217_ _02215_ net760 VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__or3_1
XANTENNA__08165__B _01508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09236_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__and2_1
X_06448_ _01373_ _01385_ _01386_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_106_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09167_ genblk2\[0\].wave_shpr.div.fin_quo\[5\] net1334 _00001_ VGND VGND VPWR VPWR
+ _03810_ sky130_fd_sc_hd__mux2_1
X_06379_ _01322_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08118_ genblk1\[4\].osc.clkdiv_C.cnt\[2\] _01326_ _01213_ genblk1\[4\].osc.clkdiv_C.cnt\[3\]
+ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09098_ _03734_ genblk2\[0\].wave_shpr.div.acc\[17\] VGND VGND VPWR VPWR _03746_
+ sky130_fd_sc_hd__or2_1
X_08049_ genblk1\[5\].osc.clkdiv_C.cnt\[11\] _01355_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__nor2_1
Xhold960 genblk2\[4\].wave_shpr.div.b1\[6\] VGND VGND VPWR VPWR net1178 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06413__B _01356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold971 genblk1\[7\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR net1189 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout95_A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11060_ net899 _05119_ _05126_ _05134_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__a22o_1
Xhold982 genblk2\[7\].wave_shpr.div.b1\[4\] VGND VGND VPWR VPWR net1200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold993 genblk2\[6\].wave_shpr.div.b1\[7\] VGND VGND VPWR VPWR net1211 sky130_fd_sc_hd__dlygate4sd3_1
X_10011_ genblk2\[3\].wave_shpr.div.b1\[14\] genblk2\[3\].wave_shpr.div.acc\[14\]
+ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11962_ genblk2\[10\].wave_shpr.div.acc\[23\] genblk2\[10\].wave_shpr.div.acc\[22\]
+ genblk2\[10\].wave_shpr.div.acc\[21\] _05783_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__or4_1
XFILLER_0_99_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13701_ clknet_leaf_99_clk _01012_ net166 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06689__B1 _01578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10913_ net1201 _01819_ _04848_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__mux2_1
X_11893_ genblk2\[9\].wave_shpr.div.acc\[25\] _05719_ VGND VGND VPWR VPWR _05721_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13632_ clknet_leaf_69_clk _00945_ net213 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10844_ genblk2\[6\].wave_shpr.div.b1\[3\] genblk2\[6\].wave_shpr.div.acc\[3\] VGND
+ VGND VPWR VPWR _04988_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_11_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13563_ clknet_leaf_57_clk net244 net184 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10775_ genblk2\[5\].wave_shpr.div.acc\[16\] _04933_ _04907_ VGND VGND VPWR VPWR
+ _04934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12514_ clknet_leaf_106_clk _00025_ net153 VGND VGND VPWR VPWR PWM.start sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13494_ clknet_leaf_86_clk _00811_ net178 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12445_ net960 _03947_ _03944_ _06104_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12376_ _05954_ _06053_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06604__A _01171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11327_ _05208_ _05319_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11258_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__and2_1
X_10209_ _04413_ _04361_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__or2b_1
X_11189_ _05234_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10712__A2 _04853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08118__B1 _01213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07420_ genblk2\[2\].wave_shpr.div.i\[1\] _02161_ genblk2\[2\].wave_shpr.div.i\[4\]
+ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__or3b_1
XFILLER_0_147_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07170__A genblk1\[9\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07351_ genblk1\[11\].osc.clkdiv_C.cnt\[4\] genblk1\[11\].osc.clkdiv_C.cnt\[3\] _02097_
+ genblk1\[11\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06302_ genblk1\[0\].osc.clkdiv_C.cnt\[12\] _01263_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07282_ _02027_ _02051_ _02052_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06233_ _01194_ _01175_ _01191_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__nor3_1
X_09021_ _03692_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06164_ _01133_ _01135_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__nand2_1
Xhold201 _00460_ VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold212 genblk2\[11\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 genblk2\[2\].wave_shpr.div.quo\[10\] VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _00393_ VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__C1 genblk1\[0\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold245 _00223_ VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 genblk2\[10\].wave_shpr.div.quo\[22\] VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 genblk2\[9\].wave_shpr.div.quo\[14\] VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _00137_ VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _04206_ _04332_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09825__A _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold289 genblk2\[5\].wave_shpr.div.quo\[18\] VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10470__S _04704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09854_ _04174_ _04175_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__xnor2_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09544__B genblk1\[1\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _03511_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__inv_2
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ genblk2\[3\].wave_shpr.div.b1\[14\] _04242_ _04238_ VGND VGND VPWR VPWR _04243_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06997_ genblk1\[7\].osc.clkdiv_C.cnt\[4\] _01827_ VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07580__A1 _01432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08736_ _03439_ _03441_ _03442_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__nand3b_2
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ _03372_ _03373_ genblk2\[4\].wave_shpr.div.fin_quo\[3\] _02362_ VGND VGND
+ VPWR VPWR _03374_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ genblk1\[11\].osc.clkdiv_C.cnt\[4\] _02064_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ genblk2\[3\].wave_shpr.div.fin_quo\[0\] _02592_ _02467_ genblk2\[3\].wave_shpr.div.fin_quo\[1\]
+ _02939_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09085__A1 _03714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07549_ net1157 net1132 PWM.start VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10560_ _04779_ _04786_ _04787_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07635__A2 _01190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_130_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09219_ _03838_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10645__S _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10491_ genblk2\[4\].wave_shpr.div.acc\[16\] _04733_ _04704_ VGND VGND VPWR VPWR
+ _04734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12230_ _05929_ _05966_ _05967_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06424__A _01365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12161_ genblk2\[10\].wave_shpr.div.acc\[21\] _05783_ _05899_ VGND VGND VPWR VPWR
+ _05908_ sky130_fd_sc_hd__or3_1
XANTENNA__07239__B _01215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10942__A2 _05052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11112_ genblk2\[7\].wave_shpr.div.acc\[9\] genblk2\[7\].wave_shpr.div.b1\[9\] VGND
+ VGND VPWR VPWR _05172_ sky130_fd_sc_hd__or2b_1
XANTENNA__10047__A1_N _03727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12092_ net977 _05844_ _05850_ _05856_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__a22o_1
Xhold790 genblk2\[4\].wave_shpr.div.acc\[11\] VGND VGND VPWR VPWR net1008 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11043_ genblk2\[6\].wave_shpr.div.acc\[12\] _05121_ _05105_ VGND VGND VPWR VPWR
+ _05122_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06374__A2 _01311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12994_ clknet_leaf_131_clk _00323_ net64 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11945_ _05738_ _05765_ _05766_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08520__B1 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11505__A _05441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11876_ genblk2\[9\].wave_shpr.div.acc\[20\] _05707_ VGND VGND VPWR VPWR _05709_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_28_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13615_ clknet_leaf_94_clk _00928_ net160 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09076__A1 _01483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10827_ genblk2\[6\].wave_shpr.div.acc\[12\] genblk2\[6\].wave_shpr.div.b1\[12\]
+ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__or2b_1
XFILLER_0_67_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13546_ clknet_leaf_109_clk _00861_ net152 VGND VGND VPWR VPWR sig_norm.b1\[0\] sky130_fd_sc_hd__dfrtp_1
X_10758_ genblk2\[5\].wave_shpr.div.acc\[12\] _04920_ _04907_ VGND VGND VPWR VPWR
+ _04921_ sky130_fd_sc_hd__mux2_1
XANTENNA__07626__A2 _01241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13597__RESET_B net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13477_ clknet_leaf_72_clk _00794_ net216 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10689_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__and2_1
XANTENNA__12336__A _03689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12428_ net1203 _06072_ _06073_ _06093_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12359_ _05947_ _05939_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__or2b_1
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06920_ genblk1\[6\].osc.clkdiv_C.cnt\[4\] _01765_ genblk1\[6\].osc.clkdiv_C.cnt\[5\]
+ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12071__A _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06851_ genblk1\[5\].osc.clkdiv_C.cnt\[10\] _01710_ _01712_ _01694_ VGND VGND VPWR
+ VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o211a_1
XANTENNA__11894__B1 _03694_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09551__A2 _04042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09083__C _01363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12479__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06500__C net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09570_ genblk2\[1\].wave_shpr.div.acc\[2\] _04078_ _04011_ VGND VGND VPWR VPWR _04079_
+ sky130_fd_sc_hd__mux2_1
X_06782_ _01655_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[16\] sky130_fd_sc_hd__clkbuf_1
X_08521_ _02216_ _02552_ genblk2\[10\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR
+ _03228_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08452_ _02682_ _02687_ _02684_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07403_ genblk2\[0\].wave_shpr.div.i\[1\] _02148_ genblk2\[0\].wave_shpr.div.i\[4\]
+ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__or3b_1
XFILLER_0_148_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08383_ _03087_ _03088_ _03089_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout145_A net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06228__B _01189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07334_ _02096_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07617__A2 _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07265_ genblk1\[10\].osc.clkdiv_C.cnt\[6\] _02039_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__and2_1
XANTENNA__10465__S _04704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13267__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09004_ net1150 sig_norm.quo\[3\] _01154_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__mux2_1
X_06216_ freq_div.state\[1\] VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__buf_4
X_07196_ genblk1\[9\].osc.clkdiv_C.cnt\[13\] _01979_ _01982_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__o21a_1
X_06147_ net1 net7 _01118_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09906_ _04198_ _04319_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__xnor2_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _04269_ genblk1\[2\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__and2_1
XANTENNA__10213__B _04480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ genblk2\[3\].wave_shpr.div.b1\[6\] _01262_ _04039_ VGND VGND VPWR VPWR _04234_
+ sky130_fd_sc_hd__mux2_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout58_A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _03420_ _03421_ _03383_ _03395_ VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__o211a_1
XANTENNA__07803__A net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ genblk2\[2\].wave_shpr.div.b1\[3\] genblk2\[2\].wave_shpr.div.acc\[3\] VGND
+ VGND VPWR VPWR _04179_ sky130_fd_sc_hd__and2b_1
XFILLER_0_69_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11730_ genblk2\[9\].wave_shpr.div.fin_quo\[4\] genblk2\[9\].wave_shpr.div.quo\[3\]
+ _00023_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__mux2_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07856__A2 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06419__A _01362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ net319 _05552_ _05553_ VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__a21oi_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13400_ clknet_leaf_119_clk net422 net143 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10612_ _01738_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11592_ _05393_ _05504_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13331_ clknet_leaf_24_clk _00652_ net92 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10543_ genblk2\[5\].wave_shpr.div.acc\[9\] genblk2\[5\].wave_shpr.div.b1\[9\] VGND
+ VGND VPWR VPWR _04771_ sky130_fd_sc_hd__or2b_1
XFILLER_0_107_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08281__A2 _02521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13262_ clknet_leaf_0_clk _00585_ net38 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10474_ genblk2\[4\].wave_shpr.div.acc\[12\] _04720_ _04704_ VGND VGND VPWR VPWR
+ _04721_ sky130_fd_sc_hd__mux2_1
X_12213_ genblk2\[11\].wave_shpr.div.b1\[5\] genblk2\[11\].wave_shpr.div.acc\[5\]
+ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13193_ clknet_leaf_118_clk _00516_ net138 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12144_ _05780_ _05731_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__or2b_1
XFILLER_0_138_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06595__A2 _01363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07792__A1 _01246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12075_ _05842_ _05843_ net1118 _05813_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__a2bb2o_1
X_11026_ genblk2\[6\].wave_shpr.div.acc\[8\] _05108_ _05105_ VGND VGND VPWR VPWR _05109_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12977_ clknet_leaf_123_clk _00306_ net72 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11235__A _05074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11928_ genblk2\[10\].wave_shpr.div.b1\[2\] genblk2\[10\].wave_shpr.div.acc\[2\]
+ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11859_ genblk2\[9\].wave_shpr.div.acc\[15\] _05696_ _05673_ VGND VGND VPWR VPWR
+ _05697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13529_ clknet_leaf_98_clk _00846_ net169 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11800__B1 _05624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07050_ genblk1\[8\].osc.clkdiv_C.cnt\[9\] _01865_ _01867_ VGND VGND VPWR VPWR _01868_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_51_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07232__B1 _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07783__A1 _01200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07952_ genblk1\[7\].osc.clkdiv_C.cnt\[0\] _01801_ _02657_ _02658_ VGND VGND VPWR
+ VPWR _02659_ sky130_fd_sc_hd__a31o_1
X_06903_ _01325_ _01327_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__nor2_2
X_07883_ _02464_ genblk2\[1\].wave_shpr.div.fin_quo\[5\] _02461_ VGND VGND VPWR VPWR
+ _02590_ sky130_fd_sc_hd__or3b_1
X_09622_ genblk2\[1\].wave_shpr.div.acc\[14\] _04118_ _04095_ VGND VGND VPWR VPWR
+ _04119_ sky130_fd_sc_hd__mux2_1
X_06834_ genblk1\[5\].osc.clkdiv_C.cnt\[4\] _01700_ _01694_ VGND VGND VPWR VPWR _01702_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09553_ genblk2\[1\].wave_shpr.div.quo\[23\] _04042_ _04046_ net340 _04067_ VGND
+ VGND VPWR VPWR _00230_ sky130_fd_sc_hd__a221o_1
X_06765_ _01599_ _01640_ _01642_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08504_ _03113_ _03118_ genblk2\[2\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR
+ _03211_ sky130_fd_sc_hd__a21oi_1
X_09484_ genblk2\[2\].wave_shpr.div.b1\[9\] _01302_ _04024_ VGND VGND VPWR VPWR _04031_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07838__A2 _02539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06239__A _01200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06696_ genblk1\[4\].osc.clkdiv_C.cnt\[3\] _01326_ _01574_ genblk1\[4\].osc.clkdiv_C.cnt\[12\]
+ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08435_ net33 _02350_ _02352_ genblk2\[11\].wave_shpr.div.fin_quo\[2\] VGND VGND
+ VPWR VPWR _03142_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08366_ _02938_ _02944_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08454__A _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07317_ genblk1\[11\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__inv_2
XANTENNA__10195__S _04507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08297_ _03002_ _02970_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__and2b_1
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08173__B _01858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07248_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] genblk1\[10\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _02029_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10358__B1 _04647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07179_ _01971_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[7\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__07223__B1 _01196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10190_ genblk2\[3\].wave_shpr.div.acc\[12\] _04520_ _04507_ VGND VGND VPWR VPWR
+ _04521_ sky130_fd_sc_hd__mux2_1
XANTENNA__06702__A _01171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09515__A2 _04043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12900_ clknet_leaf_30_clk net633 net102 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07533__A _02248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12831_ clknet_leaf_64_clk _00164_ net189 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ clknet_leaf_20_clk _00095_ net109 VGND VGND VPWR VPWR freq_div.state\[1\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11713_ _05555_ _05603_ _05604_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__o21bai_2
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[6\] net172 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11644_ net1052 _05448_ _05445_ _05542_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput16 reset VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08254__A2 _02733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11575_ _05385_ _05491_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08083__B _02789_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13314_ clknet_leaf_12_clk _00635_ net54 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10526_ genblk2\[4\].wave_shpr.div.i\[1\] genblk2\[4\].wave_shpr.div.i\[0\] genblk2\[4\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__a21o_1
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13245_ clknet_leaf_11_clk net325 net54 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09203__A1 _01302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10457_ genblk2\[4\].wave_shpr.div.acc\[8\] _04707_ _04704_ VGND VGND VPWR VPWR _04708_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08006__A2 _01735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07708__A _02225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13176_ clknet_leaf_130_clk _00501_ net65 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10388_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__and2_1
XANTENNA__07765__A1 genblk1\[0\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07765__B2 genblk1\[0\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12127_ _05815_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__clkbuf_4
X_12058_ net383 _05823_ _05825_ net440 _05833_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__a221o_1
X_11009_ genblk2\[6\].wave_shpr.div.acc\[4\] _05095_ _05023_ VGND VGND VPWR VPWR _05096_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10521__A0 _04654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06689__A2_N _01574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06550_ genblk1\[2\].osc.clkdiv_C.cnt\[9\] _01464_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06481_ genblk1\[1\].osc.clkdiv_C.cnt\[16\] _01405_ _01408_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[16\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08220_ _02925_ _02926_ _02897_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12026__B1 _05817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08151_ genblk1\[3\].osc.clkdiv_C.cnt\[4\] _01250_ _01514_ genblk1\[3\].osc.clkdiv_C.cnt\[3\]
+ _02857_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07102_ genblk1\[8\].osc.clkdiv_C.cnt\[12\] genblk1\[8\].osc.clkdiv_C.cnt\[11\] _01904_
+ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__and3_1
XANTENNA__06256__A1 genblk1\[0\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08082_ _02784_ _02788_ genblk1\[5\].osc.clkdiv_C.cnt\[16\] genblk1\[5\].osc.clkdiv_C.cnt\[17\]
+ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__a211o_4
XFILLER_0_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07033_ net848 _01850_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout108_A net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08984_ net1156 _03668_ _01158_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09833__A _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07935_ _02637_ genblk2\[8\].wave_shpr.div.fin_quo\[6\] _02638_ _02641_ _02223_ VGND
+ VGND VPWR VPWR _02642_ sky130_fd_sc_hd__a41o_1
XANTENNA__10979__A _05074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09552__B genblk1\[1\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07866_ net17 _02552_ genblk2\[1\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR
+ _02573_ sky130_fd_sc_hd__and3_1
X_09605_ net366 _04076_ _04080_ _04105_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__a22o_1
X_06817_ _01681_ _01686_ _01687_ _01688_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__and4bb_1
X_07797_ _02493_ _02500_ _02502_ _02498_ _02503_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__a32oi_1
XANTENNA__07072__B genblk1\[8\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09536_ _04058_ _01307_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__nor2_1
X_06748_ _01599_ _01628_ _01629_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09467_ _04021_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__clkbuf_1
X_06679_ genblk1\[4\].osc.clkdiv_C.cnt\[15\] _01363_ _01242_ _01568_ genblk1\[4\].osc.clkdiv_C.cnt\[17\]
+ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__a221o_1
XANTENNA__10918__S _05042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08418_ _03083_ _03124_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09398_ genblk2\[1\].wave_shpr.div.acc\[9\] genblk2\[1\].wave_shpr.div.b1\[9\] VGND
+ VGND VPWR VPWR _03962_ sky130_fd_sc_hd__or2b_1
XANTENNA__08184__A _02225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08349_ _02789_ _02792_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11360_ _05342_ _05343_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10311_ _04622_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_132_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11291_ _05193_ _05175_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__or2b_1
XFILLER_0_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13030_ clknet_leaf_122_clk _00357_ net79 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10242_ genblk2\[3\].wave_shpr.div.i\[1\] genblk2\[3\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _04558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10173_ genblk2\[3\].wave_shpr.div.acc\[8\] _04506_ _04507_ VGND VGND VPWR VPWR _04508_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout160 net162 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_4
Xfanout171 net16 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_4
Xfanout182 net185 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__buf_2
Xfanout193 net195 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_2
XFILLER_0_97_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12814_ clknet_leaf_58_clk net455 net192 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ clknet_leaf_50_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[4\] net108 VGND VGND
+ VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[7\] net82 VGND VGND
+ VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_72_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11627_ genblk2\[8\].wave_shpr.div.acc\[18\] _05529_ VGND VGND VPWR VPWR _05531_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11558_ _05377_ _05478_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold608 genblk2\[6\].wave_shpr.div.acc\[7\] VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__dlygate4sd3_1
X_10509_ genblk2\[4\].wave_shpr.div.acc\[22\] _04657_ _04722_ _04746_ VGND VGND VPWR
+ VPWR _00507_ sky130_fd_sc_hd__a22o_1
Xhold619 genblk1\[6\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__buf_1
XFILLER_0_111_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12344__A genblk2\[11\].wave_shpr.div.acc_next\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11489_ _02171_ net1239 VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__and2_1
XANTENNA__09188__B1 _03705_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13228_ clknet_leaf_125_clk net309 net69 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ clknet_leaf_121_clk net644 net78 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07157__B genblk1\[9\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07720_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] _01309_ _01208_ genblk1\[1\].osc.clkdiv_C.cnt\[14\]
+ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07651_ _02349_ _02351_ _02356_ genblk2\[11\].wave_shpr.div.fin_quo\[6\] VGND VGND
+ VPWR VPWR _02358_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06602_ genblk1\[3\].osc.clkdiv_C.cnt\[0\] _01484_ _01505_ _01506_ _01509_ VGND VGND
+ VPWR VPWR _01510_ sky130_fd_sc_hd__a221o_1
X_07582_ genblk1\[9\].osc.clkdiv_C.cnt\[1\] _01230_ _01221_ VGND VGND VPWR VPWR _02289_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_149_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09321_ _03787_ _03751_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06533_ genblk1\[2\].osc.clkdiv_C.cnt\[3\] _01454_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11470__A1 _01946_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09252_ _03719_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__buf_6
X_06464_ genblk1\[1\].osc.clkdiv_C.cnt\[10\] _01394_ genblk1\[1\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08203_ _02901_ _02905_ _02909_ _02419_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09183_ _03818_ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06395_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] _01210_ _01337_ genblk1\[1\].osc.clkdiv_C.cnt\[12\]
+ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08134_ genblk2\[4\].wave_shpr.div.fin_quo\[3\] _02840_ VGND VGND VPWR VPWR _02841_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_71_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08065_ _02770_ _02771_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07016_ genblk1\[7\].osc.clkdiv_C.cnt\[11\] genblk1\[7\].osc.clkdiv_C.cnt\[10\] _01837_
+ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07729__A1 _01360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06401__A1 _01342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06401__B2 genblk1\[1\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08967_ sig_norm.quo\[6\] _03654_ _00024_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__mux2_1
X_07918_ _01489_ genblk1\[8\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__xor2_1
X_08898_ _03581_ _03601_ net26 VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__a21o_1
X_07849_ _02461_ _02462_ genblk2\[1\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR
+ _02556_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07901__B2 genblk1\[8\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10860_ genblk2\[6\].wave_shpr.div.b1\[11\] genblk2\[6\].wave_shpr.div.acc\[11\]
+ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout40_A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09519_ _04042_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__clkbuf_4
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10791_ net566 _04918_ _04922_ _04945_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ clknet_leaf_61_clk _00082_ net188 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12461_ clknet_leaf_104_clk _00034_ net155 VGND VGND VPWR VPWR PWM.final_sample_in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11412_ genblk2\[8\].wave_shpr.div.b1\[7\] genblk2\[8\].wave_shpr.div.acc\[7\] VGND
+ VGND VPWR VPWR _05388_ sky130_fd_sc_hd__and2b_1
X_12392_ _05963_ _05931_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__or2b_1
XFILLER_0_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11343_ _05216_ _05273_ genblk2\[7\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR
+ _05332_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06162__A net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11274_ _05245_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13013_ clknet_leaf_133_clk _00342_ net60 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10225_ net710 _04518_ _04522_ _04546_ VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__a22o_1
X_10156_ genblk2\[3\].wave_shpr.div.acc\[4\] _04494_ _04420_ VGND VGND VPWR VPWR _04495_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11508__A _05444_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold5 genblk2\[10\].wave_shpr.div.quo\[11\] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dlygate4sd3_1
X_10087_ _04455_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10412__A _04672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08145__A1 _01201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10989_ genblk2\[6\].wave_shpr.div.acc\[0\] _00016_ _05079_ net283 _05080_ VGND VGND
+ VPWR VPWR _00653_ sky130_fd_sc_hd__o221a_1
XFILLER_0_57_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12728_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[5\] net113 VGND VGND
+ VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12659_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[8\] net90 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06180_ sig_norm.i\[1\] sig_norm.i\[0\] sig_norm.i\[3\] _01151_ VGND VGND VPWR VPWR
+ _01152_ sky130_fd_sc_hd__and4_1
XFILLER_0_25_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11755__A2 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold405 genblk2\[6\].wave_shpr.div.quo\[11\] VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 genblk2\[3\].wave_shpr.div.quo\[14\] VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold427 genblk2\[1\].wave_shpr.div.quo\[11\] VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 genblk2\[2\].wave_shpr.div.quo\[20\] VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 genblk2\[4\].wave_shpr.div.b1\[16\] VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ net919 _04282_ _04289_ _04292_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__a22o_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _03473_ _03527_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__or2_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1105 genblk2\[10\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net1323 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06395__B1 _01337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 genblk2\[0\].wave_shpr.div.quo\[4\] VGND VGND VPWR VPWR net1334 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1127 genblk2\[5\].wave_shpr.div.acc\[20\] VGND VGND VPWR VPWR net1345 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ _02950_ _03458_ _02647_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__a21oi_1
X_07703_ genblk2\[10\].wave_shpr.div.fin_quo\[4\] _02409_ VGND VGND VPWR VPWR _02410_
+ sky130_fd_sc_hd__nor2_1
X_08683_ _03388_ _03389_ genblk2\[2\].wave_shpr.div.fin_quo\[3\] _02468_ VGND VGND
+ VPWR VPWR _03390_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_45_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07634_ genblk1\[11\].osc.clkdiv_C.cnt\[9\] _01190_ _02339_ _02340_ VGND VGND VPWR
+ VPWR _02341_ sky130_fd_sc_hd__a211o_1
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07565_ genblk1\[9\].osc.clkdiv_C.cnt\[12\] _01328_ _01799_ genblk1\[9\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__a22oi_1
X_09304_ _03779_ _03755_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__or2b_1
X_06516_ _01200_ _01441_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__nand2_4
XFILLER_0_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07496_ _02215_ net760 _02217_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06247__A _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_810 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09235_ _03835_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__clkbuf_4
X_06447_ genblk1\[1\].osc.clkdiv_C.cnt\[4\] _01380_ genblk1\[1\].osc.clkdiv_C.cnt\[5\]
+ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09166_ _03809_ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__clkbuf_1
X_06378_ net37 _01321_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11746__A2 _05623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08117_ genblk1\[4\].osc.clkdiv_C.cnt\[2\] _01326_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09097_ _03745_ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08181__B _02885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07078__A genblk1\[8\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08048_ _02752_ _02754_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold950 PWM.final_in\[5\] VGND VGND VPWR VPWR net1168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 smpl_rt_clkdiv.clkDiv_inst.cnt\[6\] VGND VGND VPWR VPWR net1179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 genblk2\[3\].wave_shpr.div.b1\[17\] VGND VGND VPWR VPWR net1190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 genblk2\[7\].wave_shpr.div.b1\[8\] VGND VGND VPWR VPWR net1201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 genblk2\[5\].wave_shpr.div.b1\[3\] VGND VGND VPWR VPWR net1212 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10010_ _04365_ _04404_ _04405_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout88_A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07499__B_N net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09999_ genblk2\[3\].wave_shpr.div.b1\[8\] genblk2\[3\].wave_shpr.div.acc\[8\] VGND
+ VGND VPWR VPWR _04395_ sky130_fd_sc_hd__and2b_1
X_11961_ genblk2\[10\].wave_shpr.div.acc\[20\] genblk2\[10\].wave_shpr.div.acc\[19\]
+ _05782_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__or3_1
X_13700_ clknet_leaf_97_clk _01011_ net166 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10912_ _05040_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__clkbuf_1
X_11892_ net1045 _03696_ _03694_ _05720_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13631_ clknet_leaf_66_clk _00944_ net197 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10843_ _04981_ genblk2\[6\].wave_shpr.div.acc\[2\] _04986_ VGND VGND VPWR VPWR _04987_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__09088__C1 _03738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13562_ clknet_leaf_85_clk _00877_ net184 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10774_ _04932_ _04811_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12513_ clknet_leaf_84_clk _00075_ net202 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13493_ clknet_leaf_86_clk net238 net177 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12444_ _06102_ _06103_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11510__B genblk1\[8\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12375_ _05955_ _05935_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10407__A _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10945__B1 _05056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06604__B _01192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11326_ _05209_ _05167_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__or2b_1
XFILLER_0_10_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11257_ net487 _05245_ _05249_ net542 _05268_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__a221o_1
X_10208_ net948 _04518_ _04522_ _04534_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__a22o_1
XANTENNA__09563__B1 _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11188_ genblk2\[8\].wave_shpr.div.b1\[6\] _01507_ _05042_ VGND VGND VPWR VPWR _05234_
+ sky130_fd_sc_hd__mux2_1
X_10139_ genblk2\[3\].wave_shpr.div.b1\[0\] _04420_ genblk2\[3\].wave_shpr.div.acc\[0\]
+ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10228__A2 _04457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07170__B genblk1\[9\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07350_ _02108_ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__inv_2
X_06301_ _01238_ _01262_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__or2_4
XFILLER_0_128_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07281_ genblk1\[10\].osc.clkdiv_C.cnt\[11\] genblk1\[10\].osc.clkdiv_C.cnt\[10\]
+ _02048_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09020_ _02152_ genblk2\[9\].wave_shpr.div.busy _02201_ VGND VGND VPWR VPWR _03692_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_115_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06232_ freq_div.state\[0\] VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__buf_2
XFILLER_0_127_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06163_ _01130_ _01132_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12008__S _05802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold202 genblk2\[11\].wave_shpr.div.b1\[8\] VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 _01034_ VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _00302_ VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 genblk2\[5\].wave_shpr.div.quo\[12\] VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 genblk2\[4\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 _00972_ VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 genblk2\[6\].wave_shpr.div.quo\[18\] VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 sig_norm.b1\[1\] VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ _04207_ _04156_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__or2b_1
X_09853_ genblk2\[2\].wave_shpr.div.acc\[1\] _04213_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__or2_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _03442_ _03443_ _03217_ _03510_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__a211oi_2
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _01490_ _01233_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__nor2_4
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ _01823_ _01827_ _01828_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__07580__A2 _01221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08735_ _03405_ _03406_ _03202_ _03440_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__a211o_1
XANTENNA__09841__A _04269_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10987__A _05054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ genblk2\[4\].wave_shpr.div.fin_quo\[2\] _02932_ _02839_ _02316_ VGND VGND
+ VPWR VPWR _03373_ sky130_fd_sc_hd__a31o_1
XFILLER_0_68_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07617_ genblk1\[11\].osc.clkdiv_C.cnt\[3\] _01513_ _02064_ genblk1\[11\].osc.clkdiv_C.cnt\[4\]
+ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__a22o_1
X_08597_ _03302_ _03303_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__nor2_1
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07548_ net1169 VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07479_ genblk2\[10\].wave_shpr.div.i\[2\] genblk2\[10\].wave_shpr.div.i\[3\] genblk2\[10\].wave_shpr.div.i\[0\]
+ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_146_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09218_ net804 _03836_ _03804_ _03839_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10490_ _04732_ _04613_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06705__A _01489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09149_ _03734_ genblk2\[0\].wave_shpr.div.acc\[17\] VGND VGND VPWR VPWR _03797_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06424__B _01367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12160_ net1257 _05818_ _05883_ _05907_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11111_ genblk2\[7\].wave_shpr.div.acc\[10\] genblk2\[7\].wave_shpr.div.b1\[10\]
+ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__or2b_1
X_12091_ genblk2\[10\].wave_shpr.div.acc\[4\] _05855_ _05787_ VGND VGND VPWR VPWR
+ _05856_ sky130_fd_sc_hd__mux2_1
Xhold780 genblk2\[4\].wave_shpr.div.acc\[6\] VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold791 genblk2\[7\].wave_shpr.div.acc\[8\] VGND VGND VPWR VPWR net1009 sky130_fd_sc_hd__dlygate4sd3_1
X_11042_ _05005_ _05120_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09751__A _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12993_ clknet_leaf_131_clk _00322_ net64 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11944_ genblk2\[10\].wave_shpr.div.b1\[10\] genblk2\[10\].wave_shpr.div.acc\[10\]
+ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11875_ net935 _05684_ _05685_ _05708_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10826_ genblk2\[6\].wave_shpr.div.acc\[13\] genblk2\[6\].wave_shpr.div.b1\[13\]
+ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__or2b_1
X_13614_ clknet_leaf_94_clk _00927_ net159 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_95_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10757_ _04803_ _04919_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__xnor2_1
X_13545_ clknet_leaf_101_clk _00860_ net165 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_133_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_133_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10091__B1 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13476_ clknet_leaf_72_clk _00793_ net216 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10688_ genblk2\[5\].wave_shpr.div.quo\[18\] _04861_ _04862_ net235 _04871_ VGND
+ VGND VPWR VPWR _00561_ sky130_fd_sc_hd__a221o_1
XFILLER_0_124_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12427_ genblk2\[11\].wave_shpr.div.acc\[19\] _06089_ _06092_ VGND VGND VPWR VPWR
+ _06093_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12358_ _03941_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11309_ _05200_ _05305_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__xnor2_1
X_12289_ _06006_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07446__A _02147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06850_ genblk1\[5\].osc.clkdiv_C.cnt\[10\] _01710_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06781_ _01599_ _01653_ _01654_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08520_ _03141_ _03226_ net3 _02364_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__o211ai_2
XANTENNA__07314__A2 _02077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08451_ _02636_ _03157_ _02604_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07402_ genblk2\[0\].wave_shpr.div.i\[2\] genblk2\[0\].wave_shpr.div.i\[3\] genblk2\[0\].wave_shpr.div.i\[0\]
+ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08382_ genblk1\[2\].osc.clkdiv_C.cnt\[2\] _02336_ _01418_ genblk1\[2\].osc.clkdiv_C.cnt\[3\]
+ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09600__S _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07333_ _02092_ _02094_ _02095_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_124_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_124_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout138_A net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07264_ _02027_ _02039_ _02040_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_45_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09003_ _03681_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06215_ _01175_ _01176_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_115_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07195_ _01953_ _01981_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06146_ net11 _01105_ _01104_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09836__A _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13236__RESET_B net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09905_ _04199_ _04160_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__or2b_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ _04268_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__buf_2
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ _03704_ net1099 _04233_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__a21o_1
X_06979_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01363_ _01196_ _01813_ _01814_ VGND
+ VGND VPWR VPWR _01815_ sky130_fd_sc_hd__o221a_1
XFILLER_0_69_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _03383_ _03395_ _03420_ _03421_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__a211oi_2
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _04171_ genblk2\[2\].wave_shpr.div.acc\[2\] _04177_ VGND VGND VPWR VPWR _04178_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _03353_ _03355_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__xnor2_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ net319 _05552_ _03855_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10611_ _04830_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_115_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_115_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11591_ _05394_ _05365_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13330_ clknet_leaf_24_clk net386 net91 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10542_ genblk2\[5\].wave_shpr.div.acc\[10\] genblk2\[5\].wave_shpr.div.b1\[10\]
+ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__or2b_1
XFILLER_0_52_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13261_ clknet_leaf_0_clk _00584_ net38 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10473_ _04605_ _04719_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12212_ _05938_ _05948_ _05949_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__a21o_1
X_13192_ clknet_leaf_122_clk _00515_ net79 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09230__A2 _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12143_ net859 _05876_ _05883_ _05895_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12117__A2 _05844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09518__B1 _04047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07792__A2 _01439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12074_ genblk2\[10\].wave_shpr.div.b1\[0\] genblk2\[10\].wave_shpr.div.acc\[0\]
+ _05787_ _05840_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__a31o_1
X_11025_ _04997_ _05107_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07633__A2_N _01262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11516__A _05441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10420__A _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12976_ clknet_leaf_123_clk net458 net71 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11927_ _05746_ _05747_ _05748_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__a21o_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ _05601_ _05695_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_106_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_106_clk sky130_fd_sc_hd__clkbuf_16
X_10809_ genblk2\[5\].wave_shpr.div.i\[1\] genblk2\[5\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _04957_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11789_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13528_ clknet_leaf_98_clk _00845_ net169 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13459_ clknet_leaf_99_clk _00776_ net166 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12356__A2 _06009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09221__A2 _03836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11564__B1 _05446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08980__A1 _01157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07951_ genblk1\[7\].osc.clkdiv_C.cnt\[1\] _01556_ _01564_ _01732_ genblk1\[7\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06902_ _01741_ _01744_ _01746_ _01755_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__or4_1
XFILLER_0_128_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07882_ _02547_ _02586_ _02520_ _02587_ _02588_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__a2111oi_1
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09621_ _03997_ _04117_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__xnor2_1
X_06833_ _01693_ _01700_ _01701_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__07904__A genblk1\[8\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09552_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__and2_1
X_06764_ _01641_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08503_ _03196_ _03199_ _03209_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12292__A1 _01327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09483_ _04030_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06695_ genblk1\[4\].osc.clkdiv_C.cnt\[10\] _01323_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__nor2_1
X_08434_ _02349_ _02351_ _02221_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_148_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08365_ _03042_ _03047_ _03041_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_117_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07316_ genblk1\[11\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__inv_2
X_08296_ _02970_ _03002_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06274__A2 _01227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07247_ _02026_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12347__A2 _05982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07178_ _01954_ _01969_ _01970_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__and3_1
XANTENNA__10358__A1 _03704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06129_ net13 net15 VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__nand2_1
XANTENNA__07223__A1 _01174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06702__B _01591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07086__A genblk1\[8\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11307__B1 _05283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout70_A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07814__A _02308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09819_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__and2_1
X_12830_ clknet_leaf_62_clk _00163_ net189 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ clknet_leaf_20_clk _00094_ net108 VGND VGND VPWR VPWR freq_div.state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12283__A1 _01946_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _05439_ genblk2\[9\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR _05604_
+ sky130_fd_sc_hd__and2_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ clknet_leaf_53_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[5\] net172 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _05540_ _05413_ genblk2\[8\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR
+ _05542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11574_ _05386_ _05369_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__or2b_1
XFILLER_0_25_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13313_ clknet_leaf_121_clk net242 net78 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10525_ _04655_ _04755_ _04756_ _04657_ net1108 VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13244_ clknet_leaf_9_clk _00567_ net54 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10456_ _04597_ _04706_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10349__A1 _01757_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11546__B1 _05444_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13175_ clknet_leaf_129_clk _00500_ net67 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07708__B _02403_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10387_ _04651_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__buf_2
XANTENNA__10415__A _04676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06612__B _01519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11204__A2_N _01490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12126_ net858 _05876_ _05850_ _05882_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__a22o_1
XANTENNA__07765__A2 _01309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06973__B1 _01311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12057_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR _05833_
+ sky130_fd_sc_hd__and2_1
X_11008_ _05094_ _04989_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10521__A1 _04651_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10150__A _04455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12959_ clknet_leaf_136_clk _00288_ net42 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06480_ net29 _01407_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__nor2_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08150_ genblk1\[3\].osc.clkdiv_C.cnt\[3\] _01234_ _02854_ _02855_ _02856_ VGND VGND
+ VPWR VPWR _02857_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09089__C _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07101_ genblk1\[8\].osc.clkdiv_C.cnt\[11\] _01904_ _01907_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__o21a_1
X_08081_ _02752_ _02753_ _02755_ _02786_ _02787_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06256__A2 _01210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07032_ _01851_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07618__B _02064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08983_ sig_norm.quo\[8\] _01098_ _03667_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__a21bo_1
X_07934_ genblk2\[8\].wave_shpr.div.fin_quo\[4\] _02640_ VGND VGND VPWR VPWR _02641_
+ sky130_fd_sc_hd__nor2_1
X_07865_ _02216_ _02552_ genblk2\[0\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR
+ _02572_ sky130_fd_sc_hd__and3_1
XANTENNA__06796__A2_N _01666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09604_ genblk2\[1\].wave_shpr.div.acc\[10\] _04104_ _04095_ VGND VGND VPWR VPWR
+ _04105_ sky130_fd_sc_hd__mux2_1
X_06816_ genblk1\[5\].osc.clkdiv_C.cnt\[12\] _01355_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__or2_1
X_07796_ _02496_ _02497_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire30 _02635_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
X_06747_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] genblk1\[4\].osc.clkdiv_C.cnt\[6\] _01616_
+ genblk1\[4\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__a31o_1
X_09535_ _03719_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__buf_4
XANTENNA__12265__A1 _01240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10995__A _05023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09466_ net1247 _01327_ _03822_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06678_ genblk1\[4\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__inv_2
XANTENNA__06684__S _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08417_ _03085_ _03123_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__xnor2_1
X_09397_ genblk2\[1\].wave_shpr.div.acc\[10\] genblk2\[1\].wave_shpr.div.b1\[10\]
+ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__or2b_1
XFILLER_0_108_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08184__B _02885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08348_ _03054_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08279_ genblk2\[9\].wave_shpr.div.fin_quo\[4\] _02303_ _02264_ _02223_ VGND VGND
+ VPWR VPWR _02986_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10310_ genblk2\[4\].wave_shpr.div.acc\[25\] genblk2\[4\].wave_shpr.div.acc\[24\]
+ genblk2\[4\].wave_shpr.div.acc\[26\] _04621_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__or4b_4
XFILLER_0_62_899 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07995__A2 _01484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11290_ net988 _05279_ _05283_ _05291_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__a22o_1
X_10241_ genblk2\[3\].wave_shpr.div.i\[1\] genblk2\[3\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _04557_ sky130_fd_sc_hd__or2_1
X_10172_ _04419_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__buf_4
Xfanout150 net171 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_4
Xfanout161 net162 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__buf_2
Xfanout172 net173 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_4
Xfanout183 net185 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_4
Xfanout194 net195 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08172__A2 _01498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06183__A1 _01099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12813_ clknet_leaf_58_clk _00146_ net192 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10806__A2 _04858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12744_ clknet_leaf_49_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[3\] net108 VGND VGND
+ VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07132__B1 _01349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12008__A1 _01483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ clknet_leaf_90_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[6\] net141 VGND VGND
+ VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_53_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11626_ net1114 _05507_ _05445_ _05530_ VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11557_ _05378_ _05373_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__or2b_1
XFILLER_0_108_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10508_ net472 _04744_ _04745_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__a21o_1
Xhold609 genblk2\[1\].wave_shpr.div.acc\[8\] VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11488_ _03726_ _05439_ _03736_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09188__A1 _03714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10439_ _04580_ _04590_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__xor2_1
X_13227_ clknet_leaf_127_clk _00550_ net67 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10145__A _04451_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ clknet_leaf_121_clk _00483_ net78 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ net1035 _05844_ _05850_ _05869_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__a22o_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13089_ clknet_leaf_137_clk _00416_ net40 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07454__A _02147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11298__A2 _05279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08163__A2 _01498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07650_ genblk2\[11\].wave_shpr.div.fin_quo\[6\] _02349_ _02351_ _02356_ VGND VGND
+ VPWR VPWR _02357_ sky130_fd_sc_hd__and4_1
X_06601_ genblk1\[3\].osc.clkdiv_C.cnt\[12\] _01507_ _01508_ genblk1\[3\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07910__A2 _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07581_ _01186_ _01437_ _01226_ _01171_ genblk1\[9\].osc.clkdiv_C.cnt\[0\] VGND VGND
+ VPWR VPWR _02288_ sky130_fd_sc_hd__o311a_1
X_09320_ _03835_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06532_ _01452_ _01454_ _01455_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_88_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09251_ genblk2\[0\].wave_shpr.div.quo\[18\] _03845_ _03847_ net410 _03854_ VGND
+ VGND VPWR VPWR _00141_ sky130_fd_sc_hd__a221o_1
X_06463_ genblk1\[1\].osc.clkdiv_C.cnt\[10\] _01394_ _01396_ _01374_ VGND VGND VPWR
+ VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o211a_1
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08202_ _02906_ _02907_ _02908_ _02416_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09182_ net1273 _01214_ _03722_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06394_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] _01210_ _01337_ genblk1\[1\].osc.clkdiv_C.cnt\[12\]
+ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_43_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08133_ genblk2\[4\].wave_shpr.div.fin_quo\[2\] _02839_ VGND VGND VPWR VPWR _02840_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_55_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11222__A2 _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout218_A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08064_ genblk1\[5\].osc.clkdiv_C.cnt\[3\] _01195_ _01254_ VGND VGND VPWR VPWR _02771_
+ sky130_fd_sc_hd__or3_1
XANTENNA__07629__A _01174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07015_ genblk1\[7\].osc.clkdiv_C.cnt\[10\] _01837_ genblk1\[7\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06252__B _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07729__A2 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_wire33_A _02348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06401__A2 genblk1\[1\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08966_ sig_norm.quo\[5\] _03653_ _01155_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__mux2_1
X_07917_ genblk1\[8\].osc.clkdiv_C.cnt\[5\] _01858_ _02621_ _02622_ _02623_ VGND VGND
+ VPWR VPWR _02624_ sky130_fd_sc_hd__o221a_1
X_08897_ sig_norm.acc\[11\] sig_norm.acc\[12\] _03591_ _03594_ VGND VGND VPWR VPWR
+ _03602_ sky130_fd_sc_hd__nor4_2
Xclkbuf_leaf_95_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_16
X_07848_ _02509_ _02551_ _02554_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__or3_1
XANTENNA__07901__A2 _01246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07779_ _01181_ genblk1\[0\].osc.clkdiv_C.cnt\[7\] _02485_ VGND VGND VPWR VPWR _02486_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09518_ net460 _04043_ _04047_ genblk2\[1\].wave_shpr.div.quo\[7\] VGND VGND VPWR
+ VPWR _00215_ sky130_fd_sc_hd__a22o_1
X_10790_ _04943_ _04944_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09449_ _04012_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__clkbuf_1
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12460_ clknet_leaf_104_clk _00033_ net155 VGND VGND VPWR VPWR PWM.final_sample_in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11749__B1 _05624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11411_ _05369_ _05385_ _05386_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12391_ net785 _06039_ _06040_ _06065_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11342_ _05217_ _05273_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11273_ net1013 _05246_ _05250_ _05278_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__a22o_1
X_10224_ _04416_ _04480_ _04543_ net524 VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__a2bb2o_1
X_13012_ clknet_leaf_133_clk _00341_ net60 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09754__A _01436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10155_ _04376_ _04387_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold6 _00961_ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dlygate4sd3_1
X_10086_ _04453_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_86_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10988_ _03719_ genblk1\[6\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12727_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[4\] net113 VGND VGND
+ VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10660__B1 _04857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12658_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[7\] net90 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_154_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11609_ _05401_ _05517_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12589_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[10\] net72 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_10_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07959__A2 _01311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold406 _00639_ VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 _00389_ VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold428 genblk2\[9\].wave_shpr.div.acc\[22\] VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 genblk2\[3\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _03470_ _03472_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06395__B2 genblk1\[1\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 genblk2\[10\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net1324 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 genblk2\[8\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net1335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1128 genblk2\[3\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net1346 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ genblk2\[7\].wave_shpr.div.fin_quo\[0\] _02467_ VGND VGND VPWR VPWR _03458_
+ sky130_fd_sc_hd__nand2_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07615__C _01437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_77_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_136_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07702_ _02406_ _02408_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__nand2_1
X_08682_ genblk2\[2\].wave_shpr.div.fin_quo\[2\] _03113_ _03115_ _02224_ VGND VGND
+ VPWR VPWR _03389_ sky130_fd_sc_hd__a31o_1
XFILLER_0_136_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07633_ genblk1\[11\].osc.clkdiv_C.cnt\[10\] _01262_ _01494_ _02128_ VGND VGND VPWR
+ VPWR _02340_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout168_A net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07564_ _01930_ _01227_ _01732_ _02268_ _02270_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__o221a_1
XANTENNA__07631__B _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09303_ net1049 _03870_ _03877_ _03890_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__a22o_1
X_06515_ _01440_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__buf_6
XFILLER_0_8_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07495_ _02216_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__buf_2
XFILLER_0_119_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09839__A _04269_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06446_ genblk1\[1\].osc.clkdiv_C.cnt\[5\] genblk1\[1\].osc.clkdiv_C.cnt\[4\] _01380_
+ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__and3_1
X_09234_ genblk2\[0\].wave_shpr.div.quo\[11\] _03841_ _03839_ net569 _03844_ VGND
+ VGND VPWR VPWR _00134_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09165_ genblk2\[0\].wave_shpr.div.fin_quo\[4\] genblk2\[0\].wave_shpr.div.quo\[3\]
+ _00001_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06377_ _01188_ _01191_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08116_ genblk1\[4\].osc.clkdiv_C.cnt\[1\] _01866_ genblk1\[4\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09096_ _03744_ _01490_ _03741_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08047_ genblk1\[5\].osc.clkdiv_C.cnt\[12\] _01666_ _02753_ VGND VGND VPWR VPWR _02754_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold940 genblk2\[0\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR net1158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold951 _02257_ VGND VGND VPWR VPWR net1169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 genblk1\[6\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR net1180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 genblk2\[8\].wave_shpr.div.b1\[17\] VGND VGND VPWR VPWR net1191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 genblk2\[7\].wave_shpr.div.b1\[6\] VGND VGND VPWR VPWR net1202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 genblk1\[2\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR net1213 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11903__B1 _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09998_ _04371_ _04392_ _04393_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__a21o_1
X_08949_ _03638_ _03639_ sig_norm.quo\[2\] _01098_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_leaf_68_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_16
X_11960_ genblk2\[10\].wave_shpr.div.acc\[18\] _05781_ VGND VGND VPWR VPWR _05782_
+ sky130_fd_sc_hd__or2_1
XANTENNA__08532__C1 _02364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07822__A net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10911_ genblk2\[7\].wave_shpr.div.b1\[7\] _04444_ _04848_ VGND VGND VPWR VPWR _05040_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07886__B2 _02592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11891_ _05718_ _05715_ _05719_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__o21ai_1
X_13630_ clknet_leaf_67_clk _00943_ net195 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10842_ _04981_ genblk2\[6\].wave_shpr.div.acc\[2\] _04985_ VGND VGND VPWR VPWR _04986_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09088__B1 _01591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07638__A1 _01229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13561_ clknet_leaf_85_clk _00876_ net184 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10773_ _04812_ _04764_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12512_ clknet_leaf_84_clk _00074_ net202 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13492_ clknet_leaf_87_clk _00809_ net177 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12443_ genblk2\[11\].wave_shpr.div.acc\[25\] _05980_ genblk2\[11\].wave_shpr.div.acc\[24\]
+ genblk2\[11\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__or4b_1
XFILLER_0_35_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11198__A1 _05239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12374_ net997 _06039_ _06040_ _06052_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06604__C _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11325_ net805 _05311_ _05315_ _05318_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__a22o_1
XANTENNA__06613__A2 _01256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_880 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11256_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09563__A1 _04045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10207_ genblk2\[3\].wave_shpr.div.acc\[16\] _04533_ _04507_ VGND VGND VPWR VPWR
+ _04534_ sky130_fd_sc_hd__mux2_1
X_11187_ _05233_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07574__B1 genblk1\[9\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10138_ _04480_ _04380_ genblk2\[3\].wave_shpr.div.b1\[0\] VGND VGND VPWR VPWR _04481_
+ sky130_fd_sc_hd__or3b_1
Xclkbuf_leaf_59_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08118__A2 _01326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10069_ net1205 _04444_ _04440_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__mux2_1
XANTENNA__08828__A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13759_ clknet_leaf_66_clk _01070_ net213 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_06300_ _01261_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__buf_4
XFILLER_0_127_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07280_ genblk1\[10\].osc.clkdiv_C.cnt\[10\] _02048_ genblk1\[10\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06231_ _01181_ _01192_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__nand2_2
XFILLER_0_122_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06162_ net10 VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold203 genblk2\[7\].wave_shpr.div.quo\[7\] VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold214 genblk2\[10\].wave_shpr.div.quo\[9\] VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 genblk2\[11\].wave_shpr.div.quo\[12\] VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 genblk2\[0\].wave_shpr.div.quo\[23\] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _00461_ VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06518__A2_N _01442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold258 genblk2\[0\].wave_shpr.div.quo\[22\] VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ net788 _04315_ _04322_ _04331_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__a22o_1
Xhold269 genblk2\[7\].wave_shpr.div.quo\[22\] VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08357__A2 _02521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09852_ _04277_ _04278_ net782 _04248_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__a2bb2o_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07565__B1 _01799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08803_ _03204_ _03205_ _03216_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__o21ba_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _03732_ net1152 _04241_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__o21a_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06995_ genblk1\[7\].osc.clkdiv_C.cnt\[3\] _01825_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__nor2_1
XANTENNA__08109__A2 _01323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08734_ _03202_ _03440_ _03405_ _03406_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__o211ai_2
XANTENNA__07642__A net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ _02932_ _02839_ genblk2\[4\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR
+ _03372_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10479__S _04704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _02318_ _02319_ _02320_ _02321_ _02322_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__o311a_1
XFILLER_0_49_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08596_ _02798_ _03299_ _03301_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__a21oi_1
X_07547_ PWM.final_sample_in\[5\] net1168 PWM.start VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07478_ _02204_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09217_ _03838_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__clkbuf_4
X_06429_ _01372_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06705__B _01196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09148_ _03747_ _03794_ _03795_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_860 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10927__A1 _01365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09079_ _03708_ _01210_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__nand2_8
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11110_ genblk2\[7\].wave_shpr.div.acc\[11\] genblk2\[7\].wave_shpr.div.b1\[11\]
+ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__or2b_1
X_12090_ _05854_ _05753_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__xnor2_1
Xhold770 genblk2\[7\].wave_shpr.div.acc\[6\] VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold781 genblk2\[9\].wave_shpr.div.acc\[5\] VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ _05006_ _04971_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__or2b_1
Xhold792 genblk2\[7\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR net1010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09751__B _01302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12992_ clknet_leaf_131_clk _00321_ net64 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12301__B1 _06010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold929_A genblk2\[8\].wave_shpr.div.b1\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11943_ _05739_ _05763_ _05764_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__a21o_1
X_11874_ genblk2\[9\].wave_shpr.div.acc\[19\] _05608_ _05707_ VGND VGND VPWR VPWR
+ _05708_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13613_ clknet_leaf_94_clk _00926_ net159 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10825_ genblk2\[6\].wave_shpr.div.acc\[14\] genblk2\[6\].wave_shpr.div.b1\[14\]
+ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__or2b_1
XANTENNA__11802__A _03693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13544_ clknet_leaf_101_clk _00859_ net164 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10756_ _04804_ _04768_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__or2b_1
XFILLER_0_82_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11521__B genblk1\[8\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13475_ clknet_leaf_71_clk _00792_ net216 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10687_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__and2_1
XANTENNA__11013__S _05023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12426_ _05978_ net20 VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__nor2_1
XANTENNA__08036__A1 genblk2\[6\].wave_shpr.div.fin_quo\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10918__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12357_ _03942_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11308_ _05201_ _05171_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__or2b_1
X_12288_ genblk2\[1\].wave_shpr.div.b1\[12\] _06005_ _05994_ VGND VGND VPWR VPWR _06006_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08339__A2 _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11239_ _05074_ genblk1\[7\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__and2_1
XANTENNA__11894__A2 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06780_ genblk1\[4\].osc.clkdiv_C.cnt\[16\] _01652_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08450_ _03155_ _03156_ genblk2\[8\].wave_shpr.div.fin_quo\[4\] _02521_ VGND VGND
+ VPWR VPWR _03157_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_147_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07401_ genblk2\[0\].wave_shpr.div.start VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__buf_8
XFILLER_0_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08381_ genblk1\[2\].osc.clkdiv_C.cnt\[1\] _01209_ _02336_ genblk1\[2\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07332_ genblk1\[11\].osc.clkdiv_C.cnt\[1\] genblk1\[11\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _02095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06806__A _01336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07263_ genblk1\[10\].osc.clkdiv_C.cnt\[4\] _02034_ genblk1\[10\].osc.clkdiv_C.cnt\[5\]
+ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09002_ net1172 net1176 _01154_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__mux2_1
X_06214_ freq_div.state\[2\] VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__buf_4
XANTENNA__09224__B1 _03840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07194_ genblk1\[9\].osc.clkdiv_C.cnt\[13\] genblk1\[9\].osc.clkdiv_C.cnt\[12\] _01978_
+ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__and3_1
XANTENNA__10909__A1 _04432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09775__A1 _02336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06145_ _01114_ _01116_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout200_A net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09904_ net953 _04315_ _04289_ _04318_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__a22o_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09835_ _02147_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__buf_4
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09766_ _01302_ _03727_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__nor2_4
X_06978_ genblk1\[7\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__inv_2
XANTENNA__09063__S _03722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08717_ _03386_ _03392_ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__nand2_1
XANTENNA__11098__B1 _05057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ _04171_ genblk2\[2\].wave_shpr.div.acc\[2\] _04176_ VGND VGND VPWR VPWR _04177_
+ sky130_fd_sc_hd__o21a_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08648_ _03280_ _03292_ _03354_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__a21oi_1
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08579_ _03285_ _02404_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__nor2_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10610_ genblk2\[6\].wave_shpr.div.b1\[0\] _01189_ _04637_ VGND VGND VPWR VPWR _04830_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11590_ net908 _05447_ _05484_ _05503_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10073__A1 _04242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10541_ genblk2\[5\].wave_shpr.div.acc\[11\] genblk2\[5\].wave_shpr.div.b1\[11\]
+ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__or2b_1
XFILLER_0_106_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13260_ clknet_leaf_0_clk _00583_ net38 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10472_ _04606_ _04570_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__or2b_1
X_12211_ genblk2\[11\].wave_shpr.div.b1\[4\] genblk2\[11\].wave_shpr.div.acc\[4\]
+ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13191_ clknet_leaf_122_clk net735 net78 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold879_A genblk2\[5\].wave_shpr.div.b1\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12142_ genblk2\[10\].wave_shpr.div.acc\[16\] _05894_ _05865_ VGND VGND VPWR VPWR
+ _05895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07792__A3 _01344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09518__B2 genblk2\[1\].wave_shpr.div.quo\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12073_ genblk2\[10\].wave_shpr.div.b1\[0\] _05787_ genblk2\[10\].wave_shpr.div.acc\[0\]
+ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__a21oi_1
X_11024_ _04998_ _04975_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__or2b_1
XANTENNA__11089__B1 _05055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12975_ clknet_leaf_124_clk _00304_ net71 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11926_ genblk2\[10\].wave_shpr.div.b1\[1\] genblk2\[10\].wave_shpr.div.acc\[1\]
+ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__and2b_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _05602_ _05556_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__or2b_1
XFILLER_0_129_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10808_ _04956_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11788_ net306 _02203_ _03693_ net565 _05643_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__a221o_1
XANTENNA__10064__A1 _01589_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11261__B1 _05249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13527_ clknet_leaf_98_clk _00844_ net169 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10739_ _04795_ _04905_ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11800__A2 _05623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13458_ clknet_leaf_99_clk _00775_ net165 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12409_ net897 _06072_ _06073_ _06079_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13389_ clknet_leaf_78_clk _00708_ net205 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07457__A _02189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06361__A _01223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07950_ _01556_ _01564_ genblk1\[7\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _02657_
+ sky130_fd_sc_hd__a21o_1
X_06901_ _01748_ _01749_ _01752_ _01754_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__or4_1
X_07881_ _02545_ _02518_ _02424_ _02541_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_128_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09620_ _03998_ _03957_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__or2b_1
XFILLER_0_37_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06832_ genblk1\[5\].osc.clkdiv_C.cnt\[3\] _01698_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__nor2_1
XANTENNA__07904__B _01869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09551_ net340 _04042_ _04046_ net608 _04066_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__a221o_1
X_06763_ genblk1\[4\].osc.clkdiv_C.cnt\[12\] _01637_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08502_ _03198_ _03197_ VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__and2b_1
X_09482_ genblk2\[2\].wave_shpr.div.b1\[8\] _01183_ _04024_ VGND VGND VPWR VPWR _04030_
+ sky130_fd_sc_hd__mux2_1
X_06694_ genblk1\[4\].osc.clkdiv_C.cnt\[11\] _01313_ _01561_ _01582_ _01583_ VGND
+ VGND VPWR VPWR _01584_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_66_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08433_ _02310_ _03139_ _02314_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout150_A net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08364_ _02846_ _03060_ _03064_ _03066_ _03070_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10055__A1 _04436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07315_ genblk1\[11\].osc.clkdiv_C.cnt\[8\] _01211_ _02077_ genblk1\[11\].osc.clkdiv_C.cnt\[12\]
+ _02078_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__o221a_1
X_08295_ _02998_ _03001_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09847__A _04250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07246_ net1080 _02027_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__08751__A genblk2\[7\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07177_ genblk1\[9\].osc.clkdiv_C.cnt\[7\] _01967_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__or2_1
XANTENNA__07759__B1 _02224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06128_ net13 net15 VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07504__B_N net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09818_ _04250_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout63_A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09749_ genblk2\[2\].wave_shpr.div.fin_quo\[7\] net1197 _00009_ VGND VGND VPWR VPWR
+ _04222_ sky130_fd_sc_hd__mux2_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10818__B1 _04858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12760_ clknet_leaf_93_clk _00001_ net146 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _05556_ _05601_ _05602_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__a21oi_2
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12691_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[4\] net174 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ net946 _05448_ _05445_ _05541_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11573_ net932 _05447_ _05484_ _05490_ VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13312_ clknet_leaf_118_clk _00633_ net138 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10524_ genblk2\[4\].wave_shpr.div.i\[1\] genblk2\[4\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _04756_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13243_ clknet_leaf_9_clk _00566_ net55 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10455_ _04598_ _04574_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__or2b_1
XFILLER_0_33_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13174_ clknet_leaf_129_clk _00499_ net65 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10386_ net602 _04657_ _04655_ genblk2\[4\].wave_shpr.div.quo\[10\] _04660_ VGND
+ VGND VPWR VPWR _00470_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12125_ genblk2\[10\].wave_shpr.div.acc\[12\] _05881_ _05865_ VGND VGND VPWR VPWR
+ _05882_ sky130_fd_sc_hd__mux2_1
XANTENNA__09492__A _01411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12056_ net440 _05823_ _05825_ net518 _05832_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11007_ _04990_ _04979_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__or2b_1
XFILLER_0_74_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12958_ clknet_leaf_136_clk _00287_ net42 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08478__B2 _02308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11909_ genblk2\[10\].wave_shpr.div.acc\[17\] genblk2\[10\].wave_shpr.div.b1\[17\]
+ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__or2b_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ clknet_leaf_30_clk _00220_ net96 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12358__A _03941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11262__A _04676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12026__A2 _05813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09089__D _03738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07100_ _01887_ _01906_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08080_ _01200_ _01680_ _02748_ _02749_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07031_ _01822_ _01849_ _01850_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__and3b_1
XFILLER_0_130_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13550__RESET_B net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08982_ _01097_ _03570_ _03666_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__or3_1
X_07933_ genblk2\[8\].wave_shpr.div.fin_quo\[3\] _02639_ VGND VGND VPWR VPWR _02640_
+ sky130_fd_sc_hd__or2_1
XANTENNA_fanout198_A net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07864_ _02517_ _02566_ _02570_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__a21o_1
XANTENNA__10341__A _03701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09603_ _03989_ _04103_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__xnor2_1
X_06815_ genblk1\[5\].osc.clkdiv_C.cnt\[12\] _01355_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07795_ genblk1\[0\].osc.clkdiv_C.cnt\[9\] _01184_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__nand2_1
Xwire20 _06088_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
Xwire31 _02508_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_2
X_09534_ net511 _04052_ _04053_ net519 _04057_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__a221o_1
X_06746_ _01627_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__inv_2
XANTENNA__09666__B1 _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10487__S _04704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09465_ _04020_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06677_ genblk1\[4\].osc.clkdiv_C.cnt\[5\] _01565_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08416_ _03114_ _03121_ _03122_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__o21ai_1
X_09396_ genblk2\[1\].wave_shpr.div.acc\[11\] genblk2\[1\].wave_shpr.div.b1\[11\]
+ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11225__B1 _05250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08347_ _03030_ _03051_ _03052_ _03053_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08278_ _02303_ _02264_ genblk2\[9\].wave_shpr.div.fin_quo\[4\] VGND VGND VPWR VPWR
+ _02985_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07229_ _01229_ _01230_ VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__nand2_4
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10240_ _04556_ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__clkbuf_1
X_10171_ _04394_ _04505_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout140 net145 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_4
Xfanout151 net152 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_4
Xfanout162 net163 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
Xfanout173 net174 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_4
Xfanout184 net185 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__buf_2
XANTENNA__10503__A2 _04715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout195 net198 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
X_12812_ clknet_leaf_58_clk net266 net192 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_70_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ clknet_leaf_49_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[2\] net108 VGND VGND
+ VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07132__B2 genblk1\[9\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_831 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12674_ clknet_leaf_90_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[5\] net174 VGND VGND
+ VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_154_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ genblk2\[8\].wave_shpr.div.acc\[18\] _05529_ VGND VGND VPWR VPWR _05530_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__06891__B1 _01484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11556_ _05449_ _05475_ _05477_ _05448_ net699 VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__a32o_1
XFILLER_0_13_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06904__A _01576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10507_ _04619_ _04622_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11487_ net713 VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10990__A2 _05023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13226_ clknet_leaf_127_clk net254 net132 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10438_ net842 _04683_ _04690_ _04693_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__a22o_1
XANTENNA__07199__A1 genblk1\[9\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08396__B1 _01209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13157_ clknet_leaf_121_clk _00482_ net78 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10369_ _04654_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ genblk2\[10\].wave_shpr.div.acc\[8\] _05868_ _05865_ VGND VGND VPWR VPWR
+ _05869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ clknet_leaf_137_clk _00415_ net40 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08148__B1 _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12039_ _05812_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_06600_ _01241_ _01432_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__nor2_2
X_07580_ _01432_ _01221_ genblk1\[9\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _02287_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06531_ genblk1\[2\].osc.clkdiv_C.cnt\[1\] genblk1\[2\].osc.clkdiv_C.cnt\[0\] genblk1\[2\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09250_ _03853_ genblk1\[0\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06462_ genblk1\[1\].osc.clkdiv_C.cnt\[10\] _01394_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__nand2_1
X_08201_ net17 _02552_ genblk2\[10\].wave_shpr.div.fin_quo\[6\] VGND VGND VPWR VPWR
+ _02908_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06882__B1 _01735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09181_ _03817_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__clkbuf_1
X_06393_ _01336_ _01226_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__nor2_4
XFILLER_0_29_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08132_ genblk2\[4\].wave_shpr.div.fin_quo\[0\] genblk2\[4\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08063_ genblk1\[5\].osc.clkdiv_C.cnt\[2\] _01238_ net35 VGND VGND VPWR VPWR _02770_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_43_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07014_ genblk1\[7\].osc.clkdiv_C.cnt\[10\] _01837_ _01839_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[10\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08965_ _03650_ _03652_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__xnor2_1
X_07916_ genblk1\[8\].osc.clkdiv_C.cnt\[4\] _01487_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__or2_1
X_08896_ sig_norm.b1\[0\] _03578_ _03580_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__nand3_1
X_07847_ _02217_ _02553_ genblk2\[0\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR
+ _02554_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07778_ _01181_ genblk1\[0\].osc.clkdiv_C.cnt\[7\] _01198_ VGND VGND VPWR VPWR _02485_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__11446__A0 genblk2\[8\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09517_ genblk2\[1\].wave_shpr.div.quo\[7\] _04043_ _04047_ net292 VGND VGND VPWR
+ VPWR _00214_ sky130_fd_sc_hd__a22o_1
X_06729_ _01600_ _01613_ _01614_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__and3_1
XANTENNA__13532__D _00023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11997__A1 _01556_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09448_ genblk2\[1\].wave_shpr.div.fin_quo\[0\] _04011_ _00007_ VGND VGND VPWR VPWR
+ _04012_ sky130_fd_sc_hd__mux2_1
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09379_ _03942_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11410_ genblk2\[8\].wave_shpr.div.b1\[6\] genblk2\[8\].wave_shpr.div.acc\[6\] VGND
+ VGND VPWR VPWR _05386_ sky130_fd_sc_hd__and2b_1
X_12390_ genblk2\[11\].wave_shpr.div.acc\[10\] _06064_ _06055_ VGND VGND VPWR VPWR
+ _06065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11341_ net628 _05311_ _05315_ _05330_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11272_ genblk2\[7\].wave_shpr.div.acc\[1\] _05277_ _05222_ VGND VGND VPWR VPWR _05278_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13011_ clknet_leaf_133_clk _00340_ net59 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10223_ net524 _04518_ _04522_ _04545_ VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__a22o_1
XANTENNA__09754__B _01925_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10154_ net979 _04486_ _04490_ _04493_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10085_ net794 _04452_ _04420_ _04454_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__a22o_1
Xhold7 modein.delay_octave_down_in\[0\] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11524__B genblk1\[8\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10987_ _05054_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__inv_2
XANTENNA__11988__A1 _01946_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12726_ clknet_leaf_37_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[3\] net113 VGND VGND
+ VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_128_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12657_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[6\] net90 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_154_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11608_ _05402_ _05361_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__or2b_1
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08066__C1 genblk1\[5\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09802__B1 _04252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12588_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[9\] net72 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_80_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07449__B _02153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11539_ _05464_ genblk1\[8\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold407 genblk2\[5\].wave_shpr.div.b1\[5\] VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 genblk2\[0\].wave_shpr.div.quo\[20\] VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold429 _00913_ VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13209_ clknet_leaf_25_clk _00532_ net86 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06395__A2 _01210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _03455_ _03456_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__or2_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 genblk2\[8\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net1325 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 genblk2\[5\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net1336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 genblk2\[7\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net1347 sky130_fd_sc_hd__dlygate4sd3_1
X_07701_ genblk2\[10\].wave_shpr.div.fin_quo\[2\] _02407_ VGND VGND VPWR VPWR _02408_
+ sky130_fd_sc_hd__and2b_1
X_08681_ _03113_ _03115_ genblk2\[2\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR
+ _03388_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08541__B1 _02308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07632_ genblk1\[11\].osc.clkdiv_C.cnt\[10\] _01262_ _02338_ VGND VGND VPWR VPWR
+ _02339_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_136_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07563_ _01930_ _01556_ _01564_ _01801_ _01928_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__a32o_1
XANTENNA__07631__C _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09302_ genblk2\[0\].wave_shpr.div.acc\[7\] _03888_ _03889_ VGND VGND VPWR VPWR _03890_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06514_ _01191_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07494_ net17 VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__buf_2
XANTENNA__10100__B1 _04454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09233_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06445_ _01384_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09164_ _03808_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06376_ freq_div.state\[0\] _01178_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_127_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08115_ _01172_ _01180_ _01568_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06607__B1 _01514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08072__A2 _01309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09095_ _01211_ _01556_ _03743_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09855__A _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08046_ genblk1\[5\].osc.clkdiv_C.cnt\[13\] _01674_ _01666_ genblk1\[5\].osc.clkdiv_C.cnt\[12\]
+ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold930 genblk2\[3\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR net1148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold941 genblk1\[2\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR net1159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 sig_norm.quo\[4\] VGND VGND VPWR VPWR net1170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold963 genblk2\[7\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR net1181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 genblk2\[4\].wave_shpr.div.b1\[11\] VGND VGND VPWR VPWR net1192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 genblk2\[11\].wave_shpr.div.acc\[20\] VGND VGND VPWR VPWR net1203 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11903__A1 _03839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold996 genblk2\[8\].wave_shpr.div.b1\[3\] VGND VGND VPWR VPWR net1214 sky130_fd_sc_hd__dlygate4sd3_1
X_09997_ genblk2\[3\].wave_shpr.div.b1\[7\] genblk2\[3\].wave_shpr.div.acc\[7\] VGND
+ VGND VPWR VPWR _04393_ sky130_fd_sc_hd__and2b_1
XANTENNA__07583__A1 genblk1\[9\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08948_ _01098_ _03559_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__or2_1
X_08879_ _03575_ sig_norm.acc\[3\] _03584_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__o21a_1
XANTENNA__08532__B1 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10910_ _05039_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07822__B net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07886__A2 _02539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11890_ genblk2\[9\].wave_shpr.div.acc\[24\] _05646_ _05715_ VGND VGND VPWR VPWR
+ _05719_ sky130_fd_sc_hd__or3b_1
X_10841_ _04982_ _04983_ _04984_ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__o21ai_1
X_13560_ clknet_leaf_84_clk net291 net184 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10772_ net925 _04918_ _04922_ _04931_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12511_ clknet_leaf_84_clk _00073_ net202 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10642__A1 _04645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13491_ clknet_leaf_88_clk _00808_ net177 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12442_ genblk2\[11\].wave_shpr.div.acc\[24\] _05980_ genblk2\[11\].wave_shpr.div.acc\[25\]
+ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12373_ genblk2\[11\].wave_shpr.div.acc\[6\] _06051_ _05982_ VGND VGND VPWR VPWR
+ _06052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10945__A2 _05052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11324_ genblk2\[7\].wave_shpr.div.acc\[13\] _05317_ _05300_ VGND VGND VPWR VPWR
+ _05318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11255_ genblk2\[7\].wave_shpr.div.quo\[21\] _05255_ _05256_ net527 _05267_ VGND
+ VGND VPWR VPWR _00732_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10206_ _04532_ _04410_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11519__B genblk1\[8\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11186_ genblk2\[8\].wave_shpr.div.b1\[5\] _01508_ _05042_ VGND VGND VPWR VPWR _05233_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07574__A1 _01336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10137_ _04417_ _04418_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__nor2_2
X_10068_ _01325_ _01226_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__nor2_2
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12130__S _05865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13758_ clknet_leaf_66_clk _01069_ net197 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12083__B1 _05817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13394__RESET_B net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12709_ clknet_leaf_56_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[4\] net181 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
X_13689_ clknet_leaf_57_clk _00004_ net184 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06230_ _01175_ _01191_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__nand2_4
XFILLER_0_127_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06161_ _01130_ _01132_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold204 _00719_ VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold215 _00958_ VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__A2 _01577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold226 _01045_ VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold237 _00147_ VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09920_ genblk2\[2\].wave_shpr.div.acc\[16\] _04330_ _04301_ VGND VGND VPWR VPWR
+ _04331_ sky130_fd_sc_hd__mux2_1
Xhold248 genblk2\[0\].wave_shpr.div.quo\[18\] VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold259 genblk2\[6\].wave_shpr.div.quo\[9\] VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10149__B1 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06811__B _01326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09851_ genblk2\[2\].wave_shpr.div.b1\[0\] genblk2\[2\].wave_shpr.div.acc\[0\] _04214_
+ _04275_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__a31o_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _03219_ _03222_ _03220_ _03221_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__o211a_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11361__A2 _05248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06672__A2_N _01326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _03702_ _01490_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__nand2_4
X_06994_ genblk1\[7\].osc.clkdiv_C.cnt\[3\] _01825_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__and2_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _03175_ _03201_ _03200_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout180_A net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ _02798_ _03370_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ genblk1\[11\].osc.clkdiv_C.cnt\[2\] _01186_ _01437_ _01225_ VGND VGND VPWR
+ VPWR _02322_ sky130_fd_sc_hd__or4_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _02798_ _03299_ _03301_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07546_ _02256_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09490__A1 _04034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07477_ _02201_ _02153_ genblk2\[9\].wave_shpr.div.busy VGND VGND VPWR VPWR _02204_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11180__A _03708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09216_ _03837_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06428_ genblk1\[1\].osc.clkdiv_C.cnt\[0\] _01304_ _01319_ _01331_ _01371_ VGND VGND
+ VPWR VPWR _01372_ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09147_ genblk2\[0\].wave_shpr.div.b1\[16\] genblk2\[0\].wave_shpr.div.acc\[16\]
+ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08045__A2 _01675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06359_ _01179_ _01222_ _01302_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09078_ _03702_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__buf_8
XFILLER_0_102_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08029_ genblk2\[6\].wave_shpr.div.fin_quo\[2\] _02735_ VGND VGND VPWR VPWR _02736_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07817__B net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold760 genblk2\[8\].wave_shpr.div.acc\[8\] VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 genblk2\[10\].wave_shpr.div.acc\[2\] VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 genblk2\[3\].wave_shpr.div.acc\[23\] VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ _05051_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__clkbuf_4
Xhold793 _00753_ VGND VGND VPWR VPWR net1011 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11888__B1 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12991_ clknet_leaf_130_clk _00320_ net65 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08505__B1 _02224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11942_ genblk2\[10\].wave_shpr.div.b1\[9\] genblk2\[10\].wave_shpr.div.acc\[9\]
+ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11873_ genblk2\[9\].wave_shpr.div.acc\[19\] _05704_ VGND VGND VPWR VPWR _05707_
+ sky130_fd_sc_hd__or2_1
X_13612_ clknet_leaf_94_clk _00925_ net159 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10824_ genblk2\[6\].wave_shpr.div.acc\[15\] genblk2\[6\].wave_shpr.div.b1\[15\]
+ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__or2b_1
XANTENNA__12065__B1 _05815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10615__A1 _01684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13543_ clknet_leaf_101_clk _00858_ net164 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10755_ _02183_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06295__A1 _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10091__A2 _04452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13474_ clknet_leaf_71_clk _00791_ net215 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10686_ net235 _04861_ _04862_ net378 _04870_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12425_ net641 _06072_ _06073_ _06091_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08036__A2 _02539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12356_ net1020 _06009_ _06010_ _06038_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__a22o_1
X_11307_ net797 _05279_ _05283_ _05304_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12125__S _05865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10434__A _04654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12287_ _01337_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__inv_2
X_11238_ net640 _05255_ _05256_ net670 _05258_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__a221o_1
X_11169_ genblk2\[7\].wave_shpr.div.fin_quo\[3\] genblk2\[7\].wave_shpr.div.quo\[2\]
+ _00019_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06359__A _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07400_ net1220 _02145_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08380_ genblk1\[2\].osc.clkdiv_C.cnt\[1\] _01209_ _02425_ genblk1\[2\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07331_ genblk1\[11\].osc.clkdiv_C.cnt\[1\] genblk1\[11\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _02094_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08275__A2 _02361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06806__B _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07262_ genblk1\[10\].osc.clkdiv_C.cnt\[5\] genblk1\[10\].osc.clkdiv_C.cnt\[4\] _02034_
+ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09001_ _03680_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06213_ freq_div.state\[1\] VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__buf_4
X_07193_ net1296 _01978_ _01980_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06144_ _01113_ _01115_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__nand2_1
XANTENNA__07918__A _01489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10344__A _01678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09903_ genblk2\[2\].wave_shpr.div.acc\[12\] _04317_ _04301_ VGND VGND VPWR VPWR
+ _04318_ sky130_fd_sc_hd__mux2_1
Xwire5 _02589_ VGND VGND VPWR VPWR net1354 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09834_ genblk2\[2\].wave_shpr.div.quo\[20\] _04257_ _04259_ net322 _04267_ VGND
+ VGND VPWR VPWR _00311_ sky130_fd_sc_hd__a221o_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _04232_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__clkbuf_1
X_06977_ genblk1\[7\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__inv_2
X_08716_ _03387_ _03391_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__or2b_1
XANTENNA__11098__A1 _05055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09696_ _04174_ _04175_ _04172_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__o21ai_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06269__A _01229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08647_ _03289_ _03290_ _02419_ _03284_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08578_ genblk2\[10\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__inv_2
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07529_ _01099_ _02245_ _02246_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10540_ genblk2\[5\].wave_shpr.div.acc\[12\] genblk2\[5\].wave_shpr.div.b1\[12\]
+ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__or2b_1
XFILLER_0_119_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10471_ net778 _04715_ _04690_ _04718_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12210_ _05939_ _05946_ _05947_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13190_ clknet_leaf_118_clk _00513_ net138 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12141_ _05893_ _05777_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09518__A2 _04043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12072_ genblk2\[10\].wave_shpr.div.acc\[0\] _00002_ _05840_ net247 _05841_ VGND
+ VGND VPWR VPWR _00975_ sky130_fd_sc_hd__o221a_1
Xhold590 genblk2\[7\].wave_shpr.div.acc\[13\] VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__dlygate4sd3_1
X_11023_ net867 _05086_ _05093_ _05106_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__a22o_1
XANTENNA__10533__B1 _03855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12974_ clknet_leaf_124_clk net554 net71 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11925_ genblk2\[10\].wave_shpr.div.acc\[0\] genblk2\[10\].wave_shpr.div.b1\[0\]
+ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__or2b_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12038__B1 _05816_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06517__A2_N _01439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11856_ net912 _05684_ _05685_ _05694_ VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__a22o_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10807_ _04856_ _02183_ genblk2\[5\].wave_shpr.div.i\[0\] VGND VGND VPWR VPWR _04956_
+ sky130_fd_sc_hd__mux2_1
X_11787_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10738_ _04796_ _04772_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__or2b_1
X_13526_ clknet_leaf_98_clk _00843_ net169 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13457_ clknet_leaf_99_clk _00774_ net165 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_10669_ genblk2\[5\].wave_shpr.div.quo\[10\] _04858_ _04855_ net310 _04860_ VGND
+ VGND VPWR VPWR _00553_ sky130_fd_sc_hd__a221o_1
XANTENNA__11549__C1 _05472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08841__B _03544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12408_ genblk2\[11\].wave_shpr.div.acc\[14\] _06078_ _06055_ VGND VGND VPWR VPWR
+ _06079_ sky130_fd_sc_hd__mux2_1
X_13388_ clknet_leaf_78_clk _00707_ net208 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12339_ net434 _03942_ _03941_ net438 _06027_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__a221o_1
XANTENNA__06361__B _01226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06900_ _01753_ genblk1\[6\].osc.clkdiv_C.cnt\[0\] _01363_ genblk1\[6\].osc.clkdiv_C.cnt\[15\]
+ genblk1\[6\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__a221o_1
X_07880_ _02424_ _02471_ _02519_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__o21a_1
X_06831_ genblk1\[5\].osc.clkdiv_C.cnt\[3\] _01698_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__and2_1
X_09550_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__and2_1
X_06762_ genblk1\[4\].osc.clkdiv_C.cnt\[12\] _01637_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__or2_1
X_08501_ net24 _03207_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__or2b_1
X_09481_ _04029_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06693_ genblk1\[4\].osc.clkdiv_C.cnt\[11\] _01313_ _01340_ genblk1\[4\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08432_ _03137_ _03138_ genblk2\[9\].wave_shpr.div.fin_quo\[3\] _02308_ VGND VGND
+ VPWR VPWR _03139_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12029__B1 _05817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08363_ _02939_ _03069_ _02943_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout143_A net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07314_ genblk1\[11\].osc.clkdiv_C.cnt\[12\] _02077_ genblk1\[11\].osc.clkdiv_C.cnt\[17\]
+ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08294_ _02998_ _02999_ _03000_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__nor3_1
XFILLER_0_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12638__RESET_B net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07245_ _02026_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08751__B _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07176_ genblk1\[9\].osc.clkdiv_C.cnt\[7\] _01967_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06127_ _01098_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__buf_2
XFILLER_0_2_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11307__A2 _05279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09074__S _03722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09817_ net553 _04257_ _04251_ genblk2\[2\].wave_shpr.div.quo\[11\] _04258_ VGND
+ VGND VPWR VPWR _00303_ sky130_fd_sc_hd__a221o_1
X_09748_ _04221_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout56_A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10818__A1 _04855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ genblk2\[2\].wave_shpr.div.acc\[14\] genblk2\[2\].wave_shpr.div.b1\[14\]
+ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__or2b_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ genblk2\[9\].wave_shpr.div.b1\[15\] genblk2\[9\].wave_shpr.div.acc\[15\]
+ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__and2b_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ clknet_leaf_53_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[3\] net174 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_hold522_A genblk2\[10\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11641_ genblk2\[8\].wave_shpr.div.acc\[23\] _05412_ _05540_ VGND VGND VPWR VPWR
+ _05541_ sky130_fd_sc_hd__a21o_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11572_ genblk2\[8\].wave_shpr.div.acc\[5\] _05489_ _05417_ VGND VGND VPWR VPWR _05490_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13311_ clknet_leaf_118_clk net721 net137 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10523_ genblk2\[4\].wave_shpr.div.i\[1\] genblk2\[4\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _04755_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13242_ clknet_leaf_9_clk net246 net55 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10454_ net891 _04683_ _04690_ _04705_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__a22o_1
XANTENNA__06462__A genblk1\[1\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11546__A2 _05441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13173_ clknet_leaf_128_clk _00498_ net66 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10385_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__and2_1
X_12124_ _05769_ _05880_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06973__A2 _01363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12055_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR _05832_
+ sky130_fd_sc_hd__and2_1
X_11006_ _05054_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12957_ clknet_leaf_114_clk _00286_ net132 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11482__A1 _02656_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11908_ net273 _05729_ _05730_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__a21oi_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12888_ clknet_leaf_30_clk _00219_ net96 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07150__A2 _01799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09013__A _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11839_ _05594_ _05560_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__or2b_1
XFILLER_0_145_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13509_ clknet_leaf_80_clk _00826_ net205 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07030_ genblk1\[7\].osc.clkdiv_C.cnt\[16\] _01847_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__nand2_1
XANTENNA__07468__A _02147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08402__A2 _01411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08981_ _03525_ _03568_ _03569_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__and3_1
X_07932_ genblk2\[8\].wave_shpr.div.fin_quo\[0\] genblk2\[8\].wave_shpr.div.fin_quo\[1\]
+ genblk2\[8\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__or3_1
X_07863_ _02469_ _02569_ _02529_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__o21a_1
XANTENNA__07913__A1 genblk1\[8\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09602_ _03990_ _03961_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__or2b_1
X_06814_ genblk1\[5\].osc.clkdiv_C.cnt\[6\] _01242_ _01682_ _01683_ _01685_ VGND VGND
+ VPWR VPWR _01686_ sky130_fd_sc_hd__a221o_1
X_07794_ _02478_ _02492_ _02495_ _02500_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__or4b_1
XANTENNA__09622__S _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07931__A net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09533_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06745_ genblk1\[4\].osc.clkdiv_C.cnt\[8\] genblk1\[4\].osc.clkdiv_C.cnt\[7\] _01620_
+ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__and3_1
Xwire32 _02302_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09666__A1 _04045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09464_ genblk2\[2\].wave_shpr.div.b1\[0\] net35 _03822_ VGND VGND VPWR VPWR _04020_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11473__A1 _04230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06676_ genblk1\[4\].osc.clkdiv_C.cnt\[5\] _01565_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__and2_1
X_08415_ net8 _02744_ _02365_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__and3_2
XFILLER_0_65_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09395_ genblk2\[1\].wave_shpr.div.acc\[12\] genblk2\[1\].wave_shpr.div.b1\[12\]
+ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__or2b_1
XFILLER_0_80_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08346_ _02993_ _02994_ _02995_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08277_ _02977_ _02983_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__and2b_1
XFILLER_0_117_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10984__B1 _05054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07228_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _01235_ _01227_ genblk1\[10\].osc.clkdiv_C.cnt\[9\]
+ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_132_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07159_ _01957_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[1\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__07062__D1 genblk1\[8\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10170_ _04395_ _04370_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__or2b_1
Xfanout130 net131 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10532__A _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout141 net145 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout152 net158 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_4
Xfanout163 net171 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
Xfanout174 net218 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__buf_2
Xfanout185 net218 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13260__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06707__A2 _01304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout196 net198 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_4
X_12811_ clknet_leaf_59_clk _00144_ net192 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11464__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07668__B1 _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ clknet_leaf_50_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[1\] net108 VGND VGND
+ VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ clknet_leaf_90_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[4\] net173 VGND VGND
+ VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11624_ _05409_ _05416_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_92_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11555_ _05417_ _05476_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__nand2_1
XANTENNA__08391__B _01302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06904__B _01757_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10506_ genblk2\[4\].wave_shpr.div.acc\[20\] _04740_ VGND VGND VPWR VPWR _04744_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_52_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11486_ _03831_ net390 _03717_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_80_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13225_ clknet_leaf_114_clk _00548_ net133 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10437_ genblk2\[4\].wave_shpr.div.acc\[3\] _04692_ _04623_ VGND VGND VPWR VPWR _04693_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13156_ clknet_leaf_121_clk net666 net78 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _04653_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__clkbuf_4
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12107_ _05761_ _05867_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__xnor2_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ clknet_leaf_136_clk _00414_ net42 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ _04568_ _04609_ _04610_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__a21o_1
X_12038_ net223 _05818_ _05816_ net398 _05822_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06530_ genblk1\[2\].osc.clkdiv_C.cnt\[2\] genblk1\[2\].osc.clkdiv_C.cnt\[1\] genblk1\[2\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__and3_1
XANTENNA__07470__B _02153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12912__RESET_B net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08320__B2 _02362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06461_ _01373_ _01394_ _01395_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_146_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08200_ _02405_ _02403_ _02410_ _02524_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__o31a_1
XFILLER_0_145_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09180_ net1249 _01356_ _03722_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06392_ _01179_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08131_ _02221_ _02837_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__nor2_2
XFILLER_0_50_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10617__A _03701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08062_ _02766_ _02768_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__nand2_1
XANTENNA__07831__B1 _02224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07013_ genblk1\[7\].osc.clkdiv_C.cnt\[10\] _01837_ _01822_ VGND VGND VPWR VPWR _01839_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout106_A net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07595__C1 genblk1\[9\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08964_ _03651_ _03646_ _03506_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__a21oi_1
X_07915_ genblk1\[8\].osc.clkdiv_C.cnt\[3\] _01866_ _01487_ genblk1\[8\].osc.clkdiv_C.cnt\[4\]
+ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__a22o_1
X_08895_ net629 _03596_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__or2_1
X_07846_ _02552_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__clkbuf_2
XANTENNA__07898__B1 _01576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07777_ genblk1\[0\].osc.clkdiv_C.cnt\[4\] _01258_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09516_ net292 _04043_ _04047_ net771 VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__a22o_1
X_06728_ genblk1\[4\].osc.clkdiv_C.cnt\[4\] _01609_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09447_ _04010_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06659_ _01522_ _01551_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__nor2_1
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09378_ genblk2\[11\].wave_shpr.div.i\[1\] genblk2\[11\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _03946_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11749__A2 _05623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08329_ genblk2\[7\].wave_shpr.div.fin_quo\[4\] VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08075__B1 _01726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11340_ genblk2\[7\].wave_shpr.div.acc\[17\] _05329_ _05300_ VGND VGND VPWR VPWR
+ _05330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11271_ _05184_ _05276_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__nor2_1
X_13010_ clknet_leaf_133_clk _00339_ net59 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10222_ _04543_ _04544_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10153_ genblk2\[3\].wave_shpr.div.acc\[3\] _04492_ _04420_ VGND VGND VPWR VPWR _04493_
+ sky130_fd_sc_hd__mux2_1
X_10084_ _04453_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__buf_4
Xhold8 genblk2\[9\].wave_shpr.div.quo\[22\] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10488__A2 _04715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07571__A genblk1\[9\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06187__A _01157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10986_ net283 _05051_ _05054_ net668 _05078_ VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__a221o_1
X_13774_ clknet_leaf_73_clk _01085_ net213 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12725_ clknet_leaf_37_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[2\] net113 VGND VGND
+ VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10660__A2 _04853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12656_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[5\] net90 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08066__B1 _01171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11607_ net846 _05507_ _05484_ _05516_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12587_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[8\] net72 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11538_ net575 _05454_ _05458_ net660 _05466_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold408 genblk2\[4\].wave_shpr.div.quo\[20\] VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 genblk2\[4\].wave_shpr.div.quo\[13\] VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ _05431_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09566__B1 _04047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13208_ clknet_leaf_8_clk _00531_ net88 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13139_ clknet_leaf_115_clk net750 net133 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 genblk2\[5\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net1326 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1119 genblk2\[8\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net1337 sky130_fd_sc_hd__dlygate4sd3_1
X_07700_ genblk2\[10\].wave_shpr.div.fin_quo\[0\] genblk2\[10\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__nor2_1
X_08680_ _03307_ _03330_ _03328_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08541__A1 genblk2\[8\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08541__B2 genblk2\[8\].wave_shpr.div.fin_quo\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07631_ _02128_ _01179_ _01249_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07562_ genblk1\[9\].osc.clkdiv_C.cnt\[11\] _01799_ _01731_ _02268_ VGND VGND VPWR
+ VPWR _02269_ sky130_fd_sc_hd__a2bb2o_1
X_09301_ _03803_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__buf_4
XFILLER_0_75_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06513_ _01213_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__buf_4
XFILLER_0_152_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07493_ modein.delay_in\[0\] VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09232_ net569 _03841_ _03839_ net598 _03843_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06444_ _01374_ _01382_ _01383_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10545__B_N genblk2\[5\].wave_shpr.div.b1\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09163_ genblk2\[0\].wave_shpr.div.fin_quo\[3\] net1314 _00001_ VGND VGND VPWR VPWR
+ _03808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06375_ _01306_ _01315_ _01316_ _01318_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__or4b_1
X_08114_ _02811_ _02820_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__nand2_1
X_09094_ _01367_ _03739_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08072__A3 _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08045_ genblk1\[5\].osc.clkdiv_C.cnt\[13\] _01675_ _02748_ _02751_ VGND VGND VPWR
+ VPWR _02752_ sky130_fd_sc_hd__a211o_1
Xhold920 genblk2\[6\].wave_shpr.div.acc\[20\] VGND VGND VPWR VPWR net1138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold931 genblk2\[9\].wave_shpr.div.i\[2\] VGND VGND VPWR VPWR net1149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 genblk2\[4\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR net1160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 genblk2\[10\].wave_shpr.div.b1\[2\] VGND VGND VPWR VPWR net1171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 genblk1\[8\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR net1182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold975 genblk1\[3\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR net1193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 genblk2\[11\].wave_shpr.div.b1\[10\] VGND VGND VPWR VPWR net1204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 genblk2\[7\].wave_shpr.div.fin_quo\[7\] VGND VGND VPWR VPWR net1215 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10082__A _04451_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09996_ _04372_ _04390_ _04391_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07583__A2 _01234_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08947_ _03557_ _03558_ _03546_ _03551_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11906__A _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08878_ _03576_ sig_norm.acc\[2\] _03583_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07829_ _02530_ _02535_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__nor2_1
X_10840_ genblk2\[6\].wave_shpr.div.b1\[1\] genblk2\[6\].wave_shpr.div.acc\[1\] VGND
+ VGND VPWR VPWR _04984_ sky130_fd_sc_hd__or2b_1
XFILLER_0_67_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_99_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10771_ genblk2\[5\].wave_shpr.div.acc\[15\] _04930_ _04907_ VGND VGND VPWR VPWR
+ _04931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12510_ clknet_leaf_84_clk net1040 net202 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_136_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13490_ clknet_leaf_88_clk _00807_ net177 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12441_ net1078 _03947_ _03944_ _06101_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12372_ _05952_ _06050_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11323_ _05206_ _05316_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11254_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06470__A genblk1\[1\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07559__C1 genblk1\[9\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10205_ _04411_ _04362_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11185_ _03727_ _01432_ net593 _03687_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07574__A2 _01437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10136_ _03819_ net436 _00010_ genblk2\[3\].wave_shpr.div.acc\[0\] _04479_ VGND VGND
+ VPWR VPWR _00401_ sky130_fd_sc_hd__o221a_1
X_10067_ _04443_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11535__B genblk1\[8\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13757_ clknet_leaf_70_clk _01068_ net213 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_136_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_136_clk sky130_fd_sc_hd__clkbuf_16
X_10969_ net582 _05062_ _05064_ net595 _05069_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__a221o_1
XANTENNA__10094__B1 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12708_ clknet_leaf_56_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[3\] net181 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13688_ clknet_leaf_63_clk _01001_ net190 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12639_ clknet_leaf_16_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[6\] net73 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06160_ _01117_ _01131_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold205 genblk2\[5\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 genblk2\[11\].wave_shpr.div.quo\[23\] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 genblk2\[8\].wave_shpr.div.quo\[24\] VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 genblk2\[8\].wave_shpr.div.acc\[22\] VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07476__A _02203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold249 genblk2\[11\].wave_shpr.div.quo\[10\] VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09850_ genblk2\[2\].wave_shpr.div.b1\[0\] _04214_ genblk2\[2\].wave_shpr.div.acc\[0\]
+ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__a21oi_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07565__A2 _01328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08801_ _03451_ _03506_ _03507_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__o21bai_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _04240_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__clkbuf_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06993_ _01823_ _01825_ _01826_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _03431_ _03438_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__xnor2_1
X_08663_ genblk2\[5\].wave_shpr.div.fin_quo\[3\] _02521_ _02791_ _03369_ VGND VGND
+ VPWR VPWR _03370_ sky130_fd_sc_hd__a211o_1
XANTENNA__07722__C1 _01172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07614_ _01171_ _01192_ _01208_ genblk1\[11\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR
+ VPWR _02321_ sky130_fd_sc_hd__a31o_1
X_08594_ net10 _02364_ _03300_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__and3_1
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09630__S _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07545_ PWM.final_sample_in\[4\] net1150 PWM.start VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_127_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_127_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__10085__B1 _04420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07476_ _02203_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11180__B genblk2\[8\].wave_shpr.div.b1\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06427_ _01335_ _01353_ _01357_ _01370_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__or4b_1
X_09215_ _02152_ genblk2\[0\].wave_shpr.div.busy _02149_ VGND VGND VPWR VPWR _03837_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_17_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09146_ _03748_ _03792_ _03793_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__a21o_1
XANTENNA__09866__A _04250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09501__B1_N _03717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06358_ _01301_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__buf_6
XFILLER_0_16_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09077_ _03731_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__clkbuf_1
X_06289_ _01246_ _01250_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08028_ genblk2\[6\].wave_shpr.div.fin_quo\[0\] genblk2\[6\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold750 genblk2\[2\].wave_shpr.div.acc\[22\] VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 genblk2\[3\].wave_shpr.div.acc\[4\] VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 genblk2\[1\].wave_shpr.div.acc\[2\] VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 genblk2\[6\].wave_shpr.div.acc\[21\] VGND VGND VPWR VPWR net1001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold794 genblk2\[5\].wave_shpr.div.acc\[23\] VGND VGND VPWR VPWR net1012 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11888__A1 _03694_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout86_A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09950__B1 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09979_ genblk2\[3\].wave_shpr.div.acc\[4\] genblk2\[3\].wave_shpr.div.b1\[4\] VGND
+ VGND VPWR VPWR _04375_ sky130_fd_sc_hd__or2b_1
X_12990_ clknet_leaf_131_clk _00319_ net65 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07308__A2 _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12301__A2 _06009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11941_ _05740_ _05761_ _05762_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11872_ net1023 _05684_ _05685_ _05706_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__a22o_1
X_13611_ clknet_leaf_93_clk _00924_ net159 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10823_ genblk2\[6\].wave_shpr.div.b1\[16\] genblk2\[6\].wave_shpr.div.acc\[16\]
+ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_118_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_118_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13542_ clknet_leaf_101_clk _00857_ net165 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10754_ net1014 _04886_ _04890_ _04917_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__a22o_1
XANTENNA__06465__A genblk1\[1\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10685_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__and2_1
X_13473_ clknet_leaf_74_clk _00790_ net215 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06184__B _01095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12424_ _06089_ _06090_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08441__B1 _02361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12355_ genblk2\[11\].wave_shpr.div.acc\[2\] _06037_ _05982_ VGND VGND VPWR VPWR
+ _06038_ sky130_fd_sc_hd__mux2_1
X_11306_ genblk2\[7\].wave_shpr.div.acc\[9\] _05303_ _05300_ VGND VGND VPWR VPWR _05304_
+ sky130_fd_sc_hd__mux2_1
X_12286_ _03726_ _01312_ _06004_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__a21oi_1
X_11237_ _05074_ genblk1\[7\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__and2_1
X_11168_ _05225_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__clkbuf_1
X_10119_ net451 _04461_ _04462_ genblk2\[3\].wave_shpr.div.quo\[17\] _04470_ VGND
+ VGND VPWR VPWR _00393_ sky130_fd_sc_hd__a221o_1
X_11099_ _00016_ _05159_ net1177 VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09016__A _02155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11500__B1 _05446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09450__S _00007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10596__S _00015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_109_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_109_clk sky130_fd_sc_hd__clkbuf_16
X_07330_ _02093_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07261_ _02038_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09000_ net1102 net1126 _01154_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06212_ _01173_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_143_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07192_ _01953_ _01979_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__nor2_1
XANTENNA__09224__A2 _03836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06143_ net14 _01112_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07918__B genblk1\[8\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09902_ _04196_ _04316_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09833_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__and2_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ net1245 _01794_ _04039_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__mux2_1
X_06976_ genblk1\[7\].osc.clkdiv_C.cnt\[12\] _01811_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__xnor2_1
X_08715_ _03383_ _03395_ _03420_ _03421_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__a211o_1
XANTENNA__12295__A1 _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09695_ genblk2\[2\].wave_shpr.div.acc\[0\] genblk2\[2\].wave_shpr.div.b1\[0\] VGND
+ VGND VPWR VPWR _04175_ sky130_fd_sc_hd__and2b_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _03140_ _03150_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__xor2_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07171__B1 genblk1\[9\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07710__A2 _02362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08577_ _03141_ _03283_ _02901_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__o21a_1
XANTENNA__12287__A _01337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07528_ sig_norm.busy sig_norm.i\[0\] sig_norm.i\[1\] VGND VGND VPWR VPWR _02246_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07459_ _02190_ genblk2\[7\].wave_shpr.div.i\[1\] genblk2\[7\].wave_shpr.div.i\[0\]
+ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__or3b_1
X_10470_ genblk2\[4\].wave_shpr.div.acc\[11\] _04717_ _04704_ VGND VGND VPWR VPWR
+ _04718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09129_ genblk2\[0\].wave_shpr.div.b1\[7\] genblk2\[0\].wave_shpr.div.acc\[7\] VGND
+ VGND VPWR VPWR _03777_ sky130_fd_sc_hd__and2b_1
X_12140_ _05778_ _05732_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12071_ _03719_ genblk1\[10\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR _05841_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold580 _00747_ VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 genblk2\[7\].wave_shpr.div.acc\[15\] VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ genblk2\[6\].wave_shpr.div.acc\[7\] _05104_ _05105_ VGND VGND VPWR VPWR _05106_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_hold934_A genblk2\[3\].wave_shpr.div.b1\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11089__A2 _05057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12286__A1 _03726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12973_ clknet_leaf_124_clk net442 net71 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11924_ genblk2\[10\].wave_shpr.div.acc\[1\] genblk2\[10\].wave_shpr.div.b1\[1\]
+ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__xnor2_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ genblk2\[9\].wave_shpr.div.acc\[14\] _05693_ _05673_ VGND VGND VPWR VPWR
+ _05694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08394__B _01411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10806_ net392 _04858_ _04855_ _04955_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11786_ genblk2\[9\].wave_shpr.div.quo\[23\] _02203_ _03693_ net226 _05642_ VGND
+ VGND VPWR VPWR _00888_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13525_ clknet_leaf_98_clk _00842_ net169 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10737_ net927 _04886_ _04890_ _04904_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__a22o_1
XANTENNA__11261__A2 _05245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13456_ clknet_leaf_100_clk _00773_ net164 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_36_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10668_ _04672_ genblk1\[5\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12407_ _05968_ _06077_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07738__B _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07217__B2 _01342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10599_ _04824_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__clkbuf_1
X_13387_ clknet_leaf_83_clk _00706_ net200 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12338_ _03833_ _02081_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12269_ _05995_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__clkbuf_1
X_06830_ _01693_ _01698_ _01699_ VGND VGND VPWR VPWR genblk1\[5\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
X_06761_ _01639_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[11\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__12277__A1 _02001_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08500_ _02520_ _02587_ _03206_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__o21ai_1
X_09480_ genblk2\[2\].wave_shpr.div.b1\[7\] _04028_ _04024_ VGND VGND VPWR VPWR _04029_
+ sky130_fd_sc_hd__mux2_1
X_06692_ _01562_ _01573_ _01579_ _01581_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__or4b_1
XANTENNA__09180__S _03722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08431_ genblk2\[9\].wave_shpr.div.fin_quo\[2\] net32 _02262_ _02222_ VGND VGND VPWR
+ VPWR _03138_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12029__B2 genblk2\[10\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06900__B1 _01363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08362_ genblk2\[3\].wave_shpr.div.fin_quo\[5\] _02539_ _03068_ _02592_ VGND VGND
+ VPWR VPWR _03069_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11788__B1 _03693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07313_ _01308_ _01439_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__nand2_2
X_08293_ _02921_ _02997_ _02992_ _02996_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_73_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout136_A net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07244_ _01990_ _01991_ _02009_ _02010_ _02025_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_27_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07929__A _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07175_ _01953_ _01967_ _01968_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
X_06126_ _01097_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08708__B2 _02468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10802__B _04880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09816_ _04058_ _01410_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__nor2_1
X_09747_ genblk2\[2\].wave_shpr.div.fin_quo\[6\] genblk2\[2\].wave_shpr.div.quo\[5\]
+ _00009_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__mux2_1
XANTENNA__12268__A1 _01589_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06959_ genblk1\[7\].osc.clkdiv_C.cnt\[0\] net34 genblk1\[7\].osc.clkdiv_C.cnt\[10\]
+ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__and3b_1
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ genblk2\[2\].wave_shpr.div.acc\[15\] genblk2\[2\].wave_shpr.div.b1\[15\]
+ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__or2b_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout49_A net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _02734_ _02735_ genblk2\[6\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR
+ _03336_ sky130_fd_sc_hd__a21oi_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _05413_ _05416_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11571_ _05488_ _05383_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__xnor2_1
X_13310_ clknet_leaf_118_clk net272 net137 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10522_ _04754_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10453_ net1340 _04703_ _04704_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__mux2_1
X_13241_ clknet_leaf_10_clk _00564_ net55 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13172_ clknet_leaf_128_clk _00497_ net66 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10384_ net672 _04657_ _04655_ genblk2\[4\].wave_shpr.div.quo\[9\] _04659_ VGND VGND
+ VPWR VPWR _00469_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12123_ _05770_ _05736_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__or2b_1
X_12054_ net518 _05823_ _05825_ net547 _05831_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__a221o_1
X_11005_ net986 _05086_ _05056_ _05092_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__a22o_1
XANTENNA__06186__A1 _01155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12956_ clknet_leaf_136_clk _00285_ net42 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07135__B1 _01925_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11543__B genblk1\[8\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11907_ net273 _05729_ _03855_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__o21ai_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ clknet_leaf_30_clk _00218_ net96 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11838_ net807 _05652_ _05653_ _05680_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11769_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_40_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13508_ clknet_leaf_79_clk _00825_ net205 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13439_ clknet_leaf_94_clk _00758_ net162 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08980_ _01157_ _03664_ _03665_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__o21ai_1
X_07931_ net30 VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07862_ _02525_ _02567_ _02568_ _02361_ genblk2\[1\].wave_shpr.div.fin_quo\[2\] VGND
+ VGND VPWR VPWR _02569_ sky130_fd_sc_hd__a32o_1
X_09601_ net813 _04076_ _04080_ _04102_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__a22o_1
XANTENNA__07913__A2 _01309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06813_ genblk1\[5\].osc.clkdiv_C.cnt\[0\] _01684_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07793_ _02496_ _02497_ _02498_ _02499_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__and4_1
X_09532_ net519 _04052_ _04053_ net537 _04056_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__a221o_1
X_06744_ _01626_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07126__B1 _01855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire33 _02348_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_2
XFILLER_0_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08746__C genblk2\[6\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09463_ _04019_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__clkbuf_1
X_06675_ _01187_ _01564_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__nand2_4
X_08414_ genblk2\[2\].wave_shpr.div.fin_quo\[7\] _02468_ _03120_ _02592_ VGND VGND
+ VPWR VPWR _03121_ sky130_fd_sc_hd__a22o_1
X_09394_ genblk2\[1\].wave_shpr.div.acc\[13\] genblk2\[1\].wave_shpr.div.b1\[13\]
+ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__or2b_1
XFILLER_0_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08345_ _02993_ _02994_ _02995_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__nand3_1
XANTENNA__11225__A2 _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08276_ _02416_ _02982_ _02419_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__o21ai_2
XANTENNA__07659__A net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07227_ genblk1\[10\].osc.clkdiv_C.cnt\[5\] _01992_ _02008_ VGND VGND VPWR VPWR _02009_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06282__B _01242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07158_ _01954_ _01955_ _01956_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06109_ _01089_ VGND VGND VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.next_hzX sky130_fd_sc_hd__clkbuf_1
XANTENNA__07062__C1 _01490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07089_ net1185 _01897_ _01899_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__a21oi_1
Xfanout120 net122 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_2
XFILLER_0_100_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout131 net136 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_98_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_16
Xfanout142 net145 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08157__A2 _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout153 net155 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_4
Xfanout164 net165 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_4
Xfanout175 net176 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_4
Xfanout186 net188 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08562__C1 genblk2\[7\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout197 net198 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__buf_2
X_12810_ clknet_leaf_59_clk net299 net187 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12741_ clknet_leaf_49_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[0\] net108 VGND VGND
+ VPWR VPWR genblk1\[11\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08865__B1 _02248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ clknet_leaf_90_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[3\] net173 VGND VGND
+ VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_2
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ net1222 _05507_ _05445_ _05528_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_22_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11554_ _05374_ _05375_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06473__A genblk1\[1\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10505_ net472 _04715_ _04722_ _04743_ VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11485_ _03831_ net374 _03728_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12177__B1 _05818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13224_ clknet_leaf_114_clk _00547_ net132 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09784__A _01490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10436_ _04588_ _04691_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08396__A2 _01349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13155_ clknet_leaf_121_clk net627 net80 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10367_ _02152_ genblk2\[4\].wave_shpr.div.busy _02175_ VGND VGND VPWR VPWR _04653_
+ sky130_fd_sc_hd__and3_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _05762_ _05740_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__or2b_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ clknet_leaf_136_clk net943 net42 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10298_ genblk2\[4\].wave_shpr.div.b1\[14\] genblk2\[4\].wave_shpr.div.acc\[14\]
+ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__and2b_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_89_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_16
X_12037_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13388__RESET_B net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13317__RESET_B net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09024__A _02203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12939_ clknet_leaf_110_clk _00268_ net136 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10663__B1 _04857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06460_ genblk1\[1\].osc.clkdiv_C.cnt\[9\] _01392_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06391_ genblk1\[1\].osc.clkdiv_C.cnt\[10\] _01334_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_13_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08130_ _02819_ _02836_ genblk1\[4\].osc.clkdiv_C.cnt\[16\] genblk1\[4\].osc.clkdiv_C.cnt\[17\]
+ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_83_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09281__B1 _03840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08061_ genblk1\[5\].osc.clkdiv_C.cnt\[4\] net36 _02767_ VGND VGND VPWR VPWR _02768_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07012_ _01823_ _01837_ _01838_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_24_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09033__B1 _03702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07595__B1 genblk1\[9\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08963_ _03559_ _03563_ _03564_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07914_ genblk1\[8\].osc.clkdiv_C.cnt\[3\] _01866_ _02619_ _01489_ _02620_ VGND VGND
+ VPWR VPWR _02621_ sky130_fd_sc_hd__o221a_1
X_08894_ net629 _02260_ _03599_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__a21o_1
X_07845_ net18 VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__buf_2
XFILLER_0_75_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07898__B2 genblk1\[8\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07776_ _01229_ _01359_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__nand2_1
X_09515_ genblk2\[1\].wave_shpr.div.quo\[5\] _04043_ _04047_ net414 VGND VGND VPWR
+ VPWR _00212_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06727_ genblk1\[4\].osc.clkdiv_C.cnt\[4\] _01609_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06277__B _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10654__B1 _04821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09446_ genblk2\[1\].wave_shpr.div.acc\[25\] genblk2\[1\].wave_shpr.div.acc\[26\]
+ _04009_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__or3_2
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06658_ genblk1\[3\].osc.clkdiv_C.cnt\[15\] genblk1\[3\].osc.clkdiv_C.cnt\[14\] _01547_
+ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__and3_1
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06873__A2 _01726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09377_ genblk2\[11\].wave_shpr.div.i\[1\] genblk2\[11\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _03945_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06589_ _01191_ _01233_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08328_ _02688_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06293__A _01196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08259_ _02848_ _02894_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__xor2_2
XFILLER_0_104_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11270_ genblk2\[7\].wave_shpr.div.b1\[0\] _05182_ _05183_ VGND VGND VPWR VPWR _05276_
+ sky130_fd_sc_hd__and3_1
X_10221_ genblk2\[3\].wave_shpr.div.acc\[20\] _04541_ VGND VGND VPWR VPWR _04544_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10152_ _04385_ _04491_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10083_ _02170_ genblk2\[3\].wave_shpr.div.busy _02167_ VGND VGND VPWR VPWR _04453_
+ sky130_fd_sc_hd__and3_1
Xhold9 _00888_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13773_ clknet_leaf_74_clk _01084_ net213 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10985_ _05074_ genblk1\[6\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12724_ clknet_leaf_37_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[1\] net113 VGND VGND
+ VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12655_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[4\] net90 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__10718__A _04856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08066__A1 _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11606_ genblk2\[8\].wave_shpr.div.acc\[13\] _05515_ _05493_ VGND VGND VPWR VPWR
+ _05516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12586_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[7\] net74 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09802__A2 _04248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11537_ _05464_ genblk1\[8\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold409 _00480_ VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11468_ net1208 _01811_ _05237_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__mux2_1
X_13207_ clknet_leaf_25_clk _00530_ net86 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10419_ _04654_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11399_ genblk2\[8\].wave_shpr.div.acc\[0\] genblk2\[8\].wave_shpr.div.b1\[0\] VGND
+ VGND VPWR VPWR _05375_ sky130_fd_sc_hd__and2b_1
XFILLER_0_110_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ clknet_leaf_115_clk net733 net135 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ clknet_leaf_24_clk net546 net93 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1109 genblk2\[2\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net1327 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08541__A2 _02526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07630_ genblk1\[11\].osc.clkdiv_C.cnt\[8\] _02336_ net34 VGND VGND VPWR VPWR _02337_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06378__A net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07561_ genblk1\[9\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09300_ _03776_ _03887_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__xnor2_1
X_06512_ genblk1\[2\].osc.clkdiv_C.cnt\[6\] _01437_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__xor2_1
X_07492_ _02214_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10100__A2 _04457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09231_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__and2_1
X_06443_ genblk1\[1\].osc.clkdiv_C.cnt\[4\] _01380_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06825__B genblk1\[5\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09162_ _03807_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__clkbuf_1
X_06374_ _01307_ _01311_ _01312_ genblk1\[1\].osc.clkdiv_C.cnt\[11\] _01317_ VGND
+ VGND VPWR VPWR _01318_ sky130_fd_sc_hd__o221a_1
XFILLER_0_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08113_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01323_ _01592_ genblk1\[4\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_32_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09093_ _01367_ _03739_ _03741_ _01342_ _03742_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout216_A net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08044_ _01181_ _01680_ _02749_ _02750_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__o211ai_1
Xhold910 PWM.final_in\[7\] VGND VGND VPWR VPWR net1128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 genblk2\[0\].wave_shpr.div.acc\[2\] VGND VGND VPWR VPWR net1139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 PWM.final_in\[4\] VGND VGND VPWR VPWR net1150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold943 sig_norm.b1\[0\] VGND VGND VPWR VPWR net1161 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10363__A _03833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold954 PWM.final_in\[3\] VGND VGND VPWR VPWR net1172 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07656__B _02362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold965 genblk1\[10\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR net1183 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__B1 _01246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold976 genblk1\[9\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR net1194 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold987 genblk2\[4\].wave_shpr.div.b1\[12\] VGND VGND VPWR VPWR net1205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 _05230_ VGND VGND VPWR VPWR net1216 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ genblk2\[3\].wave_shpr.div.b1\[6\] genblk2\[3\].wave_shpr.div.acc\[6\] VGND
+ VGND VPWR VPWR _04391_ sky130_fd_sc_hd__and2b_1
X_08946_ _03637_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12313__B1 _03944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07672__A _01308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08877_ _03577_ _03581_ _03582_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11194__A _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07828_ _02533_ _02534_ _02518_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06288__A _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07740__B1 _01356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07759_ genblk2\[1\].wave_shpr.div.fin_quo\[5\] _02461_ _02464_ _02224_ VGND VGND
+ VPWR VPWR _02466_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12092__A2 _05844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10770_ _04809_ _04929_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09429_ _03960_ _03991_ _03992_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12440_ _06099_ _05980_ genblk2\[11\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR
+ _06101_ sky130_fd_sc_hd__mux2_1
X_12371_ _05953_ _05936_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__or2b_1
XFILLER_0_151_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11322_ _05207_ _05168_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__or2b_1
XFILLER_0_105_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11253_ genblk2\[7\].wave_shpr.div.quo\[20\] _05255_ _05256_ net231 _05266_ VGND
+ VGND VPWR VPWR _00731_ sky130_fd_sc_hd__a221o_1
XANTENNA__07559__B1 _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06470__B genblk1\[1\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10204_ net1016 _04518_ _04522_ _04531_ VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__a22o_1
X_11184_ _05232_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__clkbuf_1
X_10135_ genblk2\[3\].wave_shpr.div.acc_next\[0\] _04455_ VGND VGND VPWR VPWR _04479_
+ sky130_fd_sc_hd__or2b_1
XANTENNA__07574__A3 _01226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12304__B1 _06010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07582__A genblk1\[9\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10066_ net1192 _04229_ _04440_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13756_ clknet_leaf_69_clk _01067_ net212 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12083__A2 _05844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10968_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__and2_1
XANTENNA__10094__A1 net401 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06298__B1 _01240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12707_ clknet_leaf_56_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[2\] net181 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13687_ clknet_leaf_63_clk _01000_ net191 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10899_ _03687_ _05033_ _04233_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12638_ clknet_leaf_19_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[5\] net109 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_155_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09787__A1 _01365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12569_ clknet_leaf_27_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[8\] net90 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09448__S _00007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold206 genblk2\[11\].wave_shpr.div.b1\[15\] VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold217 _01057_ VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold228 genblk2\[10\].wave_shpr.div.quo\[24\] VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11279__A _05249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold239 genblk2\[2\].wave_shpr.div.quo\[13\] VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _03450_ _03449_ _03427_ _03422_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__o211a_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06222__B1 _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08762__A2 _02539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ net1285 _01858_ _04238_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__mux2_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06992_ net1252 net1058 genblk1\[7\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR _01826_
+ sky130_fd_sc_hd__a21oi_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07492__A _02214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08731_ _03433_ _03437_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__xnor2_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08662_ genblk2\[5\].wave_shpr.div.fin_quo\[2\] _03367_ _03368_ VGND VGND VPWR VPWR
+ _03369_ sky130_fd_sc_hd__o21a_1
XANTENNA__07722__B1 _01591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07613_ genblk1\[11\].osc.clkdiv_C.cnt\[1\] _01186_ _01354_ _01321_ genblk1\[11\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__o311a_1
X_08593_ genblk2\[4\].wave_shpr.div.fin_quo\[0\] _02526_ _02361_ genblk2\[4\].wave_shpr.div.fin_quo\[1\]
+ _02838_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout166_A net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07544_ _02255_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10085__A1 net794 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10085__B2 _04454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07475_ _02155_ _02202_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__nor2_4
XFILLER_0_45_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09214_ _03835_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06426_ _01197_ _01364_ _01368_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] _01369_ VGND VGND
+ VPWR VPWR _01370_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09227__B1 _03840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09778__A1 _01487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09145_ genblk2\[0\].wave_shpr.div.b1\[15\] genblk2\[0\].wave_shpr.div.acc\[15\]
+ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06357_ freq_div.state\[2\] freq_div.state\[0\] VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__and2b_1
XANTENNA__07667__A _01308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09076_ net1291 _01483_ _03722_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__mux2_1
X_06288_ _01248_ _01249_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__nor2_2
XANTENNA__08450__B2 _02521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08027_ _02733_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__buf_2
XFILLER_0_130_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold740 genblk2\[11\].wave_shpr.div.acc\[5\] VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 genblk2\[10\].wave_shpr.div.acc\[3\] VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold762 genblk2\[8\].wave_shpr.div.acc\[4\] VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold773 genblk2\[8\].wave_shpr.div.acc\[17\] VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 genblk2\[2\].wave_shpr.div.acc\[14\] VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 genblk2\[7\].wave_shpr.div.acc\[2\] VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13073__RESET_B net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06425__A1_N genblk1\[1\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09978_ genblk2\[3\].wave_shpr.div.b1\[4\] genblk2\[3\].wave_shpr.div.acc\[4\] VGND
+ VGND VPWR VPWR _04374_ sky130_fd_sc_hd__or2b_1
XANTENNA_fanout79_A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08929_ sig_norm.acc\[10\] _03622_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__and2b_1
X_11940_ genblk2\[10\].wave_shpr.div.b1\[8\] genblk2\[10\].wave_shpr.div.acc\[8\]
+ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11871_ _05704_ _05705_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13610_ clknet_leaf_93_clk _00923_ net159 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10822_ genblk2\[6\].wave_shpr.div.acc\[17\] genblk2\[6\].wave_shpr.div.b1\[17\]
+ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__or2b_1
XFILLER_0_67_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13541_ clknet_leaf_101_clk _00856_ net165 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11273__B1 _05250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10753_ genblk2\[5\].wave_shpr.div.acc\[11\] _04916_ _04907_ VGND VGND VPWR VPWR
+ _04917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06465__B genblk1\[1\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09218__B1 _03804_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13472_ clknet_leaf_74_clk _00789_ net212 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10684_ _04268_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_137_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06184__C _01096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12423_ _05976_ net20 genblk2\[11\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR _06090_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_124_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08441__A1 _02525_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12354_ _05944_ _06036_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07244__A2 _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11305_ _05198_ _05302_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10207__S _04507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12285_ _03702_ net1121 VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__nor2_1
X_11236_ genblk2\[7\].wave_shpr.div.quo\[12\] _05255_ _05256_ net370 _05257_ VGND
+ VGND VPWR VPWR _00723_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold7_A modein.delay_octave_down_in\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11167_ genblk2\[7\].wave_shpr.div.fin_quo\[2\] net1311 _00019_ VGND VGND VPWR VPWR
+ _05225_ sky130_fd_sc_hd__mux2_1
X_10118_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__and2_1
XANTENNA__08201__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11098_ _05055_ _05158_ _05160_ _05057_ net739 VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__a32o_1
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10049_ _04433_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06359__C _01302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09032__A _03701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13739_ clknet_leaf_46_clk _01050_ net119 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09209__B1 _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07260_ _02028_ _02036_ _02037_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06211_ freq_div.state\[0\] VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__06691__B1 _01498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07191_ genblk1\[9\].osc.clkdiv_C.cnt\[12\] _01978_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10906__A _01805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_83_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06142_ net2 VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__inv_2
XANTENNA__09178__S _03722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06391__A genblk1\[1\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08432__B2 _02308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09901_ _04197_ _04161_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__or2b_1
XFILLER_0_1_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_98_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08196__B1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ net322 _04257_ _04259_ net339 _04266_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__a221o_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10641__A _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _04231_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__clkbuf_1
X_06975_ _01365_ _01355_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__nor2_4
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08714_ _03408_ _03419_ _03418_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__a21oi_2
X_09694_ _04172_ _04173_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _03349_ _03350_ _03340_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07171__A1 genblk1\[9\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11472__A _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08576_ _02525_ _03281_ _03282_ _02361_ genblk2\[11\].wave_shpr.div.fin_quo\[2\]
+ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07527_ sig_norm.i\[1\] _02243_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07458_ genblk2\[7\].wave_shpr.div.i\[2\] genblk2\[7\].wave_shpr.div.i\[3\] genblk2\[7\].wave_shpr.div.i\[4\]
+ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_17_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06682__B1 _01340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06409_ _01338_ _01339_ _01346_ _01352_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__or4b_1
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07389_ _02081_ _02136_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09128_ _03757_ _03774_ _03775_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09059_ _01229_ genblk2\[0\].wave_shpr.div.b1\[8\] _03719_ VGND VGND VPWR VPWR _03720_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12070_ _05815_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__inv_2
Xhold570 genblk2\[2\].wave_shpr.div.acc\[17\] VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 genblk2\[9\].wave_shpr.div.acc\[14\] VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 PWM.counter\[5\] VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ _05022_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12972_ clknet_leaf_125_clk _00301_ net71 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11923_ genblk2\[10\].wave_shpr.div.acc\[2\] genblk2\[10\].wave_shpr.div.b1\[2\]
+ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__or2b_1
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11854_ _05599_ _05692_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12038__A2 _05818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ genblk2\[5\].wave_shpr.div.acc\[25\] _04953_ VGND VGND VPWR VPWR _04955_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11785_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13524_ clknet_leaf_98_clk _00841_ net169 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10736_ genblk2\[5\].wave_shpr.div.acc\[7\] _04903_ _04821_ VGND VGND VPWR VPWR _04904_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13455_ clknet_leaf_99_clk _00772_ net168 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_10667_ net310 _04858_ _04855_ net423 _04859_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12406_ _05969_ _05928_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__or2b_1
XFILLER_0_152_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07217__A2 _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08414__B2 _02592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13386_ clknet_leaf_86_clk _00705_ net183 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10598_ genblk2\[5\].wave_shpr.div.fin_quo\[2\] net1336 _00015_ VGND VGND VPWR VPWR
+ _04824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06425__B1 _01340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12337_ net438 _03942_ _03941_ net504 _06026_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12268_ net1235 _01589_ _05994_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__mux2_1
X_11219_ genblk2\[7\].wave_shpr.div.quo\[2\] _05246_ _05250_ net563 VGND VGND VPWR
+ VPWR _00713_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12199_ genblk2\[11\].wave_shpr.div.acc\[5\] genblk2\[11\].wave_shpr.div.b1\[5\]
+ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__or2b_1
X_06760_ _01599_ _01636_ _01638_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06691_ genblk1\[4\].osc.clkdiv_C.cnt\[0\] _01210_ _01498_ genblk1\[4\].osc.clkdiv_C.cnt\[14\]
+ _01580_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__o221a_1
XANTENNA__08350__B1 _02527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08430_ _02303_ _02262_ genblk2\[9\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR
+ _03137_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12029__A2 _05813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08361_ genblk2\[3\].wave_shpr.div.fin_quo\[4\] _03067_ VGND VGND VPWR VPWR _03068_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07312_ genblk1\[11\].osc.clkdiv_C.cnt\[14\] _01210_ _01578_ genblk1\[11\].osc.clkdiv_C.cnt\[16\]
+ _02075_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__o221a_1
XANTENNA__13765__RESET_B net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08292_ _02945_ _02967_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07243_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _01235_ _02020_ _02022_ _02024_ VGND
+ VGND VPWR VPWR _02025_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07929__B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07174_ genblk1\[9\].osc.clkdiv_C.cnt\[6\] _01965_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06125_ _01094_ _01095_ _01096_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__nor3_2
XFILLER_0_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10371__A _04654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09815_ _04247_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__clkbuf_4
X_09746_ _04220_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__clkbuf_1
X_06958_ _01228_ _01220_ _01233_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__a21oi_4
XANTENNA__07680__A _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ genblk2\[2\].wave_shpr.div.acc\[16\] genblk2\[2\].wave_shpr.div.b1\[16\]
+ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__or2b_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06889_ genblk1\[6\].osc.clkdiv_C.cnt\[12\] _01519_ _01742_ genblk1\[6\].osc.clkdiv_C.cnt\[10\]
+ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12298__A _03941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _03275_ _03276_ _03295_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__nand3_2
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06296__A _01238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11228__B1 _05248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08559_ _03264_ _03265_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__nor2_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11570_ _05384_ _05370_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__or2b_1
XFILLER_0_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10521_ _04654_ _04651_ genblk2\[4\].wave_shpr.div.i\[0\] VGND VGND VPWR VPWR _04754_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13240_ clknet_leaf_11_clk net234 net57 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10452_ _04622_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13171_ clknet_leaf_126_clk _00496_ net66 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10383_ _04058_ _01568_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__nor2_1
X_12122_ net957 _05876_ _05850_ _05879_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__a22o_1
X_12053_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__and2_1
X_11004_ genblk2\[6\].wave_shpr.div.acc\[3\] _05091_ _05023_ VGND VGND VPWR VPWR _05092_
+ sky130_fd_sc_hd__mux2_1
X_12955_ clknet_leaf_136_clk _00284_ net62 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07135__A1 genblk1\[9\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07135__B2 genblk1\[9\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11906_ _03690_ _05728_ _05729_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__nor3_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12886_ clknet_leaf_30_clk _00217_ net98 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11219__B1 _05250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11837_ genblk2\[9\].wave_shpr.div.acc\[10\] _05679_ _05673_ VGND VGND VPWR VPWR
+ _05680_ sky130_fd_sc_hd__mux2_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ net485 _05628_ _05629_ net541 _05633_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10719_ _04787_ _04779_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__or2b_1
X_13507_ clknet_leaf_80_clk _00824_ net205 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11699_ _05562_ _05589_ _05590_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13438_ clknet_leaf_95_clk _00757_ net159 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13369_ clknet_leaf_116_clk _00688_ net140 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09456__S _00007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07930_ genblk2\[8\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__inv_2
XANTENNA__07484__B _02153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07861_ genblk2\[1\].wave_shpr.div.fin_quo\[0\] _02458_ _02459_ genblk2\[1\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__a31o_1
X_09600_ genblk2\[1\].wave_shpr.div.acc\[9\] _04101_ _04095_ VGND VGND VPWR VPWR _04102_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08571__B1 _02316_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06812_ _01189_ _01678_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__nor2_2
XANTENNA__07913__A3 _01855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07792_ _01246_ _01439_ _01344_ _01169_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__a31o_1
X_09531_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__and2_1
X_06743_ _01599_ _01624_ _01625_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__and3_1
XANTENNA__07126__A1 genblk1\[9\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07126__B2 genblk1\[9\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09462_ genblk2\[1\].wave_shpr.div.fin_quo\[7\] genblk2\[1\].wave_shpr.div.quo\[6\]
+ _00007_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__mux2_1
X_06674_ _01563_ VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__buf_6
XFILLER_0_66_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08413_ genblk2\[2\].wave_shpr.div.fin_quo\[6\] _03119_ VGND VGND VPWR VPWR _03120_
+ sky130_fd_sc_hd__xnor2_1
X_09393_ genblk2\[1\].wave_shpr.div.acc\[14\] genblk2\[1\].wave_shpr.div.b1\[14\]
+ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__or2b_1
XFILLER_0_93_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08344_ _03048_ _03049_ _03050_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__and3_2
XFILLER_0_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07659__B _02364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08275_ genblk2\[10\].wave_shpr.div.fin_quo\[5\] _02361_ _02980_ _02981_ VGND VGND
+ VPWR VPWR _02982_ sky130_fd_sc_hd__a22o_1
XANTENNA__10366__A _04651_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10984__A2 _05051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07226_ genblk1\[10\].osc.clkdiv_C.cnt\[5\] _01992_ _02007_ VGND VGND VPWR VPWR _02008_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07157_ genblk1\[9\].osc.clkdiv_C.cnt\[1\] genblk1\[9\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01956_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06108_ net1179 net395 _01088_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07088_ genblk1\[8\].osc.clkdiv_C.cnt\[7\] _01897_ _01886_ VGND VGND VPWR VPWR _01899_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_100_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout110 net111 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_4
Xfanout121 net122 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_4
Xfanout132 net133 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_4
Xfanout143 net145 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_4
Xfanout154 net155 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__buf_2
Xfanout165 net170 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_4
Xfanout176 net218 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
Xfanout187 net188 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_4
Xfanout198 net218 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_2
XFILLER_0_97_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09729_ genblk2\[2\].wave_shpr.div.acc\[18\] _04208_ VGND VGND VPWR VPWR _04209_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_97_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12740_ clknet_leaf_48_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[17\] net119 VGND
+ VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07668__A2 _02374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ clknet_leaf_89_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[2\] net173 VGND VGND
+ VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ genblk2\[8\].wave_shpr.div.acc\[17\] _05527_ _05416_ VGND VGND VPWR VPWR
+ _05528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09814__B1 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11553_ genblk2\[8\].wave_shpr.div.acc\[1\] _05416_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10504_ genblk2\[4\].wave_shpr.div.acc\[20\] _04740_ VGND VGND VPWR VPWR _04743_
+ sky130_fd_sc_hd__xnor2_1
X_11484_ _03727_ _01490_ _03687_ net478 VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12177__A1 _05816_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13223_ clknet_leaf_114_clk _00546_ net132 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10435_ _04589_ _04581_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07053__B1 _01870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13154_ clknet_leaf_121_clk _00479_ net77 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10366_ _04651_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__buf_2
X_12105_ net954 _05844_ _05850_ _05866_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__a22o_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06800__B1 _01666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13085_ clknet_leaf_135_clk _00412_ net62 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10297_ _04569_ _04607_ _04608_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__a21o_1
X_12036_ net398 _05818_ _05816_ net432 _05821_ VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__a221o_1
XANTENNA__08553__B1 _02261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12938_ clknet_leaf_111_clk _00267_ net136 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10663__A1 net308 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ clknet_leaf_134_clk _00200_ net60 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06390_ _01333_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09805__B1 _04252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09040__A _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08060_ genblk1\[5\].osc.clkdiv_C.cnt\[5\] _01238_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07011_ genblk1\[7\].osc.clkdiv_C.cnt\[9\] _01835_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07495__A _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08962_ _03507_ _03451_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__nor2_1
XANTENNA__08103__B _01574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07913_ genblk1\[8\].osc.clkdiv_C.cnt\[0\] _01309_ _01855_ genblk1\[8\].osc.clkdiv_C.cnt\[1\]
+ genblk1\[8\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__a311o_1
X_08893_ _01099_ _03574_ _03598_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout196_A net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07844_ genblk2\[0\].wave_shpr.div.fin_quo\[2\] _02549_ _02550_ VGND VGND VPWR VPWR
+ _02551_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09215__A _02152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07775_ genblk1\[0\].osc.clkdiv_C.cnt\[2\] _01227_ _02479_ _02480_ _02481_ VGND VGND
+ VPWR VPWR _02482_ sky130_fd_sc_hd__o221a_1
X_09514_ net414 _04043_ _04047_ net701 VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06726_ _01612_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09445_ genblk2\[1\].wave_shpr.div.acc\[24\] _04008_ VGND VGND VPWR VPWR _04009_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_148_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10654__B2 _04855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06657_ net1195 _01547_ _01550_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09376_ _03940_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__clkbuf_4
X_06588_ _01437_ _01225_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__or2_4
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12296__B1_N _03735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08327_ genblk2\[8\].wave_shpr.div.fin_quo\[5\] _02467_ _03033_ _02636_ VGND VGND
+ VPWR VPWR _03034_ sky130_fd_sc_hd__a211o_1
XANTENNA__10096__A _04451_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08075__A2 _01678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09272__B2 _03836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08258_ _02958_ _02963_ _02964_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_62_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07209_ _01556_ _01564_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__nand2_8
X_08189_ _02849_ _02894_ _02895_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10220_ genblk2\[3\].wave_shpr.div.acc\[20\] _04541_ VGND VGND VPWR VPWR _04543_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_42_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07035__B1 _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10151_ _04386_ _04377_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__or2b_1
XFILLER_0_30_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10082_ _04451_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07571__C _01355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13772_ clknet_leaf_73_clk _01083_ net215 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_2
X_10984_ genblk2\[6\].wave_shpr.div.quo\[24\] _05051_ _05054_ net385 _05077_ VGND
+ VGND VPWR VPWR _00651_ sky130_fd_sc_hd__a221o_1
XFILLER_0_139_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10645__A1 _01365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12723_ clknet_leaf_37_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[0\] net113 VGND VGND
+ VPWR VPWR genblk1\[10\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12654_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[3\] net90 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11605_ _05399_ _05514_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07299__B _01235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12585_ clknet_leaf_124_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[6\] net76 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_111_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09795__A _02152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11536_ net660 _05454_ _05458_ net677 _05465_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11740__A1_N _01099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11467_ _05430_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13206_ clknet_leaf_25_clk _00529_ net88 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10418_ net643 _04651_ _04654_ genblk2\[4\].wave_shpr.div.quo\[24\] _04678_ VGND
+ VGND VPWR VPWR _00484_ sky130_fd_sc_hd__a221o_1
XANTENNA__09566__A2 _04043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11398_ genblk2\[8\].wave_shpr.div.acc\[1\] genblk2\[8\].wave_shpr.div.b1\[1\] VGND
+ VGND VPWR VPWR _05374_ sky130_fd_sc_hd__xor2_1
X_13137_ clknet_leaf_115_clk _00462_ net135 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ net1266 _01757_ _04637_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__mux2_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ clknet_leaf_24_clk net297 net93 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11565__A _05444_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12019_ _05814_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10333__B1 _01262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09035__A _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07560_ genblk1\[9\].osc.clkdiv_C.cnt\[13\] _01245_ _01328_ genblk1\[9\].osc.clkdiv_C.cnt\[12\]
+ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__o22a_1
X_06511_ _01332_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07491_ _02211_ _02152_ genblk2\[11\].wave_shpr.div.busy VGND VGND VPWR VPWR _02214_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_76_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06304__A2 _01235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09230_ genblk2\[0\].wave_shpr.div.quo\[9\] _03841_ _03839_ net277 _03842_ VGND VGND
+ VPWR VPWR _00132_ sky130_fd_sc_hd__a221o_1
X_06442_ genblk1\[1\].osc.clkdiv_C.cnt\[4\] _01380_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09161_ genblk2\[0\].wave_shpr.div.fin_quo\[2\] net1322 _00001_ VGND VGND VPWR VPWR
+ _03807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06373_ genblk1\[1\].osc.clkdiv_C.cnt\[2\] _01240_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08112_ _02804_ _02806_ _02808_ _02817_ _02818_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__o221a_1
X_09092_ _01367_ _03740_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08043_ genblk1\[5\].osc.clkdiv_C.cnt\[14\] _01360_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout111_A net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold900 genblk2\[10\].wave_shpr.div.acc\[1\] VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 genblk2\[4\].wave_shpr.div.acc\[1\] VGND VGND VPWR VPWR net1129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold922 genblk2\[7\].wave_shpr.div.b1\[1\] VGND VGND VPWR VPWR net1140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout209_A net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12010__B1 _03733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold933 _03682_ VGND VGND VPWR VPWR net1151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 genblk1\[8\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR net1162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 genblk2\[10\].wave_shpr.div.b1\[6\] VGND VGND VPWR VPWR net1173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 genblk2\[0\].wave_shpr.div.b1\[10\] VGND VGND VPWR VPWR net1184 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__B2 genblk1\[9\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold977 genblk1\[3\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR net1195 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ _04373_ _04388_ _04389_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__a21o_1
Xhold988 genblk2\[4\].wave_shpr.div.b1\[8\] VGND VGND VPWR VPWR net1206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 genblk2\[11\].wave_shpr.div.b1\[9\] VGND VGND VPWR VPWR net1217 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06240__A1 _01201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08945_ sig_norm.quo\[2\] _03636_ _00024_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__mux2_1
X_08876_ sig_norm.b1\[2\] sig_norm.acc\[2\] VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__xor2_1
X_07827_ genblk2\[0\].wave_shpr.div.fin_quo\[4\] _02309_ _02509_ VGND VGND VPWR VPWR
+ _02534_ sky130_fd_sc_hd__a21o_1
XANTENNA__06288__B _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07740__A1 genblk1\[1\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13208__RESET_B net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07740__B2 genblk1\[1\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07758_ _02461_ _02464_ genblk2\[1\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR
+ _02465_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06709_ _01558_ _01560_ _01584_ _01598_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__or4_4
XANTENNA__09493__A1 _04036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07689_ genblk1\[10\].osc.clkdiv_C.cnt\[10\] _02005_ _02394_ _02395_ VGND VGND VPWR
+ VPWR _02396_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_66_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09428_ genblk2\[1\].wave_shpr.div.b1\[11\] genblk2\[1\].wave_shpr.div.acc\[11\]
+ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__and2b_1
XFILLER_0_125_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09359_ net933 _03903_ _03910_ _03932_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12370_ net841 _06039_ _06040_ _06049_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11321_ _05249_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11252_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__and2_1
XANTENNA__07559__A1 _01200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10203_ genblk2\[3\].wave_shpr.div.acc\[15\] _04530_ _04507_ VGND VGND VPWR VPWR
+ _04531_ sky130_fd_sc_hd__mux2_1
X_11183_ net1214 _04242_ _05042_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10134_ genblk2\[3\].wave_shpr.div.acc_next\[0\] _04451_ _04455_ net561 _04478_ VGND
+ VGND VPWR VPWR _00400_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10065_ _04442_ VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09484__A1 _01302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10967_ net595 _05062_ _05064_ net594 _05068_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__a221o_1
X_13755_ clknet_leaf_68_clk _01066_ net212 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06298__A1 genblk1\[0\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10094__A2 _04452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12706_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[1\] net183 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
X_13686_ clknet_leaf_63_clk _00999_ net191 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10898_ net1140 VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12637_ clknet_leaf_16_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[4\] net73 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12568_ clknet_leaf_27_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[7\] net90 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_135_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11519_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12499_ clknet_leaf_103_clk _00061_ net156 VGND VGND VPWR VPWR sig_norm.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold207 genblk2\[1\].wave_shpr.div.b1\[16\] VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold218 genblk1\[3\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__buf_1
XFILLER_0_124_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold229 _00973_ VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09464__S _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06222__A1 _01172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ genblk1\[7\].osc.clkdiv_C.cnt\[2\] genblk1\[7\].osc.clkdiv_C.cnt\[1\] genblk1\[7\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__and3_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08730_ _03114_ _03436_ _03122_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__o21a_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06389__A _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08661_ _03176_ _02789_ _03177_ _02525_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__o31a_1
X_07612_ _01186_ _01354_ genblk1\[11\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _02319_
+ sky130_fd_sc_hd__o21a_1
X_08592_ genblk2\[5\].wave_shpr.div.fin_quo\[0\] _02527_ _02521_ genblk2\[5\].wave_shpr.div.fin_quo\[1\]
+ _02791_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07543_ PWM.final_sample_in\[3\] net1172 PWM.start VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09475__A1 _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12074__A3 _05787_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10085__A2 _04452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07474_ genblk2\[9\].wave_shpr.div.busy _02201_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__and2_2
X_09213_ _02151_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__buf_2
X_06425_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] _01368_ _01340_ genblk1\[1\].osc.clkdiv_C.cnt\[1\]
+ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_146_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09144_ _03749_ _03790_ _03791_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__a21o_1
X_06356_ genblk1\[0\].osc.clkdiv_C.cnt\[17\] _01298_ _01300_ _01270_ VGND VGND VPWR
+ VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[17\] sky130_fd_sc_hd__o211a_1
XFILLER_0_32_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09075_ _03730_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06287_ _01173_ _01188_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__nor2_4
XFILLER_0_114_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08026_ _02712_ _02731_ _02732_ VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__o21a_4
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold730 genblk2\[3\].wave_shpr.div.acc\[17\] VGND VGND VPWR VPWR net948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 genblk2\[10\].wave_shpr.div.b1\[16\] VGND VGND VPWR VPWR net959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold752 genblk2\[4\].wave_shpr.div.acc\[5\] VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 genblk2\[5\].wave_shpr.div.acc\[13\] VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold774 genblk2\[7\].wave_shpr.div.acc\[3\] VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_889 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold785 genblk2\[6\].wave_shpr.div.acc\[10\] VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 genblk2\[5\].wave_shpr.div.acc\[12\] VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07683__A _01174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09950__A2 _04253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09977_ genblk2\[3\].wave_shpr.div.acc\[5\] genblk2\[3\].wave_shpr.div.b1\[5\] VGND
+ VGND VPWR VPWR _04373_ sky130_fd_sc_hd__or2b_1
XANTENNA__06407__A2_N _01349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08928_ net663 _02260_ _03624_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08859_ _03427_ _03505_ _03500_ _03504_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__a211oi_1
X_11870_ _05607_ _05646_ genblk2\[9\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR
+ _05705_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10821_ net856 _04965_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09466__A1 _01327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10752_ _04801_ _04915_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__xnor2_1
X_13540_ clknet_leaf_101_clk _00855_ net164 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13471_ clknet_leaf_75_clk _00788_ net204 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10683_ net378 _04861_ _04862_ net551 _04868_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__a221o_1
XANTENNA__09218__A1 net804 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09218__B2 _03839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12422_ _05977_ net20 VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07858__A _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12353_ genblk2\[11\].wave_shpr.div.b1\[2\] genblk2\[11\].wave_shpr.div.acc\[2\]
+ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__xor2_1
X_11304_ _05199_ _05172_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__or2b_1
XFILLER_0_133_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12284_ _06003_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11235_ _05074_ genblk1\[7\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09284__S _03804_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09941__A2 _04253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11166_ _05224_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__clkbuf_1
X_10117_ genblk2\[3\].wave_shpr.div.quo\[17\] _04461_ _04462_ net376 _04469_ VGND
+ VGND VPWR VPWR _00392_ sky130_fd_sc_hd__a221o_1
X_11097_ _05159_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__inv_2
X_10048_ genblk2\[4\].wave_shpr.div.b1\[3\] _01223_ _04238_ VGND VGND VPWR VPWR _04433_
+ sky130_fd_sc_hd__mux2_1
Xhold90 genblk2\[5\].wave_shpr.div.quo\[7\] VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_89_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11843__A _02203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11999_ _03687_ net420 _03705_ VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__a21bo_1
X_13738_ clknet_leaf_46_clk net352 net119 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09209__A1 _03714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13669_ clknet_leaf_41_clk _00982_ net125 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_06210_ _01171_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__clkbuf_8
X_07190_ _01953_ _01977_ _01978_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_14_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06141_ net14 _01112_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06391__B _01334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09900_ _04247_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08599__A net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09194__S _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__and2_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ net1290 _04230_ _04039_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__mux2_1
X_06974_ genblk1\[7\].osc.clkdiv_C.cnt\[14\] _01675_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__xor2_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _03408_ _03418_ _03419_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__and3_2
X_09693_ genblk2\[2\].wave_shpr.div.acc\[1\] genblk2\[2\].wave_shpr.div.b1\[1\] VGND
+ VGND VPWR VPWR _04173_ sky130_fd_sc_hd__or2b_1
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08644_ _03340_ _03349_ _03350_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__nand3_1
XFILLER_0_96_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08575_ genblk2\[11\].wave_shpr.div.fin_quo\[0\] genblk2\[11\].wave_shpr.div.fin_quo\[1\]
+ _02349_ _02351_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__nand4_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10369__A _04654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09448__A1 _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07526_ sig_norm.busy net939 _01099_ _02244_ VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08120__A1 _01224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07457_ _02189_ VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06408_ genblk1\[1\].osc.clkdiv_C.cnt\[3\] _01323_ _01347_ _01348_ _01351_ VGND VGND
+ VPWR VPWR _01352_ sky130_fd_sc_hd__o221a_1
XFILLER_0_146_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07388_ _02081_ _02136_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06582__A _01489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09127_ genblk2\[0\].wave_shpr.div.b1\[6\] genblk2\[0\].wave_shpr.div.acc\[6\] VGND
+ VGND VPWR VPWR _03775_ sky130_fd_sc_hd__and2b_1
X_06339_ genblk1\[0\].osc.clkdiv_C.cnt\[11\] genblk1\[0\].osc.clkdiv_C.cnt\[10\] _01286_
+ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09058_ _02170_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__buf_6
X_08009_ _02713_ _02714_ _02715_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__o21ba_1
Xhold560 genblk2\[4\].wave_shpr.div.acc\[12\] VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10518__B1 _04655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold571 genblk2\[9\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout91_A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold582 genblk2\[5\].wave_shpr.div.b1\[14\] VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ _04995_ _05103_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09384__B1 _03947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold593 _01165_ VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__dlygate4sd3_1
X_12971_ clknet_leaf_125_clk net301 net71 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11922_ genblk2\[10\].wave_shpr.div.acc\[3\] genblk2\[10\].wave_shpr.div.b1\[3\]
+ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__or2b_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _05600_ _05557_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__or2b_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06476__B genblk1\[1\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ net1041 _04858_ _04855_ _04954_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11784_ net226 _02203_ _03693_ net416 _05641_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__a221o_1
X_13523_ clknet_leaf_98_clk _00840_ net169 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10735_ _04793_ _04902_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13454_ clknet_leaf_99_clk _00771_ net164 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_10666_ _04672_ genblk1\[5\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__and2_1
XANTENNA__06492__A _01229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12405_ net993 _06072_ _06073_ _06076_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__a22o_1
X_13385_ clknet_leaf_83_clk _00704_ net200 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10597_ _04823_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08414__A2 _02468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12336_ _03689_ genblk1\[11\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR _06026_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_23_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12267_ _03707_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__buf_4
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11218_ net563 _05246_ _05250_ net822 VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__a22o_1
X_12198_ genblk2\[11\].wave_shpr.div.acc\[6\] genblk2\[11\].wave_shpr.div.b1\[6\]
+ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__or2b_1
XANTENNA__11182__B1 _04241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11149_ genblk2\[7\].wave_shpr.div.b1\[14\] genblk2\[7\].wave_shpr.div.acc\[14\]
+ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11485__A1 _03831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06690_ genblk1\[4\].osc.clkdiv_C.cnt\[0\] _01209_ _01578_ genblk1\[4\].osc.clkdiv_C.cnt\[16\]
+ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06667__A _01556_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08360_ _02885_ _02886_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__or2b_1
XFILLER_0_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07311_ genblk1\[11\].osc.clkdiv_C.cnt\[8\] _01211_ _01262_ genblk1\[11\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11788__A2 _02203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08291_ _02992_ _02996_ _02921_ _02997_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10996__B1 _05057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07242_ genblk1\[10\].osc.clkdiv_C.cnt\[0\] _01321_ _01183_ _02023_ VGND VGND VPWR
+ VPWR _02024_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07173_ genblk1\[9\].osc.clkdiv_C.cnt\[6\] _01965_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08405__A2 _01578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08106__B _01574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06124_ genblk2\[1\].wave_shpr.div.done genblk2\[0\].wave_shpr.div.done genblk2\[3\].wave_shpr.div.done
+ genblk2\[2\].wave_shpr.div.done VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__or4_2
XFILLER_0_131_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06967__A2 _01574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10652__A _02170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09366__B1 _03839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09814_ genblk2\[2\].wave_shpr.div.quo\[11\] _04253_ _04251_ net441 _04256_ VGND
+ VGND VPWR VPWR _00302_ sky130_fd_sc_hd__a221o_1
X_09745_ genblk2\[2\].wave_shpr.div.fin_quo\[5\] genblk2\[2\].wave_shpr.div.quo\[4\]
+ _00009_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06957_ genblk1\[7\].osc.clkdiv_C.cnt\[2\] _01227_ _01732_ genblk1\[7\].osc.clkdiv_C.cnt\[3\]
+ _01792_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_69_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ genblk2\[2\].wave_shpr.div.acc\[17\] _04041_ VGND VGND VPWR VPWR _04156_
+ sky130_fd_sc_hd__or2_1
X_06888_ _01658_ _01675_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__nand2_2
XFILLER_0_96_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _03293_ _03294_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__or2b_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10099__A _04269_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ genblk2\[8\].wave_shpr.div.fin_quo\[0\] genblk2\[8\].wave_shpr.div.fin_quo\[1\]
+ _02638_ _02223_ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07509_ _02228_ PWM.final_sample_in\[6\] VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__and2_1
X_08489_ _03182_ _03186_ _03195_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_135_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10520_ net763 _04657_ _04655_ _04753_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10451_ _04595_ _04702_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09054__C1 _03717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13170_ clknet_leaf_126_clk _00495_ net68 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06407__B2 _01342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10382_ genblk2\[4\].wave_shpr.div.quo\[9\] _04657_ _04655_ net251 _04658_ VGND VGND
+ VPWR VPWR _00468_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12121_ genblk2\[10\].wave_shpr.div.acc\[11\] _05878_ _05865_ VGND VGND VPWR VPWR
+ _05879_ sky130_fd_sc_hd__mux2_1
XANTENNA__07080__A1 genblk1\[8\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12052_ genblk2\[10\].wave_shpr.div.quo\[17\] _05823_ _05825_ net353 _05830_ VGND
+ VGND VPWR VPWR _00966_ sky130_fd_sc_hd__a221o_1
Xhold390 genblk2\[1\].wave_shpr.div.quo\[21\] VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ _04987_ _05090_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10911__A0 genblk2\[7\].wave_shpr.div.b1\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06591__B1 _01498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_82_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12954_ clknet_leaf_136_clk _00283_ net62 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1090 genblk2\[6\].wave_shpr.div.b1\[8\] VGND VGND VPWR VPWR net1308 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07135__A2 _01311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11905_ genblk2\[0\].wave_shpr.div.i\[3\] _02150_ _05726_ VGND VGND VPWR VPWR _05729_
+ sky130_fd_sc_hd__and3_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ clknet_leaf_30_clk _00216_ net97 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _05591_ _05678_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__xnor2_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__and2_1
X_13506_ clknet_leaf_98_clk _00823_ net167 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10718_ _04856_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07843__B1 _02527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11698_ genblk2\[9\].wave_shpr.div.b1\[9\] genblk2\[9\].wave_shpr.div.acc\[9\] VGND
+ VGND VPWR VPWR _05590_ sky130_fd_sc_hd__and2b_1
XFILLER_0_126_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07111__A genblk1\[8\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13437_ clknet_leaf_95_clk _00756_ net161 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10649_ _02171_ genblk2\[6\].wave_shpr.div.b1\[17\] VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09737__S _00009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13368_ clknet_leaf_116_clk _00687_ net139 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12319_ net342 _06014_ _06015_ net443 _06017_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__a221o_1
X_13299_ clknet_leaf_84_clk _00620_ net202 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09038__A _02336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07860_ genblk2\[1\].wave_shpr.div.fin_quo\[0\] genblk2\[1\].wave_shpr.div.fin_quo\[1\]
+ _02458_ _02459_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__nand4_1
X_06811_ genblk1\[5\].osc.clkdiv_C.cnt\[8\] _01326_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__or2_1
X_07791_ genblk1\[0\].osc.clkdiv_C.cnt\[11\] _01263_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__nand2_1
X_06742_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] _01620_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__or2_1
XANTENNA__11458__A1 _02064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09530_ _03707_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__clkbuf_2
XANTENNA__07126__A2 _01925_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09461_ _04018_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06828__C genblk1\[5\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire35 _01239_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
X_06673_ _01175_ _01194_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__or2b_1
X_08412_ _03118_ genblk2\[2\].wave_shpr.div.fin_quo\[5\] net25 VGND VGND VPWR VPWR
+ _03119_ sky130_fd_sc_hd__or3b_1
XFILLER_0_148_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09392_ genblk2\[1\].wave_shpr.div.acc\[15\] genblk2\[1\].wave_shpr.div.b1\[15\]
+ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__or2b_1
XFILLER_0_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08343_ _03013_ _03029_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout141_A net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08274_ _02979_ _02404_ _02978_ _02525_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__o31a_1
XANTENNA__07659__C _02365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07225_ _01994_ _02000_ _02004_ _02006_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07156_ genblk1\[9\].osc.clkdiv_C.cnt\[1\] genblk1\[9\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01955_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06107_ smpl_rt_clkdiv.clkDiv_inst.cnt\[5\] smpl_rt_clkdiv.clkDiv_inst.cnt\[4\] _01087_
+ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__and3_1
XANTENNA__07062__A1 genblk1\[8\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07087_ _01887_ _01897_ _01898_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_2_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout100 net101 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_2
Xfanout111 net112 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
Xfanout122 net126 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_2
Xfanout133 net135 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_4
Xfanout144 net145 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_2
Xfanout155 net157 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_4
Xfanout166 net170 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_4
Xfanout177 net180 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_4
Xfanout188 net198 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__buf_2
Xfanout199 net210 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_4
X_07989_ _02692_ _02693_ _02694_ _02695_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__a211o_1
X_09728_ _04156_ _04206_ _04207_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout54_A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09511__B1 _04047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09659_ _04009_ genblk2\[1\].wave_shpr.div.acc\[25\] genblk2\[1\].wave_shpr.div.acc\[26\]
+ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__or3b_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ clknet_leaf_90_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[1\] net173 VGND VGND
+ VPWR VPWR genblk1\[7\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _05407_ _05526_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08617__A2 _02362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07825__B1 _02223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11552_ _05473_ _05474_ net1116 _05442_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08027__A _02733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10503_ net694 _04715_ _04722_ _04742_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11483_ _05438_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13222_ clknet_leaf_114_clk net880 net132 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10434_ _04654_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07866__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10365_ _02177_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__clkbuf_4
X_13153_ clknet_leaf_121_clk net256 net77 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07053__B2 genblk1\[8\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12104_ genblk2\[10\].wave_shpr.div.acc\[7\] _05864_ _05865_ VGND VGND VPWR VPWR
+ _05866_ sky130_fd_sc_hd__mux2_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13084_ clknet_leaf_135_clk _00411_ net62 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ genblk2\[4\].wave_shpr.div.b1\[13\] genblk2\[4\].wave_shpr.div.acc\[13\]
+ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12035_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__and2_1
XANTENNA__08002__B1 _01666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08553__A1 genblk2\[6\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07817__A_N net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12937_ clknet_leaf_111_clk _00266_ net130 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_125_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10663__A2 _04853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ clknet_leaf_134_clk _00199_ net60 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11819_ _05583_ _05665_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10467__A _04651_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ clknet_leaf_59_clk net278 net192 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11997__S _05802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09018__C1 _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07010_ genblk1\[7\].osc.clkdiv_C.cnt\[9\] _01835_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07776__A _01229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08241__B1 _02527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08961_ _03649_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__clkbuf_1
X_07912_ _01233_ _02617_ _02618_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__o21ba_1
X_08892_ sig_norm.acc\[0\] _03597_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__xnor2_1
X_07843_ genblk2\[0\].wave_shpr.div.fin_quo\[2\] _02549_ _02527_ VGND VGND VPWR VPWR
+ _02550_ sky130_fd_sc_hd__o21ai_1
X_07774_ genblk1\[0\].osc.clkdiv_C.cnt\[3\] _01215_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09513_ net701 _04043_ _04047_ net755 VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__a22o_1
X_06725_ _01600_ _01610_ _01611_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11761__A _03693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09444_ genblk2\[1\].wave_shpr.div.acc\[23\] genblk2\[1\].wave_shpr.div.acc\[22\]
+ genblk2\[1\].wave_shpr.div.acc\[21\] _04007_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__or4_1
XANTENNA__10654__A2 _04853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06656_ _01523_ _01549_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__nor2_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06587_ genblk1\[3\].osc.clkdiv_C.cnt\[7\] _01494_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__xnor2_1
X_09375_ _03943_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__clkbuf_1
X_08326_ _03031_ _03032_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08257_ _02946_ _02957_ _02951_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__or3_1
XFILLER_0_105_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07208_ genblk1\[10\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__inv_2
X_08188_ _02799_ _02847_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11367__B1 _05248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07139_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01246_ _01196_ _01937_ _01938_ VGND
+ VGND VPWR VPWR _01939_ sky130_fd_sc_hd__o221a_1
XFILLER_0_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10150_ _04455_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__clkbuf_4
X_10081_ _02169_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__buf_4
XFILLER_0_100_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10342__A1 _01326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12631__RESET_B net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13771_ clknet_leaf_73_clk _01082_ net215 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10983_ _05074_ genblk1\[6\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12722_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[17\] net183 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold902_A genblk1\[5\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12653_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[2\] net89 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_1
X_11604_ _05400_ _05362_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__or2b_1
XFILLER_0_93_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12584_ clknet_leaf_124_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[5\] net76 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08471__B1 _02789_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11535_ _05464_ genblk1\[8\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07596__A net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11466_ net1268 _02433_ _05237_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13205_ clknet_leaf_8_clk _00528_ net48 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10417_ _04672_ genblk1\[4\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__and2_1
X_11397_ genblk2\[8\].wave_shpr.div.acc\[2\] genblk2\[8\].wave_shpr.div.b1\[2\] VGND
+ VGND VPWR VPWR _05373_ sky130_fd_sc_hd__or2b_1
XFILLER_0_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13136_ clknet_leaf_115_clk net465 net133 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _04641_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__clkbuf_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _04580_ _04590_ _04578_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__o21ai_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ clknet_leaf_22_clk _00394_ net93 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12018_ _02152_ genblk2\[10\].wave_shpr.div.busy _02206_ VGND VGND VPWR VPWR _05814_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10333__A1 _03714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10333__B2 _03705_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10896__S _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_139_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_139_clk sky130_fd_sc_hd__clkbuf_16
X_06510_ _01349_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07490_ _02213_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09051__A _03702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06441_ _01373_ _01380_ _01381_ VGND VGND VPWR VPWR genblk1\[1\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_8_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09160_ _03806_ VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06372_ genblk1\[1\].osc.clkdiv_C.cnt\[5\] _01305_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08111_ genblk1\[4\].osc.clkdiv_C.cnt\[14\] _01361_ _02802_ _02803_ VGND VGND VPWR
+ VPWR _02818_ sky130_fd_sc_hd__o31a_1
XFILLER_0_145_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09091_ _01201_ _03741_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08042_ genblk1\[5\].osc.clkdiv_C.cnt\[14\] _01359_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold901 genblk1\[10\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 genblk2\[6\].wave_shpr.div.i\[1\] VGND VGND VPWR VPWR net1130 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12010__A1 _03732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold923 sig_norm.acc\[11\] VGND VGND VPWR VPWR net1141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 genblk2\[3\].wave_shpr.div.b1\[13\] VGND VGND VPWR VPWR net1152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout104_A net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold945 genblk2\[11\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR net1163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 genblk2\[1\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR net1174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 genblk1\[8\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR net1185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 genblk1\[0\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR net1196 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ genblk2\[3\].wave_shpr.div.b1\[5\] genblk2\[3\].wave_shpr.div.acc\[5\] VGND
+ VGND VPWR VPWR _04389_ sky130_fd_sc_hd__and2b_1
Xhold989 genblk1\[2\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR net1207 sky130_fd_sc_hd__dlygate4sd3_1
X_08944_ sig_norm.quo\[1\] _01098_ _03635_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__a21o_1
XANTENNA__12313__A2 _03947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08875_ sig_norm.b1\[0\] _03578_ _03580_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__a21o_1
XANTENNA__09190__A1 _03706_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07826_ _02531_ _02532_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__nor2_1
XANTENNA__07740__A2 _01334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07757_ genblk2\[1\].wave_shpr.div.fin_quo\[4\] _02463_ VGND VGND VPWR VPWR _02464_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_79_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10088__B1 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06708_ _01585_ _01587_ _01590_ _01597_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__or4b_1
X_07688_ genblk1\[10\].osc.clkdiv_C.cnt\[9\] _01215_ _02011_ genblk1\[10\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09427_ _03961_ _03989_ _03990_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__a21o_1
X_06639_ genblk1\[3\].osc.clkdiv_C.cnt\[7\] _01535_ genblk1\[3\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09358_ genblk2\[0\].wave_shpr.div.acc\[21\] _03930_ _03931_ VGND VGND VPWR VPWR
+ _03932_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_75_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08309_ genblk2\[11\].wave_shpr.div.fin_quo\[4\] _02361_ VGND VGND VPWR VPWR _03016_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08453__B1 _02526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09289_ genblk2\[0\].wave_shpr.div.acc\[4\] _03879_ _03804_ VGND VGND VPWR VPWR _03880_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11320_ net808 _05311_ _05283_ _05314_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11251_ net231 _05255_ _05256_ net400 _05265_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__a221o_1
XANTENNA__08205__B1 _02316_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07559__A2 genblk1\[9\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10202_ _04408_ _04529_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__xnor2_1
X_11182_ _03732_ net389 _04241_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__o21a_1
XANTENNA__07568__A1_N genblk1\[9\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10133_ _04477_ genblk1\[3\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__and2_1
XANTENNA__12261__S _05802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12304__A2 _06009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10064_ net1232 _01589_ _04440_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__mux2_1
XANTENNA__07582__C _01221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06519__B1 _01418_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09570__S _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07731__A2 _01360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13754_ clknet_leaf_68_clk _01065_ net212 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10966_ _04676_ _01753_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__nor2_1
X_12705_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[0\] net181 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__13600__RESET_B net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06298__A2 _01256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13685_ clknet_leaf_63_clk _00998_ net191 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10897_ _05032_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12636_ clknet_leaf_19_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[3\] net109 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_72_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12567_ clknet_leaf_27_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[6\] net89 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_108_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10251__B1 _03855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11518_ net482 _05454_ _05449_ net506 _05455_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__a221o_1
X_12498_ clknet_leaf_103_clk _00060_ net156 VGND VGND VPWR VPWR sig_norm.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold208 genblk2\[1\].wave_shpr.div.quo\[18\] VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold219 _00401_ VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__dlygate4sd3_1
X_11449_ _05421_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09745__S _00009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11751__B1 _05624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ clknet_leaf_2_clk _00444_ net51 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06222__A2 _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ _01823_ _01824_ VGND VGND VPWR VPWR genblk1\[7\].osc.clkdiv_C.next_cnt\[1\]
+ sky130_fd_sc_hd__nor2_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07970__A2 _01577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11503__B1 _05446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13759__RESET_B net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08660_ _02789_ _03177_ VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__nor2_1
XANTENNA__07722__A2 _01262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07611_ _01186_ _01437_ _01225_ genblk1\[11\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR
+ VPWR _02318_ sky130_fd_sc_hd__o31a_1
X_08591_ _03246_ _03258_ _03296_ _03297_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__a211o_2
X_07542_ _02254_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07473_ genblk2\[9\].wave_shpr.div.i\[1\] _02200_ genblk2\[9\].wave_shpr.div.i\[4\]
+ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__or3b_1
XFILLER_0_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09212_ _03834_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06424_ _01365_ _01367_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09227__A2 _03836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09143_ genblk2\[0\].wave_shpr.div.b1\[14\] genblk2\[0\].wave_shpr.div.acc\[14\]
+ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__and2b_1
X_06355_ genblk1\[0\].osc.clkdiv_C.cnt\[17\] _01298_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09074_ genblk2\[0\].wave_shpr.div.b1\[13\] _01592_ _03722_ VGND VGND VPWR VPWR _03730_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06286_ _01247_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__buf_4
X_08025_ genblk1\[6\].osc.clkdiv_C.cnt\[16\] genblk1\[6\].osc.clkdiv_C.cnt\[17\] VGND
+ VGND VPWR VPWR _02732_ sky130_fd_sc_hd__nor2_1
Xhold720 genblk2\[9\].wave_shpr.div.acc\[6\] VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 genblk2\[11\].wave_shpr.div.acc\[13\] VGND VGND VPWR VPWR net949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold742 genblk2\[11\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR net960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 genblk2\[4\].wave_shpr.div.acc\[7\] VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 genblk2\[5\].wave_shpr.div.acc\[20\] VGND VGND VPWR VPWR net982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 genblk2\[11\].wave_shpr.div.acc\[14\] VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 genblk2\[0\].wave_shpr.div.acc\[11\] VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 genblk2\[6\].wave_shpr.div.acc\[3\] VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10390__A _04654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09976_ genblk2\[3\].wave_shpr.div.acc\[6\] genblk2\[3\].wave_shpr.div.b1\[6\] VGND
+ VGND VPWR VPWR _04372_ sky130_fd_sc_hd__or2b_1
X_08927_ _01099_ _01156_ _03623_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__and3_1
X_08858_ _03559_ _03563_ _03564_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07809_ _02514_ _02515_ genblk2\[0\].wave_shpr.div.fin_quo\[6\] _02468_ VGND VGND
+ VPWR VPWR _02516_ sky130_fd_sc_hd__a2bb2o_1
X_08789_ _03491_ _03495_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__xnor2_1
X_10820_ net855 _02181_ _04962_ _03708_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__a31o_1
XANTENNA__07204__A genblk1\[9\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10751_ _04802_ _04769_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__or2b_1
XANTENNA__11273__A2 _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13470_ clknet_leaf_74_clk _00787_ net203 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10682_ _04672_ genblk1\[5\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__and2_1
XANTENNA__09218__A2 _03836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12421_ genblk2\[11\].wave_shpr.div.acc\[25\] genblk2\[11\].wave_shpr.div.acc\[24\]
+ genblk2\[11\].wave_shpr.div.acc\[26\] _05980_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__nor4_1
XFILLER_0_118_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12352_ _03944_ _06033_ _06035_ _03947_ net1127 VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__a32o_1
XANTENNA__08035__A _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11303_ net916 _05279_ _05283_ _05301_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__a22o_1
X_12283_ genblk2\[1\].wave_shpr.div.b1\[10\] _01946_ _05994_ VGND VGND VPWR VPWR _06003_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08729__B2 _02468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09565__S _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11234_ _05249_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__buf_2
XFILLER_0_31_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12930__D _00009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11165_ genblk2\[7\].wave_shpr.div.fin_quo\[1\] net1347 _00019_ VGND VGND VPWR VPWR
+ _05224_ sky130_fd_sc_hd__mux2_1
XANTENNA__07952__A2 _01801_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10116_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__and2_1
X_11096_ genblk2\[6\].wave_shpr.div.i\[1\] genblk2\[6\].wave_shpr.div.i\[0\] genblk2\[6\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10047_ _03727_ _04432_ net1075 _03687_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__a2bb2o_1
Xhold80 genblk2\[0\].wave_shpr.div.quo\[19\] VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 _00551_ VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12020__A _05815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11998_ _05804_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07114__A genblk1\[8\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13737_ clknet_leaf_47_clk _01048_ net119 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10949_ _04869_ genblk1\[6\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_70_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_900 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13668_ clknet_leaf_42_clk _00981_ net123 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_144_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12619_ clknet_leaf_17_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[4\] net83 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__06691__A2 _01210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13599_ clknet_leaf_77_clk _00914_ net208 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06140_ _01103_ _01111_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06979__B1 _01196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07928__C1 genblk1\[8\].osc.clkdiv_C.cnt\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08196__A2 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09830_ net339 _04257_ _04259_ net393 _04265_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__a221o_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07943__A2 _01925_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _01436_ _04229_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__nand2_4
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01363_ _01311_ genblk1\[7\].osc.clkdiv_C.cnt\[11\]
+ _01808_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__a221o_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _03406_ _03407_ _03359_ _03381_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__a211o_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ genblk2\[2\].wave_shpr.div.b1\[1\] genblk2\[2\].wave_shpr.div.acc\[1\] VGND
+ VGND VPWR VPWR _04172_ sky130_fd_sc_hd__or2b_1
X_08643_ _02604_ _03344_ _03348_ _02648_ VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout171_A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08574_ genblk2\[11\].wave_shpr.div.fin_quo\[0\] net33 _02350_ genblk2\[11\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07525_ _02243_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08656__B1 _02885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_61_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08120__A2 _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07456_ _02186_ _02153_ genblk2\[6\].wave_shpr.div.busy VGND VGND VPWR VPWR _02189_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06407_ genblk1\[1\].osc.clkdiv_C.cnt\[16\] _01349_ _01350_ _01342_ VGND VGND VPWR
+ VPWR _01351_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06682__A2 _01439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10385__A _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07387_ _02137_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[13\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09126_ _03758_ _03772_ _03773_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__a21o_1
X_06338_ genblk1\[0\].osc.clkdiv_C.cnt\[10\] _01286_ genblk1\[0\].osc.clkdiv_C.cnt\[11\]
+ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12475__RESET_B net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06269_ _01229_ _01230_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__nor2_4
XFILLER_0_103_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09057_ _03718_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08008_ genblk1\[6\].osc.clkdiv_C.cnt\[3\] _01730_ _01758_ _01729_ VGND VGND VPWR
+ VPWR _02715_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_103_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold550 genblk2\[8\].wave_shpr.div.b1\[7\] VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 genblk2\[3\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 genblk2\[3\].wave_shpr.div.acc\[10\] VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 genblk2\[7\].wave_shpr.div.i\[2\] VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09384__A1 _03944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold594 genblk2\[2\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11191__A1 _01556_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout84_A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09959_ _04251_ _04355_ _04357_ _04253_ net711 VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__a32o_1
X_12970_ clknet_leaf_113_clk net276 net128 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11921_ genblk2\[10\].wave_shpr.div.acc\[4\] genblk2\[10\].wave_shpr.div.b1\[4\]
+ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__and2b_1
XANTENNA__13263__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07860__C _02458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ net799 _05684_ _05685_ _05691_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__a22o_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _04952_ _04949_ _04953_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11783_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_52_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08111__A2 _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13522_ clknet_leaf_79_clk _00839_ net206 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_138_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10734_ _04794_ _04773_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__or2b_1
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07870__A1 _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13453_ clknet_leaf_99_clk _00770_ net168 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_24_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10665_ _02182_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06492__B _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12404_ genblk2\[11\].wave_shpr.div.acc\[13\] _06075_ _06055_ VGND VGND VPWR VPWR
+ _06076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13384_ clknet_leaf_83_clk _00703_ net200 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10596_ genblk2\[5\].wave_shpr.div.fin_quo\[1\] genblk2\[5\].wave_shpr.div.quo\[0\]
+ _00015_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12335_ genblk2\[11\].wave_shpr.div.quo\[21\] _06014_ _06015_ net239 _06025_ VGND
+ VGND VPWR VPWR _01054_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12266_ _05993_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__clkbuf_1
X_11217_ _05249_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12197_ genblk2\[11\].wave_shpr.div.acc\[7\] genblk2\[11\].wave_shpr.div.b1\[7\]
+ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__or2b_1
XANTENNA__11182__A1 _03732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11148_ _05168_ _05206_ _05207_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__a21o_1
X_11079_ genblk2\[6\].wave_shpr.div.acc\[22\] _05146_ VGND VGND VPWR VPWR _05148_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__07138__B1 genblk1\[9\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06667__B _01344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_43_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_16
X_07310_ genblk1\[11\].osc.clkdiv_C.cnt\[10\] _02002_ VGND VGND VPWR VPWR _02074_
+ sky130_fd_sc_hd__xnor2_1
X_08290_ _02747_ _02919_ _02920_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__a21o_1
XANTENNA__09850__A2 _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10996__A1 _05055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07241_ genblk1\[10\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07172_ _01953_ _01965_ _01966_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_82_891 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06123_ genblk2\[5\].wave_shpr.div.done genblk2\[4\].wave_shpr.div.done genblk2\[7\].wave_shpr.div.done
+ genblk2\[6\].wave_shpr.div.done VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__or4_4
XFILLER_0_14_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13774__RESET_B net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09813_ _04058_ _01414_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__nor2_1
XANTENNA__10920__A1 _02433_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11764__A _02155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09744_ _04219_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07961__B _01360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06956_ genblk1\[7\].osc.clkdiv_C.cnt\[11\] _01311_ _01732_ genblk1\[7\].osc.clkdiv_C.cnt\[3\]
+ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__o22ai_1
X_09675_ net285 _04154_ _04155_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__a21oi_1
X_06887_ genblk1\[6\].osc.clkdiv_C.cnt\[1\] _01738_ _01740_ VGND VGND VPWR VPWR _01741_
+ sky130_fd_sc_hd__a21bo_1
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _03331_ _03332_ _03298_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__nand3b_2
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ genblk2\[8\].wave_shpr.div.fin_quo\[0\] _02638_ genblk2\[8\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_34_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07508_ PWM.counter\[6\] VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08488_ _03187_ _03194_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07439_ _02147_ _02176_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10450_ _04596_ _04575_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__or2b_1
XFILLER_0_17_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09109_ genblk2\[0\].wave_shpr.div.acc\[6\] genblk2\[0\].wave_shpr.div.b1\[6\] VGND
+ VGND VPWR VPWR _03757_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10381_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12120_ _05767_ _05877_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12051_ _03833_ _02003_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold380 genblk2\[0\].wave_shpr.div.quo\[9\] VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 genblk2\[6\].wave_shpr.div.quo\[22\] VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11002_ _04988_ _04980_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__or2b_1
XANTENNA__10911__A1 _04444_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12953_ clknet_leaf_136_clk _00282_ net62 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1080 genblk2\[3\].wave_shpr.div.b1\[8\] VGND VGND VPWR VPWR net1298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1091 genblk2\[4\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net1309 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ _00000_ _05726_ net1158 VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__a21oi_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12884_ clknet_leaf_30_clk net461 net97 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11219__A2 _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11835_ _05592_ _05561_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__or2b_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07599__A _02261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ genblk2\[9\].wave_shpr.div.quo\[13\] _05628_ _05629_ net243 _05632_ VGND
+ VGND VPWR VPWR _00878_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ clknet_leaf_98_clk _00822_ net167 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10717_ net961 _04886_ _04857_ _04889_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__a22o_1
X_11697_ _05563_ _05587_ _05588_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__a21o_1
X_13436_ clknet_leaf_95_clk _00755_ net159 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07111__B genblk1\[8\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10648_ _03726_ _04851_ _03736_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13367_ clknet_leaf_116_clk _00686_ net139 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_106_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10579_ _04767_ _04805_ _04806_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__a21o_1
X_12318_ _05835_ genblk1\[11\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__and2_1
X_13298_ clknet_leaf_84_clk _00619_ net202 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12249_ genblk2\[11\].wave_shpr.div.fin_quo\[2\] net769 _00005_ VGND VGND VPWR VPWR
+ _05985_ sky130_fd_sc_hd__mux2_1
XANTENNA__09038__B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12352__B1 _03947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10902__A1 _01923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06810_ genblk1\[5\].osc.clkdiv_C.cnt\[8\] _01326_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__nand2_1
X_07790_ genblk1\[0\].osc.clkdiv_C.cnt\[10\] _01996_ _01801_ VGND VGND VPWR VPWR _02497_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06741_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] _01620_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__nand2_1
Xwire25 _03112_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
X_09460_ genblk2\[1\].wave_shpr.div.fin_quo\[6\] genblk2\[1\].wave_shpr.div.quo\[5\]
+ _00007_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__mux2_1
X_06672_ genblk1\[4\].osc.clkdiv_C.cnt\[3\] _01326_ _01498_ genblk1\[4\].osc.clkdiv_C.cnt\[14\]
+ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08893__A _01099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08411_ genblk2\[2\].wave_shpr.div.fin_quo\[4\] _03117_ VGND VGND VPWR VPWR _03118_
+ sky130_fd_sc_hd__or2_1
X_09391_ genblk2\[1\].wave_shpr.div.acc\[16\] genblk2\[1\].wave_shpr.div.b1\[16\]
+ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_16_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__10418__B1 _04654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08342_ _03041_ _03042_ _03047_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08273_ _02404_ _02978_ _02979_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08117__B _01326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07224_ genblk1\[10\].osc.clkdiv_C.cnt\[11\] _02005_ VGND VGND VPWR VPWR _02006_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07155_ _01952_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06106_ smpl_rt_clkdiv.clkDiv_inst.cnt\[3\] _01086_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__and2_1
XANTENNA__07062__A2 _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07086_ genblk1\[8\].osc.clkdiv_C.cnt\[6\] _01895_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout101 net107 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12343__B1 _03941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout112 net127 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_2
Xfanout123 net125 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_4
Xfanout134 net135 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_4
Xfanout145 net171 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_4
Xfanout156 net157 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_4
Xfanout167 net170 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10602__S _00015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout178 net180 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_2
Xfanout189 net191 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_4
X_07988_ _02217_ _02553_ genblk2\[7\].wave_shpr.div.fin_quo\[7\] VGND VGND VPWR VPWR
+ _02695_ sky130_fd_sc_hd__and3_1
XANTENNA__06588__A _01437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09727_ genblk2\[2\].wave_shpr.div.acc\[17\] _04041_ VGND VGND VPWR VPWR _04207_
+ sky130_fd_sc_hd__and2_1
X_06939_ genblk1\[6\].osc.clkdiv_C.cnt\[12\] genblk1\[6\].osc.clkdiv_C.cnt\[11\] _01777_
+ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10657__B1 _04857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09511__B2 net764 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09658_ net1228 _04048_ _04045_ _04144_ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__a22o_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout47_A net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08609_ _03314_ _02789_ _03315_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _03984_ _03964_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__or2b_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _05408_ _05358_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12490__RESET_B net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09814__A2 _04253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11551_ genblk2\[8\].wave_shpr.div.b1\[0\] genblk2\[8\].wave_shpr.div.acc\[0\] _05417_
+ _05471_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10502_ _04740_ _04741_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11482_ genblk2\[9\].wave_shpr.div.b1\[12\] _02656_ _05433_ VGND VGND VPWR VPWR _05438_
+ sky130_fd_sc_hd__mux2_1
X_13221_ clknet_leaf_114_clk _00544_ net132 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10433_ net1068 _04683_ _04656_ _04689_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13152_ clknet_leaf_17_clk _00477_ net80 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10364_ _04650_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12103_ _05786_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ clknet_leaf_135_clk _00410_ net61 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10295_ _04570_ _04605_ _04606_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__a21o_1
X_12034_ net432 _05818_ _05816_ genblk2\[10\].wave_shpr.div.quo\[8\] _05820_ VGND
+ VGND VPWR VPWR _00958_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08553__A2 genblk2\[6\].wave_shpr.div.fin_quo\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10648__B1 _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12936_ clknet_leaf_113_clk _00265_ net130 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_87_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12867_ clknet_leaf_134_clk _00198_ net60 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11818_ _05584_ _05565_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__or2b_1
XFILLER_0_56_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09266__B1 _03838_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ clknet_leaf_57_clk _00131_ net183 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09805__A2 _04248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11749_ net586 _05623_ _05624_ net700 VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10820__B1 _03708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06961__A _01432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13419_ clknet_leaf_91_clk _00738_ net147 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07776__B _01359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11376__A1 _05248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08960_ sig_norm.quo\[5\] _03648_ _00024_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_5_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_16
X_07911_ _01228_ _01308_ _01440_ _01889_ _01879_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__o41a_1
X_08891_ sig_norm.b1\[0\] _03596_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__nand2_1
X_07842_ genblk2\[0\].wave_shpr.div.fin_quo\[0\] genblk2\[0\].wave_shpr.div.fin_quo\[1\]
+ _02510_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__o21a_1
XANTENNA__11422__A_N genblk2\[8\].wave_shpr.div.b1\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07773_ genblk1\[0\].osc.clkdiv_C.cnt\[2\] _01556_ _01564_ _01190_ genblk1\[0\].osc.clkdiv_C.cnt\[1\]
+ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09512_ genblk2\[1\].wave_shpr.div.quo\[2\] _04043_ _04047_ net684 VGND VGND VPWR
+ VPWR _00209_ sky130_fd_sc_hd__a22o_1
X_06724_ genblk1\[4\].osc.clkdiv_C.cnt\[3\] _01605_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__or2_1
XANTENNA__12930__RESET_B net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09443_ genblk2\[1\].wave_shpr.div.acc\[20\] genblk2\[1\].wave_shpr.div.acc\[19\]
+ _04006_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__or3_1
X_06655_ genblk1\[3\].osc.clkdiv_C.cnt\[14\] _01547_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09374_ _03941_ _03942_ genblk2\[11\].wave_shpr.div.i\[0\] VGND VGND VPWR VPWR _03943_
+ sky130_fd_sc_hd__mux2_1
X_06586_ _01342_ _01248_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__nor2_4
XFILLER_0_47_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08325_ genblk2\[8\].wave_shpr.div.fin_quo\[4\] _02638_ _02640_ _02223_ VGND VGND
+ VPWR VPWR _03032_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10811__B1 _04858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08256_ _02742_ _02962_ _02745_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07207_ net1194 _01988_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__11489__A _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08187_ _02890_ _02891_ _02892_ _02893_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__a31o_1
XANTENNA__10393__A _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07138_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01246_ genblk1\[9\].osc.clkdiv_C.cnt\[17\]
+ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07069_ _01886_ VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__clkbuf_4
X_10080_ _04450_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13770_ clknet_leaf_71_clk _01081_ net215 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10982_ net385 _05051_ _05054_ net609 _05076_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12721_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[16\] net183 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_97_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12652_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[1\] net89 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08038__A net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11603_ net833 _05507_ _05484_ _05513_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__a22o_1
X_12583_ clknet_leaf_124_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[4\] net72 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11534_ _04268_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11465_ _05429_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_49_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13204_ clknet_leaf_8_clk _00527_ net48 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10416_ net714 _04651_ _04654_ net698 _04677_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11396_ genblk2\[8\].wave_shpr.div.acc\[3\] genblk2\[8\].wave_shpr.div.b1\[3\] VGND
+ VGND VPWR VPWR _05372_ sky130_fd_sc_hd__or2b_1
X_13135_ clknet_leaf_114_clk net419 net133 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10347_ net1283 _01658_ _04637_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12307__B1 _06010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ clknet_leaf_22_clk net452 net93 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10278_ _04581_ _04588_ _04589_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__a21oi_1
X_12017_ _05812_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_cap1 _05138_ VGND VGND VPWR VPWR net1350 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11294__B1 _05283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12919_ clknet_leaf_39_clk _00250_ net115 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06675__B _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06440_ genblk1\[1\].osc.clkdiv_C.cnt\[3\] _01378_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06371_ _01307_ _01311_ _01312_ genblk1\[1\].osc.clkdiv_C.cnt\[11\] _01314_ VGND
+ VGND VPWR VPWR _01315_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08110_ genblk1\[4\].osc.clkdiv_C.cnt\[10\] _01313_ _02809_ _02810_ _02816_ VGND
+ VGND VPWR VPWR _02817_ sky130_fd_sc_hd__o311a_1
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13547__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09090_ _03739_ _03740_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08041_ genblk1\[5\].osc.clkdiv_C.cnt\[15\] _01576_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold902 genblk1\[5\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 sig_norm.acc\[0\] VGND VGND VPWR VPWR net1131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold924 PWM.final_sample_in\[7\] VGND VGND VPWR VPWR net1142 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_6_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold935 genblk2\[10\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR net1153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold946 genblk2\[8\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR net1164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 genblk2\[0\].wave_shpr.div.acc\[20\] VGND VGND VPWR VPWR net1175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 genblk2\[4\].wave_shpr.div.b1\[9\] VGND VGND VPWR VPWR net1186 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ _04376_ _04387_ _04374_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__o21ai_1
Xhold979 genblk2\[2\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net1197 sky130_fd_sc_hd__dlygate4sd3_1
X_08943_ _03545_ _03634_ _03546_ _01155_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__o211a_1
XANTENNA__11756__B genblk1\[9\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
X_08874_ _03577_ _03579_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07725__B1 _01313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07825_ genblk2\[0\].wave_shpr.div.fin_quo\[3\] _02510_ _02511_ _02223_ VGND VGND
+ VPWR VPWR _02532_ sky130_fd_sc_hd__a31o_1
X_07756_ genblk2\[1\].wave_shpr.div.fin_quo\[2\] genblk2\[1\].wave_shpr.div.fin_quo\[3\]
+ _02462_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__or3_1
XANTENNA__10088__B2 net794 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06707_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] _01304_ _01593_ _01594_ _01596_ VGND VGND
+ VPWR VPWR _01597_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_79_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10388__A _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07687_ genblk1\[10\].osc.clkdiv_C.cnt\[11\] _02011_ _02005_ genblk1\[10\].osc.clkdiv_C.cnt\[10\]
+ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__o22ai_2
X_09426_ genblk2\[1\].wave_shpr.div.b1\[10\] genblk2\[1\].wave_shpr.div.acc\[10\]
+ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__and2b_1
X_06638_ genblk1\[3\].osc.clkdiv_C.cnt\[8\] genblk1\[3\].osc.clkdiv_C.cnt\[7\] _01535_
+ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09357_ genblk2\[0\].wave_shpr.div.acc\[21\] genblk2\[0\].wave_shpr.div.acc\[20\]
+ _03800_ net1352 VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__or4_1
XFILLER_0_136_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06569_ net1167 _01476_ _01479_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07697__A _02403_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08308_ genblk2\[11\].wave_shpr.div.fin_quo\[3\] _02349_ _02351_ _02353_ _02222_
+ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__a41o_1
XFILLER_0_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09288_ _03878_ _03770_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06464__B1 genblk1\[1\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08239_ _02646_ _02647_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11250_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10201_ _04409_ _04363_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__or2b_1
X_11181_ _03819_ _01242_ _02064_ _05231_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__o31a_1
XFILLER_0_31_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10132_ _04268_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__buf_2
XFILLER_0_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10063_ _04441_ VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10062__S _04440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07731__A3 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13753_ clknet_leaf_68_clk _01064_ net211 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10965_ net594 _05062_ _05064_ net498 _05067_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__a221o_1
X_12704_ clknet_leaf_89_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[17\] net173 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_1
X_13684_ clknet_leaf_63_clk _00997_ net191 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10896_ genblk2\[7\].wave_shpr.div.b1\[0\] _01514_ _04848_ VGND VGND VPWR VPWR _05032_
+ sky130_fd_sc_hd__mux2_1
X_12635_ clknet_leaf_16_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[2\] net74 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12566_ clknet_leaf_28_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[5\] net89 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07400__A net1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11517_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__and2_1
X_12497_ clknet_leaf_102_clk _00059_ net156 VGND VGND VPWR VPWR sig_norm.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12018__A _02152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold209 _00225_ VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ genblk2\[8\].wave_shpr.div.fin_quo\[3\] net1337 _00021_ VGND VGND VPWR VPWR
+ _05421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11379_ _03690_ _05355_ _05356_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__nor3_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ clknet_leaf_125_clk _00443_ net69 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ clknet_leaf_112_clk _00376_ net132 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08380__B1 _02425_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07610_ genblk1\[11\].osc.clkdiv_C.cnt\[7\] _01211_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__nand2_1
X_08590_ _03275_ _03276_ _03295_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09062__A _03701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07541_ PWM.final_sample_in\[2\] net1102 PWM.start VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07472_ genblk2\[9\].wave_shpr.div.i\[2\] genblk2\[9\].wave_shpr.div.i\[3\] genblk2\[9\].wave_shpr.div.i\[0\]
+ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__nand3b_1
XANTENNA__08683__B2 _02468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09211_ _03833_ net1302 VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06423_ _01366_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__clkbuf_4
X_09142_ _03750_ _03788_ _03789_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08435__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06354_ net1196 _01296_ _01299_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[16\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07238__A2 _02011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06254__A1_N genblk1\[0\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08406__A net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10703__B_N _04856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09073_ _03729_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06285_ _01173_ _01191_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout214_A net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11990__A1 _04230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08024_ _02711_ _02724_ _02727_ _02730_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__a31o_1
Xhold710 genblk2\[4\].wave_shpr.div.acc\[9\] VGND VGND VPWR VPWR net928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold721 sig_norm.i\[0\] VGND VGND VPWR VPWR net939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 genblk2\[8\].wave_shpr.div.acc\[7\] VGND VGND VPWR VPWR net950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 genblk2\[5\].wave_shpr.div.acc\[3\] VGND VGND VPWR VPWR net961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold754 _00492_ VGND VGND VPWR VPWR net972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 genblk2\[1\].wave_shpr.div.acc\[19\] VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold776 _01073_ VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11742__A1 _02248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold787 genblk2\[8\].wave_shpr.div.b1\[13\] VGND VGND VPWR VPWR net1005 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ genblk2\[3\].wave_shpr.div.acc\[7\] genblk2\[3\].wave_shpr.div.b1\[7\] VGND
+ VGND VPWR VPWR _04371_ sky130_fd_sc_hd__or2b_1
Xhold798 genblk2\[3\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR net1016 sky130_fd_sc_hd__dlygate4sd3_1
X_08926_ sig_norm.acc\[9\] _03589_ _03622_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__a21o_1
X_08857_ _03562_ _03557_ _03560_ _03561_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07808_ genblk2\[0\].wave_shpr.div.fin_quo\[5\] _02510_ _02513_ _02224_ VGND VGND
+ VPWR VPWR _02515_ sky130_fd_sc_hd__a31o_1
XANTENNA__10610__S _04637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08788_ _03114_ _03494_ _03122_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__o21a_1
X_07739_ genblk1\[1\].osc.clkdiv_C.cnt\[9\] _01334_ _01312_ genblk1\[1\].osc.clkdiv_C.cnt\[10\]
+ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08123__B1 _01565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10750_ net1061 _04886_ _04890_ _04914_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09409_ _03970_ _03971_ _03972_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__a21o_1
X_10681_ genblk2\[5\].wave_shpr.div.quo\[15\] _04861_ _04862_ net249 _04867_ VGND
+ VGND VPWR VPWR _00558_ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12420_ net576 _06072_ _06073_ _06087_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07220__A _01365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12351_ _05982_ _06034_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10057__S _04238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08035__B _02733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11302_ genblk2\[7\].wave_shpr.div.acc\[8\] _05299_ _05300_ VGND VGND VPWR VPWR _05301_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12282_ _06002_ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11233_ _05245_ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__buf_2
X_11164_ _05223_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__clkbuf_1
X_10115_ net376 _04461_ _04462_ net514 _04468_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__a221o_1
X_11095_ genblk2\[6\].wave_shpr.div.i\[1\] genblk2\[6\].wave_shpr.div.i\[0\] genblk2\[6\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__a21o_1
X_10046_ _01325_ _01996_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__nor2_2
XFILLER_0_117_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold70 genblk2\[11\].wave_shpr.div.i\[4\] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 _00143_ VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 genblk2\[5\].wave_shpr.div.quo\[9\] VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11997_ net1275 _01556_ _05802_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10948_ _05051_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__clkbuf_4
X_13736_ clknet_leaf_47_clk net343 net119 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09610__A _04042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13667_ clknet_leaf_42_clk _00980_ net124 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10879_ _05022_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__buf_4
XFILLER_0_85_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12618_ clknet_leaf_17_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[3\] net80 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
X_13598_ clknet_leaf_76_clk net647 net208 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_775 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12549_ clknet_leaf_60_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[6\] net186 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 _04242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08196__A3 _02350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _01325_ _01423_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__nor2_4
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06972_ genblk1\[7\].osc.clkdiv_C.cnt\[13\] _01214_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__xnor2_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _03410_ _03417_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__xor2_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11488__B1 _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09691_ genblk2\[2\].wave_shpr.div.b1\[2\] VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__inv_2
X_08642_ _02604_ _02648_ _03344_ _03348_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__nand4_1
XFILLER_0_89_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08573_ _02310_ _03279_ _02314_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07524_ _01152_ sig_norm.i\[0\] sig_norm.busy VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__and3b_1
XFILLER_0_49_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09520__A _03855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07455_ _02188_ VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__inv_2
XANTENNA__11660__B1 _03855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10666__A _04672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06406_ _01201_ genblk1\[1\].osc.clkdiv_C.cnt\[13\] genblk1\[1\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07386_ _02091_ _02135_ _02136_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07040__A _01489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09125_ genblk2\[0\].wave_shpr.div.b1\[5\] genblk2\[0\].wave_shpr.div.acc\[5\] VGND
+ VGND VPWR VPWR _03773_ sky130_fd_sc_hd__and2b_1
X_06337_ genblk1\[0\].osc.clkdiv_C.cnt\[10\] _01286_ _01288_ _01270_ VGND VGND VPWR
+ VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o211a_1
XFILLER_0_127_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09081__A1 _03704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09056_ net1289 _01201_ _03708_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__mux2_1
X_06268_ _01220_ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11497__A _05444_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08007_ _01729_ _01758_ _01735_ genblk1\[6\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR
+ VPWR _02714_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_103_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold540 genblk2\[7\].wave_shpr.div.b1\[16\] VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__dlygate4sd3_1
X_06199_ PWM.counter\[5\] PWM.counter\[4\] _01161_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__and3_1
Xhold551 genblk2\[11\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10518__A2 _04657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07919__B1 _01858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold562 _00379_ VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 genblk2\[3\].wave_shpr.div.acc\[11\] VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 genblk2\[8\].wave_shpr.div.acc\[16\] VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 genblk2\[1\].wave_shpr.div.acc\[10\] VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08592__B1 _02521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09958_ _04356_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout77_A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08909_ _03587_ net26 VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__or2_1
X_09889_ _04190_ _04306_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__xnor2_1
X_11920_ genblk2\[10\].wave_shpr.div.acc\[5\] genblk2\[10\].wave_shpr.div.b1\[5\]
+ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07860__D _02459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ genblk2\[9\].wave_shpr.div.acc\[13\] _05690_ _05673_ VGND VGND VPWR VPWR
+ _05691_ sky130_fd_sc_hd__mux2_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ genblk2\[5\].wave_shpr.div.acc\[24\] _04880_ _04949_ VGND VGND VPWR VPWR
+ _04953_ sky130_fd_sc_hd__or3b_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11782_ net416 _05628_ _05629_ net533 _05640_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__a221o_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09844__B1 _04250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10733_ net1037 _04886_ _04890_ _04901_ VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__a22o_1
X_13521_ clknet_leaf_79_clk _00838_ net206 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13452_ clknet_leaf_99_clk _00769_ net166 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_10664_ genblk2\[5\].wave_shpr.div.quo\[8\] _04853_ _04857_ net308 VGND VGND VPWR
+ VPWR _00551_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_14_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12403_ _05966_ _06074_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09072__A1 _01340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13383_ clknet_leaf_83_clk _00702_ net200 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10595_ _04822_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07885__A _02526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07083__B1 genblk1\[8\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12334_ _03689_ genblk1\[11\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR _06025_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_50_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12265_ net1295 _01240_ _05802_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__mux2_1
XANTENNA__10509__A2 _04657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11216_ _05247_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__clkbuf_4
X_12196_ genblk2\[11\].wave_shpr.div.acc\[8\] genblk2\[11\].wave_shpr.div.b1\[8\]
+ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__or2b_1
X_11147_ genblk2\[7\].wave_shpr.div.b1\[13\] genblk2\[7\].wave_shpr.div.acc\[13\]
+ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11078_ net1031 _05119_ _05126_ _05147_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__a22o_1
XANTENNA__07138__A1 genblk1\[9\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10029_ genblk2\[3\].wave_shpr.div.fin_quo\[1\] genblk2\[3\].wave_shpr.div.quo\[0\]
+ _04422_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13719_ clknet_leaf_36_clk _01030_ net105 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11185__A1_N _03727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07240_ genblk1\[10\].osc.clkdiv_C.cnt\[3\] _02013_ _02021_ VGND VGND VPWR VPWR _02022_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__07861__A2 _02458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07171_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01960_ genblk1\[9\].osc.clkdiv_C.cnt\[5\]
+ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07304__A2_N _02064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06122_ genblk2\[9\].wave_shpr.div.done genblk2\[8\].wave_shpr.div.done genblk2\[11\].wave_shpr.div.done
+ genblk2\[10\].wave_shpr.div.done VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__or4_2
XFILLER_0_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09366__A2 _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09812_ net441 _04253_ _04251_ net574 _04255_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__a221o_1
X_09743_ genblk2\[2\].wave_shpr.div.fin_quo\[4\] net1327 _00009_ VGND VGND VPWR VPWR
+ _04219_ sky130_fd_sc_hd__mux2_1
X_06955_ net1063 _01790_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10160__S _04420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09674_ net285 _04154_ _03819_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__o21ai_1
X_06886_ genblk1\[6\].osc.clkdiv_C.cnt\[1\] _01738_ _01739_ genblk1\[6\].osc.clkdiv_C.cnt\[8\]
+ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__o22a_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _03296_ _03297_ _03246_ _03258_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__o211ai_2
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _02742_ _03261_ _03262_ _02745_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__o31a_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07507_ PWM.counter\[7\] VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__inv_2
XANTENNA__09250__A _03853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12087__S _05787_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08487_ _02939_ _03193_ _02943_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07438_ genblk2\[4\].wave_shpr.div.busy _02175_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07852__A2 _02309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07369_ _02123_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__inv_2
XANTENNA__09054__A1 _03714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09108_ genblk2\[0\].wave_shpr.div.acc\[7\] genblk2\[0\].wave_shpr.div.b1\[7\] VGND
+ VGND VPWR VPWR _03756_ sky130_fd_sc_hd__or2b_1
XANTENNA__07604__A2 _02309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10380_ _04651_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12625__RESET_B net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09039_ _02147_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12050_ net353 _05823_ _05825_ net357 _05829_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__a221o_1
Xhold370 genblk2\[1\].wave_shpr.div.acc_next\[0\] VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 genblk2\[0\].wave_shpr.div.quo\[11\] VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ net1015 _05086_ _05056_ _05089_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__a22o_1
Xhold392 genblk2\[1\].wave_shpr.div.quo\[10\] VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__dlygate4sd3_1
X_12952_ clknet_leaf_125_clk _00281_ net61 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1070 genblk2\[7\].wave_shpr.div.b1\[2\] VGND VGND VPWR VPWR net1288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 genblk2\[1\].wave_shpr.div.b1\[13\] VGND VGND VPWR VPWR net1299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1092 genblk2\[11\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net1310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06879__B1 _01732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11903_ _03839_ _05725_ _05727_ _03841_ net775 VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__a32o_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ clknet_leaf_55_clk net293 net176 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ net884 _05652_ _05653_ _05677_ VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__a22o_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09817__B1 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ genblk2\[5\].wave_shpr.div.acc\[2\] _04888_ _04821_ VGND VGND VPWR VPWR _04889_
+ sky130_fd_sc_hd__mux2_1
X_13504_ clknet_leaf_81_clk _00821_ net199 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11696_ genblk2\[9\].wave_shpr.div.b1\[8\] genblk2\[9\].wave_shpr.div.acc\[8\] VGND
+ VGND VPWR VPWR _05588_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10647_ net1096 VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__inv_2
X_13435_ clknet_leaf_95_clk _00754_ net161 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09045__A1 _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13366_ clknet_leaf_91_clk _00685_ net143 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_10578_ genblk2\[5\].wave_shpr.div.b1\[13\] genblk2\[5\].wave_shpr.div.acc\[13\]
+ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12317_ net443 _06014_ _06015_ genblk2\[11\].wave_shpr.div.quo\[11\] _06016_ VGND
+ VGND VPWR VPWR _01045_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13297_ clknet_leaf_86_clk _00618_ net179 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12248_ _05984_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12352__A1 _03944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12179_ genblk2\[10\].wave_shpr.div.i\[1\] genblk2\[10\].wave_shpr.div.i\[0\] genblk2\[10\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08308__B1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06740_ _01623_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06671_ genblk1\[4\].osc.clkdiv_C.cnt\[2\] _01559_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__nor2_1
X_08410_ genblk2\[2\].wave_shpr.div.fin_quo\[3\] _03116_ VGND VGND VPWR VPWR _03117_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09390_ genblk2\[1\].wave_shpr.div.acc\[17\] genblk2\[1\].wave_shpr.div.b1\[17\]
+ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09070__A _03702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08341_ _03041_ _03042_ _03047_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__nand3_1
XFILLER_0_86_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08272_ genblk2\[10\].wave_shpr.div.fin_quo\[4\] VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07223_ _01174_ _01230_ _01196_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_105_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout127_A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07154_ net1136 _01953_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06105_ smpl_rt_clkdiv.clkDiv_inst.cnt\[1\] smpl_rt_clkdiv.clkDiv_inst.cnt\[0\] smpl_rt_clkdiv.clkDiv_inst.cnt\[2\]
+ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07085_ genblk1\[8\].osc.clkdiv_C.cnt\[6\] _01895_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12343__A1 genblk2\[11\].wave_shpr.div.acc_next\[0\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfanout102 net104 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08547__B1 _02309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout113 net114 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11775__A _04676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout124 net125 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08011__A2 _01367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout135 net136 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_2
Xfanout146 net150 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_4
Xfanout157 net158 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
Xfanout168 net170 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_4
X_07987_ _02225_ _02681_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__and2_1
Xfanout179 net180 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_4
X_09726_ _04157_ _04204_ _04205_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__a21o_1
X_06938_ genblk1\[6\].osc.clkdiv_C.cnt\[11\] _01777_ _01780_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09511__A2 _04043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09657_ _04009_ _04129_ _04143_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__o21ai_1
X_06869_ _01694_ _01723_ _01724_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ genblk2\[5\].wave_shpr.div.fin_quo\[1\] VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__inv_2
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ net995 _04076_ _04080_ _04092_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__a22o_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08539_ _03235_ _03245_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__or2b_1
XFILLER_0_49_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11550_ genblk2\[8\].wave_shpr.div.b1\[0\] _05417_ genblk2\[8\].wave_shpr.div.acc\[0\]
+ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10501_ genblk2\[4\].wave_shpr.div.acc\[18\] _04738_ net591 VGND VGND VPWR VPWR _04741_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11481_ _05437_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13220_ clknet_leaf_136_clk _00543_ net62 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10432_ genblk2\[4\].wave_shpr.div.acc\[2\] _04688_ _04623_ VGND VGND VPWR VPWR _04689_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08786__B1 _02224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13151_ clknet_leaf_17_clk net532 net80 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10363_ _03833_ net1223 VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__and2_1
XANTENNA__08043__B _01360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12102_ _05759_ _05863_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13082_ clknet_leaf_126_clk _00409_ net61 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10294_ genblk2\[4\].wave_shpr.div.b1\[12\] genblk2\[4\].wave_shpr.div.acc\[12\]
+ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__and2b_1
X_12033_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__and2_1
XANTENNA__08002__A2 _01675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10896__A1 _01514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07210__B1 _01241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06498__B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10648__A1 _03726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12935_ clknet_leaf_30_clk _00264_ net102 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ clknet_leaf_135_clk _00197_ net61 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08069__A2 _01592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11817_ net938 _05652_ _05653_ _05664_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__a22o_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ clknet_leaf_57_clk net270 net183 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ genblk2\[9\].wave_shpr.div.quo\[3\] _05623_ _05624_ net686 VGND VGND VPWR
+ VPWR _00868_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06961__B _01221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11679_ genblk2\[9\].wave_shpr.div.acc\[2\] genblk2\[9\].wave_shpr.div.b1\[2\] VGND
+ VGND VPWR VPWR _05571_ sky130_fd_sc_hd__or2b_1
XFILLER_0_114_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13418_ clknet_leaf_119_clk _00737_ net141 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13349_ clknet_leaf_4_clk _00670_ net45 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09764__S _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11595__A _05441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07910_ _01230_ _01564_ _01889_ _01238_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__a211oi_1
X_08890_ _03595_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__buf_2
XFILLER_0_75_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07841_ _02530_ _02535_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07772_ genblk1\[0\].osc.clkdiv_C.cnt\[1\] _01190_ net34 genblk1\[0\].osc.clkdiv_C.cnt\[0\]
+ _02336_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__o2111a_1
X_09511_ net684 _04043_ _04047_ net764 VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__a22o_1
XANTENNA__10639__A1 _04225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06723_ _01609_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10939__A _05054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09442_ genblk2\[1\].wave_shpr.div.acc\[18\] _04005_ VGND VGND VPWR VPWR _04006_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_78_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_2_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06654_ genblk1\[3\].osc.clkdiv_C.cnt\[13\] _01545_ _01548_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07313__A _01308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09373_ _02213_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__buf_4
X_06585_ _01490_ genblk1\[3\].osc.clkdiv_C.cnt\[13\] _01363_ genblk1\[3\].osc.clkdiv_C.cnt\[15\]
+ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_47_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08324_ _02638_ _02640_ genblk2\[8\].wave_shpr.div.fin_quo\[4\] VGND VGND VPWR VPWR
+ _03031_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08255_ _02960_ _02961_ genblk2\[6\].wave_shpr.div.fin_quo\[6\] _02539_ VGND VGND
+ VPWR VPWR _02962_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_46_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10811__A1 _04855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12365__S _05982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10674__A _04672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07206_ _01989_ VGND VGND VPWR VPWR genblk1\[9\].osc.clkdiv_C.next_cnt\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12013__B1 _03735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08186_ net9 _02744_ _02365_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__nand3_1
XFILLER_0_6_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07137_ genblk1\[9\].osc.clkdiv_C.cnt\[16\] _01936_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06243__A1 genblk1\[0\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07068_ _01862_ _01885_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__nor2_2
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10613__S _04637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06599__A _01441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09709_ genblk2\[2\].wave_shpr.div.b1\[8\] genblk2\[2\].wave_shpr.div.acc\[8\] VGND
+ VGND VPWR VPWR _04189_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10981_ _05074_ genblk1\[6\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12720_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[15\] net183 VGND VGND
+ VPWR VPWR genblk1\[9\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12651_ clknet_leaf_28_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[0\] net89 VGND VGND
+ VPWR VPWR genblk1\[6\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11602_ genblk2\[8\].wave_shpr.div.acc\[12\] _05512_ _05493_ VGND VGND VPWR VPWR
+ _05513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12582_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[3\] net74 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11533_ genblk2\[8\].wave_shpr.div.quo\[19\] _05454_ _05458_ net617 _05463_ VGND
+ VGND VPWR VPWR _00814_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12004__A0 genblk2\[11\].wave_shpr.div.b1\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11464_ net1230 net34 _05237_ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13203_ clknet_leaf_8_clk _00526_ net48 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10415_ _04676_ _01650_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08223__A2 _02308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11395_ genblk2\[8\].wave_shpr.div.acc\[4\] genblk2\[8\].wave_shpr.div.b1\[4\] VGND
+ VGND VPWR VPWR _05371_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13134_ clknet_leaf_115_clk _00459_ net133 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10346_ _04640_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__clkbuf_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12307__A1 net355 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ clknet_leaf_22_clk net377 net95 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10277_ genblk2\[4\].wave_shpr.div.b1\[3\] genblk2\[4\].wave_shpr.div.acc\[3\] VGND
+ VGND VPWR VPWR _04589_ sky130_fd_sc_hd__and2b_1
XFILLER_0_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12016_ _02208_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap2 _04335_ VGND VGND VPWR VPWR net1351 sky130_fd_sc_hd__buf_1
XANTENNA__09487__A1 _04032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12918_ clknet_leaf_39_clk _00249_ net115 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ clknet_leaf_58_clk _00180_ net194 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06370_ genblk1\[1\].osc.clkdiv_C.cnt\[4\] _01313_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__xnor2_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08040_ _02697_ _02698_ _02746_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__nand3_1
XFILLER_0_127_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold903 genblk2\[1\].wave_shpr.div.b1\[11\] VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 PWM.final_in\[6\] VGND VGND VPWR VPWR net1132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 genblk1\[10\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR net1143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold936 genblk2\[5\].wave_shpr.div.i\[2\] VGND VGND VPWR VPWR net1154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 genblk2\[6\].wave_shpr.div.acc\[2\] VGND VGND VPWR VPWR net1165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 sig_norm.quo\[2\] VGND VGND VPWR VPWR net1176 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13516__RESET_B net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09991_ _04377_ _04385_ _04386_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__a21oi_1
Xhold969 genblk2\[9\].wave_shpr.div.b1\[6\] VGND VGND VPWR VPWR net1187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08942_ _03551_ _03633_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__and2_1
X_08873_ sig_norm.acc\[1\] sig_norm.b1\[1\] VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07824_ _02510_ _02511_ genblk2\[0\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR
+ _02531_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07755_ genblk2\[1\].wave_shpr.div.fin_quo\[0\] genblk2\[1\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__or2_1
XANTENNA__10088__A2 _04452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06706_ genblk1\[4\].osc.clkdiv_C.cnt\[13\] _01595_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__xnor2_1
X_07686_ _02023_ _02386_ _02388_ _02389_ _02392_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__o221a_1
XANTENNA__08139__A net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09425_ _03962_ _03987_ _03988_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__a21o_1
X_06637_ net1095 _01535_ _01537_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09356_ genblk2\[0\].wave_shpr.div.acc\[20\] _03800_ net1352 VGND VGND VPWR VPWR
+ _03930_ sky130_fd_sc_hd__or3_1
X_06568_ _01451_ _01478_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08307_ _02349_ _02351_ _02353_ genblk2\[11\].wave_shpr.div.fin_quo\[3\] VGND VGND
+ VPWR VPWR _03014_ sky130_fd_sc_hd__a31oi_1
XANTENNA__12095__S _05787_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09287_ _03771_ _03759_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__or2b_1
XANTENNA__10608__S _00015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06499_ genblk1\[2\].osc.clkdiv_C.cnt\[13\] genblk1\[2\].osc.clkdiv_C.cnt\[0\] net35
+ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__nor3_1
XFILLER_0_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08238_ _02798_ _02931_ _02936_ _02938_ _02944_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06464__A1 genblk1\[1\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07661__B1 _01235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08169_ genblk1\[3\].osc.clkdiv_C.cnt\[8\] _01423_ _02870_ _02871_ _02875_ VGND VGND
+ VPWR VPWR _02876_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10200_ net930 _04518_ _04522_ _04528_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__a22o_1
X_11180_ _03708_ genblk2\[8\].wave_shpr.div.b1\[1\] VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10131_ genblk2\[3\].wave_shpr.div.quo\[24\] _04451_ _04455_ net490 _04476_ VGND
+ VGND VPWR VPWR _00399_ sky130_fd_sc_hd__a221o_1
X_10062_ net1186 _01240_ _04440_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__mux2_1
XANTENNA_hold838_A genblk2\[5\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09469__A1 _01231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12892__RESET_B net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13752_ clknet_leaf_68_clk _01063_ net211 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10964_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__and2_1
XANTENNA__06495__C _01327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12703_ clknet_leaf_89_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[16\] net173 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
X_13683_ clknet_leaf_63_clk _00996_ net190 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10895_ _05031_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09579__S _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12634_ clknet_leaf_16_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[1\] net74 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12565_ clknet_leaf_28_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[4\] net89 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11516_ _05441_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__buf_2
XFILLER_0_13_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12496_ clknet_leaf_102_clk _00058_ net158 VGND VGND VPWR VPWR sig_norm.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11447_ _05420_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11200__A1 _01565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09944__A2 _04253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11378_ genblk2\[7\].wave_shpr.div.i\[3\] _02192_ _05353_ VGND VGND VPWR VPWR _05356_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_21_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11751__A2 _05623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _04632_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__clkbuf_1
X_13117_ clknet_leaf_13_clk _00442_ net52 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ clknet_leaf_135_clk _00375_ net62 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07540_ _02253_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11179__B1_N _03705_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07471_ _02199_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11812__S _05613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09210_ _02170_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__clkbuf_8
X_06422_ _01233_ _01249_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__nor2_1
XANTENNA__07798__A genblk1\[0\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09141_ genblk2\[0\].wave_shpr.div.b1\[13\] genblk2\[0\].wave_shpr.div.acc\[13\]
+ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__and2b_1
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06353_ _01268_ _01298_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__nor2_1
XANTENNA__13768__RESET_B net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08435__A2 _02350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09072_ genblk2\[0\].wave_shpr.div.b1\[12\] _01340_ _03722_ VGND VGND VPWR VPWR _03729_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07310__B _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06284_ _01245_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__buf_4
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08023_ _01229_ _01749_ _02729_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold700 genblk2\[2\].wave_shpr.div.acc\[3\] VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold711 genblk2\[10\].wave_shpr.div.acc\[7\] VGND VGND VPWR VPWR net929 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout207_A net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold722 _00026_ VGND VGND VPWR VPWR net940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold733 genblk2\[10\].wave_shpr.div.acc\[10\] VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 genblk2\[2\].wave_shpr.div.acc\[26\] VGND VGND VPWR VPWR net962 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11767__B genblk1\[9\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold755 genblk2\[1\].wave_shpr.div.acc\[17\] VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 genblk2\[9\].wave_shpr.div.acc\[7\] VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 genblk2\[1\].wave_shpr.div.acc\[7\] VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 genblk2\[9\].wave_shpr.div.acc\[3\] VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ genblk2\[3\].wave_shpr.div.acc\[8\] genblk2\[3\].wave_shpr.div.b1\[8\] VGND
+ VGND VPWR VPWR _04370_ sky130_fd_sc_hd__or2b_1
Xhold799 genblk2\[3\].wave_shpr.div.acc\[13\] VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10950__B1 _05055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08925_ _03590_ _03602_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__nor2_1
X_08856_ _03560_ _03561_ _03562_ _03557_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__a211o_1
XANTENNA__10702__B1 _04856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09253__A _03855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07807_ _02510_ _02513_ genblk2\[0\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR
+ _02514_ sky130_fd_sc_hd__a21oi_1
X_08787_ _03492_ _03493_ genblk2\[2\].wave_shpr.div.fin_quo\[2\] _02468_ VGND VGND
+ VPWR VPWR _03494_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10399__A _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_48_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07738_ _02444_ _02013_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__nor2_1
X_07669_ _01188_ _01440_ genblk1\[10\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR _02376_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_149_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11722__S _00023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09408_ genblk2\[1\].wave_shpr.div.b1\[1\] genblk2\[1\].wave_shpr.div.acc\[1\] VGND
+ VGND VPWR VPWR _03972_ sky130_fd_sc_hd__and2b_1
X_10680_ _04676_ _01670_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09339_ _03917_ _03794_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07220__B _01189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12350_ _05941_ _05942_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11301_ _05221_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_889 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12281_ genblk2\[1\].wave_shpr.div.b1\[9\] _02013_ _05994_ VGND VGND VPWR VPWR _06002_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11232_ net370 _05251_ _05248_ net736 _05254_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10073__S _04440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11163_ genblk2\[7\].wave_shpr.div.fin_quo\[0\] _05222_ _00019_ VGND VGND VPWR VPWR
+ _05223_ sky130_fd_sc_hd__mux2_1
XANTENNA__10941__B1 _05056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10114_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__and2_1
X_11094_ _05055_ _05156_ _05157_ _05057_ net1130 VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__a32o_1
X_10045_ _03714_ _04431_ _03717_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_4_10_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold60 _00132_ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold71 genblk2\[10\].wave_shpr.div.i\[4\] VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 genblk2\[2\].wave_shpr.div.quo\[8\] VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__08362__B2 _02592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold93 _00553_ VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11996_ _05803_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__clkbuf_1
X_13735_ clknet_leaf_46_clk _01046_ net119 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10947_ net515 _05052_ _05056_ net523 VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13666_ clknet_leaf_41_clk net869 net123 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10878_ genblk2\[6\].wave_shpr.div.acc\[25\] genblk2\[6\].wave_shpr.div.acc\[24\]
+ genblk2\[6\].wave_shpr.div.acc\[26\] _05021_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__or4_2
XFILLER_0_38_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12617_ clknet_leaf_18_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[2\] net80 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
X_13597_ clknet_leaf_77_clk _00912_ net208 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07625__B1 _01576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12548_ clknet_leaf_61_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[5\] net186 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__06979__A2 _01363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12479_ clknet_leaf_108_clk _00041_ net152 VGND VGND VPWR VPWR sig_norm.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_2 _04242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09772__S _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ genblk1\[7\].osc.clkdiv_C.cnt\[6\] _01802_ _01805_ genblk1\[7\].osc.clkdiv_C.cnt\[5\]
+ _01806_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__o221a_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _03412_ _03416_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__xnor2_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10711__S _04821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11488__A1 _03726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09690_ genblk2\[2\].wave_shpr.div.acc\[3\] genblk2\[2\].wave_shpr.div.b1\[3\] VGND
+ VGND VPWR VPWR _04170_ sky130_fd_sc_hd__or2b_1
XFILLER_0_83_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08641_ _03345_ _03346_ _03347_ _02694_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__a211o_1
X_08572_ _03277_ _03278_ genblk2\[9\].wave_shpr.div.fin_quo\[2\] _02362_ VGND VGND
+ VPWR VPWR _03279_ sky130_fd_sc_hd__a2bb2o_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07523_ _02227_ net286 _02242_ VGND VGND VPWR VPWR PWM.next_pwm_out sky130_fd_sc_hd__a21o_1
XFILLER_0_76_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout157_A net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07454_ _02147_ _02187_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10666__B genblk1\[5\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06405_ _01172_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__buf_4
XFILLER_0_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07385_ genblk1\[11\].osc.clkdiv_C.cnt\[13\] _02132_ VGND VGND VPWR VPWR _02136_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09124_ _03759_ _03770_ _03771_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__a21o_1
XANTENNA__07040__B _01344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06336_ genblk1\[0\].osc.clkdiv_C.cnt\[10\] _01286_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09055_ _03704_ net394 _03715_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_4_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06267_ _01228_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__buf_6
XANTENNA__12373__S _05982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10682__A _04672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08006_ genblk1\[6\].osc.clkdiv_C.cnt\[1\] _01735_ _01738_ genblk1\[6\].osc.clkdiv_C.cnt\[0\]
+ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__o211a_1
Xhold530 genblk2\[10\].wave_shpr.div.i\[2\] VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__dlygate4sd3_1
X_06198_ _01163_ _01161_ VGND VGND VPWR VPWR PWM.next_counter\[4\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold541 genblk2\[10\].wave_shpr.div.b1\[14\] VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 genblk2\[5\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07919__A1 genblk1\[8\].osc.clkdiv_C.cnt\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold563 genblk2\[4\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07919__B2 genblk1\[8\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold574 genblk2\[6\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__clkbuf_2
Xhold585 genblk2\[1\].wave_shpr.div.acc\[23\] VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 genblk2\[3\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__dlygate4sd3_1
X_09957_ genblk2\[2\].wave_shpr.div.i\[1\] genblk2\[2\].wave_shpr.div.i\[0\] genblk2\[2\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__and3_1
X_08908_ _03610_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10621__S _04834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _04191_ _04164_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__or2b_1
X_08839_ _03540_ _03545_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__nand2_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _05597_ _05689_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__xnor2_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ genblk2\[5\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[12\] VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13520_ clknet_leaf_79_clk _00837_ net206 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10732_ genblk2\[5\].wave_shpr.div.acc\[6\] _04900_ _04821_ VGND VGND VPWR VPWR _04901_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13451_ clknet_leaf_119_clk _00768_ net143 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10663_ net308 _04853_ _04857_ net770 VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12402_ _05967_ _05929_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__or2b_1
X_10594_ genblk2\[5\].wave_shpr.div.fin_quo\[0\] _04821_ _00015_ VGND VGND VPWR VPWR
+ _04822_ sky130_fd_sc_hd__mux2_1
X_13382_ clknet_leaf_83_clk _00701_ net200 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07083__A1 genblk1\[8\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12333_ net239 _06014_ _06015_ net483 _06024_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12264_ _05992_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08032__B1 _02261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11215_ net822 _05246_ _05222_ _05248_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__a22o_1
X_12195_ genblk2\[11\].wave_shpr.div.acc\[9\] genblk2\[11\].wave_shpr.div.b1\[9\]
+ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__or2b_1
XFILLER_0_102_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09592__S _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11146_ _05169_ _05204_ _05205_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11077_ genblk2\[6\].wave_shpr.div.acc\[21\] _05145_ _05146_ VGND VGND VPWR VPWR
+ _05147_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07138__A2 _01246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10028_ _04423_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06346__B1 genblk1\[0\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08099__B1 _02805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11979_ _05794_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06964__B _01799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13718_ clknet_leaf_36_clk _01029_ net105 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13649_ clknet_leaf_38_clk _00962_ net126 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07861__A3 _02459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07170_ genblk1\[9\].osc.clkdiv_C.cnt\[5\] genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01960_
+ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__and3_1
X_06121_ smpl_rt_clkdiv.clkDiv_inst.next_hzX _01093_ VGND VGND VPWR VPWR smpl_rt_clkdiv.clkDiv_inst.next_cnt\[7\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_120_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_120_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09396__B_N genblk2\[1\].wave_shpr.div.b1\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09811_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[1\] VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__and2_1
XANTENNA__06585__B1 _01363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09742_ _04218_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__clkbuf_1
X_06954_ _01791_ VGND VGND VPWR VPWR genblk1\[6\].osc.clkdiv_C.next_cnt\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09523__B1 _04045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09673_ _03690_ _04153_ _04154_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__nor3_1
X_06885_ _01349_ _01209_ _01439_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__and3_2
XFILLER_0_118_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _03307_ _03330_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _02217_ _02553_ genblk2\[6\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR
+ _03262_ sky130_fd_sc_hd__and3_1
XANTENNA__11272__S _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06874__B _01578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07506_ _02218_ _02221_ _02224_ _02226_ VGND VGND VPWR VPWR FSM.next_mode\[1\] sky130_fd_sc_hd__a31oi_1
X_08486_ genblk2\[3\].wave_shpr.div.fin_quo\[4\] _02467_ _03192_ _02592_ VGND VGND
+ VPWR VPWR _03193_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07051__A _01336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07437_ genblk2\[4\].wave_shpr.div.i\[1\] _02174_ genblk2\[4\].wave_shpr.div.i\[4\]
+ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__or3b_1
XFILLER_0_64_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07368_ genblk1\[11\].osc.clkdiv_C.cnt\[9\] _02119_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__and2_1
XANTENNA__07065__A1 genblk1\[8\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09107_ genblk2\[0\].wave_shpr.div.acc\[8\] genblk2\[0\].wave_shpr.div.b1\[8\] VGND
+ VGND VPWR VPWR _03755_ sky130_fd_sc_hd__or2b_1
X_06319_ _01269_ _01276_ _01277_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_111_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_111_clk sky130_fd_sc_hd__clkbuf_16
X_07299_ genblk1\[11\].osc.clkdiv_C.cnt\[9\] _01235_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09038_ _02336_ net34 VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__nand2_2
XFILLER_0_60_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold360 genblk2\[0\].wave_shpr.div.acc_next\[0\] VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 _00232_ VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08565__A1 _02261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold382 genblk2\[0\].wave_shpr.div.quo\[4\] VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ genblk2\[6\].wave_shpr.div.acc\[2\] _05088_ _05023_ VGND VGND VPWR VPWR _05089_
+ sky130_fd_sc_hd__mux2_1
Xhold393 genblk2\[8\].wave_shpr.div.quo\[15\] VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12113__A2 _05844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09514__B1 _04047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12951_ clknet_leaf_125_clk _00280_ net71 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1060 genblk2\[11\].wave_shpr.div.b1\[17\] VGND VGND VPWR VPWR net1278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1071 genblk2\[0\].wave_shpr.div.b1\[7\] VGND VGND VPWR VPWR net1289 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ _05726_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__inv_2
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1082 sig_norm.quo\[7\] VGND VGND VPWR VPWR net1300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1093 genblk2\[7\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net1311 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ clknet_leaf_91_clk _00213_ net146 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold918_A genblk1\[9\].osc.clkdiv_C.cnt\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ genblk2\[9\].wave_shpr.div.acc\[9\] _05676_ _05673_ VGND VGND VPWR VPWR _05677_
+ sky130_fd_sc_hd__mux2_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _02155_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__clkbuf_2
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13503_ clknet_leaf_87_clk _00820_ net180 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _04784_ _04887_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__xnor2_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11695_ _05564_ _05585_ _05586_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09587__S _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07896__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13434_ clknet_leaf_81_clk net1011 net199 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10646_ _04850_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_102_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_102_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13365_ clknet_leaf_12_clk _00684_ net53 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10577_ _04768_ _04803_ _04804_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12316_ _05835_ genblk1\[11\].osc.clkdiv_C.cnt\[3\] VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13296_ clknet_leaf_87_clk _00617_ net179 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12247_ genblk2\[11\].wave_shpr.div.fin_quo\[1\] net1310 _00005_ VGND VGND VPWR VPWR
+ _05984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12178_ genblk2\[10\].wave_shpr.div.i\[1\] genblk2\[10\].wave_shpr.div.i\[0\] genblk2\[10\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__a21o_1
XANTENNA__11560__B1 _05446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06959__B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11129_ _05180_ _05187_ _05188_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12042__A _05815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07136__A genblk1\[9\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06670_ genblk1\[4\].osc.clkdiv_C.cnt\[2\] _01559_ _01557_ genblk1\[4\].osc.clkdiv_C.cnt\[6\]
+ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__a22o_1
XANTENNA__11791__B_N _03693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire27 _01692_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_1
XANTENNA__06975__A _01365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08340_ _03045_ _03046_ _02745_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__o21a_1
XANTENNA__10418__A2 _04651_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09070__B _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08271_ _02409_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11820__S _05613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07222_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] _02001_ _02002_ _02003_ VGND VGND VPWR
+ VPWR _02004_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07153_ _01952_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07084_ _01887_ _01895_ _01896_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08156__A2_N _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08547__A1 genblk2\[6\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout103 net104 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08547__B2 genblk2\[6\].wave_shpr.div.fin_quo\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12343__A2 _03942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09526__A _04042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout114 net126 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_4
Xfanout125 net126 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__buf_2
Xfanout136 net171 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_4
Xfanout147 net171 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_2
Xfanout158 net171 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
X_07986_ _02691_ _02682_ _02690_ _02527_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__o31a_1
Xfanout169 net170 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07770__A2 _01240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09725_ genblk2\[2\].wave_shpr.div.b1\[16\] genblk2\[2\].wave_shpr.div.acc\[16\]
+ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__and2b_1
X_06937_ net28 _01779_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__nor2_1
XANTENNA__11303__B1 _05283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09656_ genblk2\[1\].wave_shpr.div.acc\[24\] _04008_ VGND VGND VPWR VPWR _04143_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__10657__A2 _04853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06868_ genblk1\[5\].osc.clkdiv_C.cnt\[16\] _01721_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__nand2_1
XANTENNA__06885__A _01349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09261__A _03853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08607_ genblk2\[5\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__inv_2
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ genblk2\[1\].wave_shpr.div.acc\[6\] _04091_ _04011_ VGND VGND VPWR VPWR _04092_
+ sky130_fd_sc_hd__mux2_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06799_ genblk1\[5\].osc.clkdiv_C.cnt\[14\] _01210_ _01304_ genblk1\[5\].osc.clkdiv_C.cnt\[1\]
+ _01670_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__a221o_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _03243_ _03244_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08469_ genblk2\[5\].wave_shpr.div.fin_quo\[2\] VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__inv_2
XANTENNA__11730__S _00023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10500_ _04618_ _04738_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11480_ genblk2\[9\].wave_shpr.div.b1\[11\] _01732_ _05433_ VGND VGND VPWR VPWR _05437_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07038__A1 _01436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10431_ _04586_ _04687_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08235__B1 _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12127__A _05815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13150_ clknet_leaf_121_clk net681 net80 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10362_ _03726_ _04649_ _03736_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__o21ai_1
X_12101_ _05760_ _05741_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__or2b_1
XANTENNA__11790__B1 _03693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13081_ clknet_leaf_126_clk _00408_ net63 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10293_ _04571_ _04603_ _04604_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12032_ _02155_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__clkbuf_2
Xhold190 genblk2\[4\].wave_shpr.div.quo\[7\] VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07210__A1 _01359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07303__A2_N _01256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12934_ clknet_leaf_30_clk _00263_ net102 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12865_ clknet_leaf_135_clk _00196_ net61 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11816_ genblk2\[9\].wave_shpr.div.acc\[5\] _05663_ _05613_ VGND VGND VPWR VPWR _05664_
+ sky130_fd_sc_hd__mux2_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap34_A _01794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12796_ clknet_leaf_92_clk _00129_ net149 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ genblk2\[9\].wave_shpr.div.quo\[2\] _05623_ _05624_ net649 VGND VGND VPWR
+ VPWR _00867_ sky130_fd_sc_hd__a22o_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12270__A1 _04229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11678_ genblk2\[9\].wave_shpr.div.acc\[3\] genblk2\[9\].wave_shpr.div.b1\[3\] VGND
+ VGND VPWR VPWR _05570_ sky130_fd_sc_hd__or2b_1
X_13417_ clknet_leaf_119_clk _00736_ net141 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10629_ _04841_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13348_ clknet_leaf_5_clk _00669_ net45 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13279_ clknet_leaf_11_clk _00600_ net56 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10336__A1 _01256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07840_ _02536_ _02546_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__nor2_1
XANTENNA__09780__S _04238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07752__A2 _01577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07771_ _02475_ _02477_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09510_ _04046_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__buf_4
X_06722_ genblk1\[4\].osc.clkdiv_C.cnt\[3\] _01605_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09441_ _03954_ _04003_ _04004_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06653_ _01523_ _01547_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07313__B _01439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09372_ _03940_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__buf_4
XFILLER_0_47_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06584_ genblk1\[3\].osc.clkdiv_C.cnt\[10\] _01231_ _01488_ _01490_ _01491_ VGND
+ VGND VPWR VPWR _01492_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08323_ _03013_ _03029_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12261__A1 _01329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08254_ genblk2\[6\].wave_shpr.div.fin_quo\[5\] _02733_ _02959_ _02261_ VGND VGND
+ VPWR VPWR _02961_ sky130_fd_sc_hd__a31o_1
XFILLER_0_145_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07205_ _01954_ _01987_ _01988_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__and3_1
XANTENNA__06491__A2 _01363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12013__A1 _03726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08185_ genblk2\[3\].wave_shpr.div.fin_quo\[7\] _02539_ VGND VGND VPWR VPWR _02892_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08144__B _01576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07136_ genblk1\[9\].osc.clkdiv_C.cnt\[15\] _01361_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07067_ _01863_ _01872_ _01873_ _01884_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__or4b_1
XANTENNA__06243__A2 _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08160__A _01489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06599__B _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07969_ _02650_ _02667_ _02675_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__a21oi_2
X_09708_ _04166_ _04186_ _04187_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__a21o_1
X_10980_ net609 _05051_ _05064_ net616 _05075_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__a221o_1
XANTENNA__07504__A net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09639_ _04130_ _04131_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12650_ clknet_leaf_10_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[17\] net57 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10566__A_N genblk2\[5\].wave_shpr.div.b1\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08038__C _02365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11601_ _05397_ _05511_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12581_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[2\] net70 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11532_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[10\] VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12004__A1 _01500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11463_ _05428_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08054__B _01223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13202_ clknet_leaf_8_clk _00525_ net55 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10414_ _03719_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__buf_6
X_11394_ genblk2\[8\].wave_shpr.div.acc\[5\] genblk2\[8\].wave_shpr.div.b1\[5\] VGND
+ VGND VPWR VPWR _05370_ sky130_fd_sc_hd__or2b_1
XFILLER_0_110_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13133_ clknet_leaf_0_clk _00458_ net41 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10345_ net1303 _04639_ _04637_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__mux2_1
XANTENNA__12307__A2 _06009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ clknet_leaf_29_clk _00391_ net95 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10276_ _04582_ _04586_ _04587_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__a21o_1
XANTENNA__11515__B1 _05449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12015_ _05811_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10105__A _04269_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06302__B _01263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap3 _03923_ VGND VGND VPWR VPWR net1352 sky130_fd_sc_hd__buf_1
X_12917_ clknet_leaf_35_clk _00248_ net105 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11294__A2 _05279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12848_ clknet_leaf_58_clk _00179_ net194 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12779_ clknet_leaf_41_clk _00112_ net116 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06972__B _01214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09775__S _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold904 genblk2\[6\].wave_shpr.div.acc\[1\] VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 genblk1\[0\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR net1133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold926 genblk2\[4\].wave_shpr.div.acc\[24\] VGND VGND VPWR VPWR net1144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 sig_norm.acc\[6\] VGND VGND VPWR VPWR net1155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold948 genblk1\[2\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR net1166 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ genblk2\[3\].wave_shpr.div.b1\[3\] genblk2\[3\].wave_shpr.div.acc\[3\] VGND
+ VGND VPWR VPWR _04386_ sky130_fd_sc_hd__and2b_1
Xhold959 genblk2\[6\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR net1177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08941_ _03540_ _03550_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11506__B1 _05446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08872_ sig_norm.acc\[0\] VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07823_ _02469_ _02528_ _02529_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__o21ai_1
X_07754_ _02460_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__clkbuf_2
X_06705_ _01489_ _01196_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__nor2_4
XFILLER_0_67_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07685_ _02390_ _02391_ _01995_ _02016_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08139__B _02364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08150__A2 _01234_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09424_ genblk2\[1\].wave_shpr.div.b1\[9\] genblk2\[1\].wave_shpr.div.acc\[9\] VGND
+ VGND VPWR VPWR _03988_ sky130_fd_sc_hd__and2b_1
XANTENNA_hold1002_A genblk1\[11\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06636_ genblk1\[3\].osc.clkdiv_C.cnt\[7\] _01535_ _01524_ VGND VGND VPWR VPWR _01537_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09355_ net1032 _03903_ _03910_ _03929_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__a22o_1
X_06567_ genblk1\[2\].osc.clkdiv_C.cnt\[15\] genblk1\[2\].osc.clkdiv_C.cnt\[14\] _01474_
+ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08306_ _03012_ _02989_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__xnor2_1
X_09286_ _03838_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06498_ genblk1\[2\].osc.clkdiv_C.cnt\[2\] net36 VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08237_ _02939_ _02942_ _02943_ VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08168_ _02872_ _02873_ _02874_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__nand3_1
XFILLER_0_31_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11745__B1 _05624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07119_ genblk1\[9\].osc.clkdiv_C.cnt\[10\] _01227_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10624__S _04834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08099_ genblk1\[4\].osc.clkdiv_C.cnt\[13\] _01498_ _02805_ genblk1\[4\].osc.clkdiv_C.cnt\[12\]
+ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10130_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__and2_1
XANTENNA__06403__A genblk1\[1\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10061_ _03701_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13751_ clknet_leaf_74_clk _01062_ net212 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10963_ net498 _05062_ _05064_ genblk2\[6\].wave_shpr.div.quo\[13\] _05066_ VGND
+ VGND VPWR VPWR _00641_ sky130_fd_sc_hd__a221o_1
XANTENNA__08049__B _01355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_82_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12702_ clknet_leaf_89_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[15\] net173 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_97_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13682_ clknet_leaf_42_clk _00995_ net190 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10894_ genblk2\[6\].wave_shpr.div.fin_quo\[7\] net1349 _00017_ VGND VGND VPWR VPWR
+ _05031_ sky130_fd_sc_hd__mux2_1
X_12633_ clknet_leaf_16_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[0\] net74 VGND VGND
+ VPWR VPWR genblk1\[5\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10236__B1 _04454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12564_ clknet_leaf_29_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[3\] net96 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11515_ genblk2\[8\].wave_shpr.div.quo\[11\] _05448_ _05449_ net469 _05453_ VGND
+ VGND VPWR VPWR _00806_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12495_ clknet_leaf_104_clk _00057_ net153 VGND VGND VPWR VPWR sig_norm.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11446_ genblk2\[8\].wave_shpr.div.fin_quo\[2\] genblk2\[8\].wave_shpr.div.quo\[1\]
+ _00021_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11377_ _00018_ _05353_ net1181 VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12315__A _03941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13116_ clknet_leaf_2_clk _00441_ net52 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ genblk2\[5\].wave_shpr.div.b1\[0\] _01735_ _04440_ VGND VGND VPWR VPWR _04632_
+ sky130_fd_sc_hd__mux2_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09157__A1 _03804_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ clknet_leaf_129_clk _00374_ net65 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ genblk2\[4\].wave_shpr.div.acc\[11\] genblk2\[4\].wave_shpr.div.b1\[11\]
+ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__or2b_1
XFILLER_0_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08380__A2 _01209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_73_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07470_ _02196_ _02153_ genblk2\[8\].wave_shpr.div.busy VGND VGND VPWR VPWR _02199_
+ sky130_fd_sc_hd__and3b_1
XANTENNA__06983__A _01436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06421_ _01336_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__buf_8
XANTENNA__06694__A2 _01313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07798__B genblk1\[0\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09140_ _03751_ _03786_ _03787_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__a21o_1
X_06352_ genblk1\[0\].osc.clkdiv_C.cnt\[16\] genblk1\[0\].osc.clkdiv_C.cnt\[15\] _01295_
+ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06283_ _01173_ _01187_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__or2_2
XFILLER_0_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09071_ _03726_ net1084 _01302_ _03727_ _03728_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__o221a_1
XFILLER_0_32_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08022_ _02709_ _02708_ _02728_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07134__A2_N _01311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold701 genblk2\[2\].wave_shpr.div.acc\[5\] VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold712 genblk2\[3\].wave_shpr.div.acc\[15\] VGND VGND VPWR VPWR net930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold723 genblk2\[3\].wave_shpr.div.acc\[6\] VGND VGND VPWR VPWR net941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold734 genblk2\[2\].wave_shpr.div.acc\[10\] VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 genblk2\[3\].wave_shpr.div.acc\[5\] VGND VGND VPWR VPWR net963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold756 genblk2\[9\].wave_shpr.div.acc\[9\] VGND VGND VPWR VPWR net974 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A2 _01574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold767 genblk2\[11\].wave_shpr.div.acc\[4\] VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 PWM.counter\[3\] VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ genblk2\[3\].wave_shpr.div.acc\[9\] genblk2\[3\].wave_shpr.div.b1\[9\] VGND
+ VGND VPWR VPWR _04369_ sky130_fd_sc_hd__or2b_1
Xhold789 genblk2\[11\].wave_shpr.div.b1\[0\] VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07149__A2_N _01799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08924_ net717 _02260_ _03621_ _03574_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__a22o_1
X_08855_ _03498_ _03553_ _03554_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__nor3_1
XANTENNA__11783__B genblk1\[9\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06877__B _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07806_ genblk2\[0\].wave_shpr.div.fin_quo\[4\] _02512_ VGND VGND VPWR VPWR _02513_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_137_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08786_ genblk2\[2\].wave_shpr.div.fin_quo\[0\] genblk2\[2\].wave_shpr.div.fin_quo\[1\]
+ _03113_ _02224_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__a31o_1
X_07737_ genblk1\[1\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_64_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08123__A2 _01224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06893__A _01308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07668_ genblk1\[10\].osc.clkdiv_C.cnt\[3\] _02374_ _02013_ genblk1\[10\].osc.clkdiv_C.cnt\[2\]
+ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09407_ genblk2\[1\].wave_shpr.div.acc\[0\] genblk2\[1\].wave_shpr.div.b1\[0\] VGND
+ VGND VPWR VPWR _03971_ sky130_fd_sc_hd__or2b_1
X_06619_ genblk1\[3\].osc.clkdiv_C.cnt\[1\] genblk1\[3\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01526_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07599_ _02261_ _02305_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09338_ _03795_ _03747_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07501__B net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09269_ net715 _00000_ _03863_ net578 _03864_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11300_ _05196_ _05298_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12280_ _06001_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11231_ _05074_ genblk1\[7\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07229__A _01229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11162_ _05221_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06133__A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10113_ net514 _04461_ _04462_ net634 _04467_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__a221o_1
X_11093_ genblk2\[6\].wave_shpr.div.i\[1\] genblk2\[6\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _05157_ sky130_fd_sc_hd__nand2_1
X_10044_ net1100 VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__inv_2
Xhold50 _00872_ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06787__B _01658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08362__A2 _02539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold61 sig_norm.i\[3\] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 genblk2\[9\].wave_shpr.div.quo\[9\] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 _00300_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 genblk2\[8\].wave_shpr.div.quo\[13\] VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__dlygate4sd3_1
X_11995_ net1242 _02805_ _05802_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_55_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13734_ clknet_leaf_46_clk net444 net119 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10946_ genblk2\[6\].wave_shpr.div.quo\[7\] _05052_ _05056_ net241 VGND VGND VPWR
+ VPWR _00634_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13665_ clknet_leaf_43_clk _00978_ net123 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10877_ genblk2\[6\].wave_shpr.div.acc\[23\] _05020_ VGND VGND VPWR VPWR _05021_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_85_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12616_ clknet_leaf_18_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[1\] net80 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13596_ clknet_leaf_77_clk net936 net208 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06428__A2 _01304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12547_ clknet_leaf_61_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[4\] net186 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12478_ clknet_leaf_108_clk _00040_ net152 VGND VGND VPWR VPWR sig_norm.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_3 _04242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11429_ _05360_ _05403_ _05404_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08242__B _02309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11185__B2 _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06970_ genblk1\[7\].osc.clkdiv_C.cnt\[5\] _01805_ _01801_ genblk1\[7\].osc.clkdiv_C.cnt\[1\]
+ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__o2bb2a_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08640_ _02216_ _02553_ genblk2\[7\].wave_shpr.div.fin_quo\[3\] VGND VGND VPWR VPWR
+ _03347_ sky130_fd_sc_hd__and3_1
XANTENNA__10696__B1 _04856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08571_ genblk2\[9\].wave_shpr.div.fin_quo\[0\] genblk2\[9\].wave_shpr.div.fin_quo\[1\]
+ _02303_ _02316_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_46_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_16
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07522_ _02227_ net286 _02229_ _02241_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__o22a_1
XANTENNA__07602__A _02308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07453_ genblk2\[6\].wave_shpr.div.busy _02186_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06404_ genblk1\[1\].osc.clkdiv_C.cnt\[14\] _01327_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__and2_1
XANTENNA__07321__B _01359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07384_ genblk1\[11\].osc.clkdiv_C.cnt\[13\] _02132_ VGND VGND VPWR VPWR _02135_
+ sky130_fd_sc_hd__or2_1
X_09123_ genblk2\[0\].wave_shpr.div.b1\[4\] genblk2\[0\].wave_shpr.div.acc\[4\] VGND
+ VGND VPWR VPWR _03771_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06335_ _01269_ _01286_ _01287_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_115_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_863 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09054_ _03714_ net727 _03715_ _03717_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__o211a_1
X_06266_ _01194_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08005_ _02700_ _02703_ _02711_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__a21boi_1
Xhold520 _00378_ VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 genblk2\[4\].wave_shpr.div.quo\[4\] VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__dlygate4sd3_1
X_06197_ net1307 VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__inv_2
Xhold542 modein.delay_in\[1\] VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07919__A2 _01430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold553 genblk2\[1\].wave_shpr.div.quo\[5\] VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 genblk2\[2\].wave_shpr.div.acc\[1\] VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 genblk2\[4\].wave_shpr.div.quo\[2\] VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold586 genblk2\[0\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold597 _00381_ VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08592__A2 _02527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09956_ genblk2\[2\].wave_shpr.div.i\[1\] genblk2\[2\].wave_shpr.div.i\[0\] genblk2\[2\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__a21o_1
XANTENNA__10902__S _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06888__A _01658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08907_ _03609_ net1240 _01157_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__mux2_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ net895 _04282_ _04289_ _04305_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__a22o_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _03542_ _03544_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__and2_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ _03457_ _03459_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__or2b_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _04819_ _04855_ _04951_ _04858_ net1038 VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__a32o_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11780_ genblk2\[9\].wave_shpr.div.quo\[20\] _05628_ _05629_ net362 _05639_ VGND
+ VGND VPWR VPWR _00885_ sky130_fd_sc_hd__a221o_1
XANTENNA__07304__B1 _01925_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09844__A2 _04247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09203__S _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10731_ _04791_ _04899_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10349__S _04637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13450_ clknet_leaf_119_clk _00767_ net143 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10662_ genblk2\[5\].wave_shpr.div.quo\[6\] _04853_ _04857_ net253 VGND VGND VPWR
+ VPWR _00549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06128__A net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12401_ _03941_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__clkbuf_4
X_13381_ clknet_leaf_96_clk _00700_ net167 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10593_ _04820_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__buf_4
XFILLER_0_91_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12332_ _03833_ _02128_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06297__A2_N _01190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12263_ genblk2\[1\].wave_shpr.div.b1\[1\] _01263_ _05802_ VGND VGND VPWR VPWR _05992_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09873__S _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11214_ _05247_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__clkbuf_4
X_12194_ genblk2\[11\].wave_shpr.div.acc\[10\] genblk2\[11\].wave_shpr.div.b1\[10\]
+ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__or2b_1
XANTENNA__09780__A1 _01858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08583__A2 _02308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11145_ genblk2\[7\].wave_shpr.div.b1\[12\] genblk2\[7\].wave_shpr.div.acc\[12\]
+ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11076_ genblk2\[6\].wave_shpr.div.acc\[21\] genblk2\[6\].wave_shpr.div.acc\[20\]
+ _05019_ net1350 VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10027_ genblk2\[3\].wave_shpr.div.fin_quo\[0\] _04420_ _04422_ VGND VGND VPWR VPWR
+ _04423_ sky130_fd_sc_hd__mux2_1
XANTENNA__11209__A _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06897__A2 _01367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11978_ genblk2\[10\].wave_shpr.div.fin_quo\[6\] net1324 _00003_ VGND VGND VPWR VPWR
+ _05794_ sky130_fd_sc_hd__mux2_1
XANTENNA__07422__A _02147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13717_ clknet_leaf_36_clk _01028_ net105 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10929_ net758 VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__inv_2
XANTENNA__11642__A2 _05448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13648_ clknet_leaf_38_clk net224 net126 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13579_ clknet_leaf_76_clk _00894_ net207 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06120_ net365 _01088_ net395 VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13329__RESET_B net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08023__A1 _01229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09220__B1 _03840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09810_ genblk2\[2\].wave_shpr.div.quo\[9\] _04253_ _04251_ net300 _04254_ VGND VGND
+ VPWR VPWR _00300_ sky130_fd_sc_hd__a221o_1
XANTENNA__08574__A2 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09084__A _03735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09741_ genblk2\[2\].wave_shpr.div.fin_quo\[3\] net1329 _00009_ VGND VGND VPWR VPWR
+ _04218_ sky130_fd_sc_hd__mux2_1
X_06953_ _01760_ _01789_ _01790_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__and3b_1
XFILLER_0_94_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10669__B1 _04855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09672_ genblk2\[1\].wave_shpr.div.i\[3\] _02158_ _04151_ VGND VGND VPWR VPWR _04154_
+ sky130_fd_sc_hd__and3_1
X_06884_ _01241_ _01660_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__nor2_2
X_08623_ _03328_ _03329_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_19_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _03259_ _03260_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__nor2_1
X_07505_ _02215_ net760 _02225_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__o21a_1
XANTENNA__11094__B1 _05057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08485_ genblk2\[3\].wave_shpr.div.fin_quo\[3\] _03191_ VGND VGND VPWR VPWR _03192_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07436_ genblk2\[4\].wave_shpr.div.i\[2\] genblk2\[4\].wave_shpr.div.i\[3\] genblk2\[4\].wave_shpr.div.i\[0\]
+ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07051__B _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07367_ _02122_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09106_ genblk2\[0\].wave_shpr.div.acc\[9\] genblk2\[0\].wave_shpr.div.b1\[9\] VGND
+ VGND VPWR VPWR _03754_ sky130_fd_sc_hd__or2b_1
XANTENNA__09259__A _03853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06318_ genblk1\[0\].osc.clkdiv_C.cnt\[3\] _01274_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07065__A2 _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07298_ net695 _02061_ VGND VGND VPWR VPWR genblk1\[10\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09037_ _03704_ net861 _03705_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__a21bo_1
X_06249_ _01182_ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold350 _00648_ VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold361 _00148_ VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 genblk2\[10\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09762__A1 _04230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11728__S _00023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold383 _00128_ VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 sig_norm.acc\[7\] VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10632__S _04834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07773__B1 _01190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09939_ net968 _04315_ _04322_ _04344_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
X_12950_ clknet_leaf_125_clk _00279_ net71 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1050 genblk2\[9\].wave_shpr.div.b1\[4\] VGND VGND VPWR VPWR net1268 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12634__RESET_B net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1061 genblk2\[5\].wave_shpr.div.b1\[12\] VGND VGND VPWR VPWR net1279 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ genblk2\[0\].wave_shpr.div.i\[1\] genblk2\[0\].wave_shpr.div.i\[0\] genblk2\[0\].wave_shpr.div.i\[2\]
+ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__and3_1
Xhold1072 genblk2\[3\].wave_shpr.div.b1\[3\] VGND VGND VPWR VPWR net1290 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ clknet_leaf_91_clk net415 net146 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1083 genblk2\[7\].wave_shpr.div.b1\[12\] VGND VGND VPWR VPWR net1301 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 genblk2\[1\].wave_shpr.div.quo\[1\] VGND VGND VPWR VPWR net1312 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11832_ _05589_ _05675_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__xnor2_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11085__B1 _05055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ net243 _05628_ _05629_ net481 _05630_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__a221o_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__08057__B _01223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _04785_ _04780_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__or2b_1
X_13502_ clknet_leaf_87_clk _00819_ net180 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ genblk2\[9\].wave_shpr.div.b1\[7\] genblk2\[9\].wave_shpr.div.acc\[7\] VGND
+ VGND VPWR VPWR _05586_ sky130_fd_sc_hd__and2b_1
X_13433_ clknet_leaf_82_clk _00752_ net201 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07896__B net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10645_ genblk2\[6\].wave_shpr.div.b1\[15\] _01365_ _04848_ VGND VGND VPWR VPWR _04850_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13364_ clknet_leaf_12_clk _00683_ net53 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10576_ genblk2\[5\].wave_shpr.div.b1\[12\] genblk2\[5\].wave_shpr.div.acc\[12\]
+ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12315_ _03941_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__clkbuf_4
X_13295_ clknet_leaf_53_clk _00616_ net112 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12337__B1 _03941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12246_ _05983_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__10899__B1 _04233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12177_ _05816_ _05917_ _05918_ _05818_ net1090 VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__a32o_1
X_11128_ genblk2\[7\].wave_shpr.div.b1\[3\] genblk2\[7\].wave_shpr.div.acc\[3\] VGND
+ VGND VPWR VPWR _05188_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11059_ genblk2\[6\].wave_shpr.div.acc\[16\] _05133_ _05105_ VGND VGND VPWR VPWR
+ _05134_ sky130_fd_sc_hd__mux2_1
XANTENNA__07136__B _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire28 net1356 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_99_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06975__B _01355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09778__S _04238_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08270_ _02366_ _02976_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07221_ genblk1\[10\].osc.clkdiv_C.cnt\[8\] VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07152_ _01919_ _01922_ _01927_ _01951_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__and4_2
XANTENNA__09079__A _03708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06255__B1 _01215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07083_ genblk1\[8\].osc.clkdiv_C.cnt\[4\] _01892_ genblk1\[8\].osc.clkdiv_C.cnt\[5\]
+ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08547__A2 _02527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout104 net107 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout115 net118 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_4
Xfanout126 net127 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__buf_2
Xfanout137 net145 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_4
Xfanout148 net150 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_4
X_07985_ _02682_ _02690_ _02691_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__o21ai_1
Xfanout159 net162 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06231__A _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09724_ _04158_ _04202_ _04203_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06936_ genblk1\[6\].osc.clkdiv_C.cnt\[11\] _01777_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__and2_1
XANTENNA__07046__B _01328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09655_ _04045_ _04141_ _04142_ _04048_ net448 VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__a32o_1
X_06867_ genblk1\[5\].osc.clkdiv_C.cnt\[16\] _01721_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06885__B _01209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08606_ _02891_ _03311_ _03312_ _02893_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__a31o_1
XFILLER_0_145_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__09261__B genblk1\[0\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _03981_ _04090_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__xnor2_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06798_ genblk1\[5\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _03240_ _03242_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10814__B1 _04858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08468_ _03154_ _03173_ _03051_ _03174_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_65_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07419_ genblk2\[2\].wave_shpr.div.i\[2\] genblk2\[2\].wave_shpr.div.i\[3\] genblk2\[2\].wave_shpr.div.i\[0\]
+ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08399_ _03103_ _03104_ _03105_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__or3b_1
XFILLER_0_107_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08605__B _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10430_ _04587_ _04582_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__or2b_1
XFILLER_0_33_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08235__A1 _02592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07038__A2 _01855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10361_ net834 VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06125__B _01095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12100_ net929 _05844_ _05850_ _05862_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__a22o_1
X_13080_ clknet_leaf_125_clk _00407_ net63 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10292_ genblk2\[4\].wave_shpr.div.b1\[11\] genblk2\[4\].wave_shpr.div.acc\[11\]
+ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__and2b_1
XFILLER_0_131_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12886__RESET_B net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12031_ _05812_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09735__A1 _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold180 genblk2\[10\].wave_shpr.div.quo\[10\] VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 genblk2\[1\].wave_shpr.div.b1\[17\] VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08943__C1 _01155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06141__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07210__A2 _01224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12933_ clknet_leaf_31_clk _00262_ net102 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ clknet_leaf_129_clk _00195_ net64 VGND VGND VPWR VPWR genblk2\[2\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _05662_ _05581_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__xnor2_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12795_ clknet_leaf_92_clk net601 net148 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ net649 _05623_ _05624_ net746 VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11677_ _05567_ _05568_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13416_ clknet_leaf_119_clk net535 net141 VGND VGND VPWR VPWR genblk2\[7\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10628_ net1211 _01189_ _04834_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13347_ clknet_leaf_5_clk _00668_ net45 VGND VGND VPWR VPWR genblk2\[6\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11230__B1 _05248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10559_ genblk2\[5\].wave_shpr.div.b1\[3\] genblk2\[5\].wave_shpr.div.acc\[3\] VGND
+ VGND VPWR VPWR _04787_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13278_ clknet_leaf_11_clk _00599_ net56 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12229_ genblk2\[11\].wave_shpr.div.b1\[13\] genblk2\[11\].wave_shpr.div.acc\[13\]
+ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07147__A _01241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07770_ genblk1\[0\].osc.clkdiv_C.cnt\[12\] _01240_ _02476_ VGND VGND VPWR VPWR _02477_
+ sky130_fd_sc_hd__a21bo_1
X_06721_ _01608_ VGND VGND VPWR VPWR genblk1\[4\].osc.clkdiv_C.next_cnt\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09440_ genblk2\[1\].wave_shpr.div.b1\[17\] genblk2\[1\].wave_shpr.div.acc\[17\]
+ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__and2b_1
X_06652_ genblk1\[3\].osc.clkdiv_C.cnt\[13\] genblk1\[3\].osc.clkdiv_C.cnt\[12\] _01543_
+ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09371_ _02170_ genblk2\[11\].wave_shpr.div.busy _02211_ VGND VGND VPWR VPWR _03940_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_59_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06583_ genblk1\[3\].osc.clkdiv_C.cnt\[5\] _01250_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08322_ _02419_ _03018_ _03022_ _03024_ _03028_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__a32o_1
XANTENNA__09662__A0 _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08253_ _02734_ _02959_ genblk2\[6\].wave_shpr.div.fin_quo\[5\] VGND VGND VPWR VPWR
+ _02960_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07204_ genblk1\[9\].osc.clkdiv_C.cnt\[16\] _01985_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08184_ _02225_ _02885_ VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__11221__B1 _05250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07135_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01311_ _01925_ genblk1\[9\].osc.clkdiv_C.cnt\[5\]
+ _01934_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07066_ genblk1\[8\].osc.clkdiv_C.cnt\[16\] _01578_ _01870_ genblk1\[8\].osc.clkdiv_C.cnt\[11\]
+ _01883_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07968_ _02672_ _02674_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__or2_1
XANTENNA__06896__A _01342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09707_ genblk2\[2\].wave_shpr.div.b1\[7\] genblk2\[2\].wave_shpr.div.acc\[7\] VGND
+ VGND VPWR VPWR _04187_ sky130_fd_sc_hd__and2b_1
X_06919_ genblk1\[6\].osc.clkdiv_C.cnt\[5\] genblk1\[6\].osc.clkdiv_C.cnt\[4\] _01765_
+ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__and3_1
X_07899_ _01181_ _01852_ _01245_ genblk1\[8\].osc.clkdiv_C.cnt\[13\] VGND VGND VPWR
+ VPWR _02606_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08153__B1 _01494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09638_ _04005_ _04129_ genblk2\[1\].wave_shpr.div.acc\[18\] VGND VGND VPWR VPWR
+ _04131_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09569_ _03973_ _04077_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11600_ _05398_ _05363_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__or2b_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12580_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[1\] net70 VGND VGND
+ VPWR VPWR genblk1\[2\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_833 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11531_ genblk2\[8\].wave_shpr.div.quo\[18\] _05454_ _05458_ net263 _05462_ VGND
+ VGND VPWR VPWR _00813_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_831 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11462_ net1294 _01797_ _05237_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06136__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13201_ clknet_leaf_114_clk _00524_ net132 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08759__A2 _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10413_ net698 _04651_ _04654_ net665 _04675_ VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11393_ genblk2\[8\].wave_shpr.div.acc\[6\] genblk2\[8\].wave_shpr.div.b1\[6\] VGND
+ VGND VPWR VPWR _05369_ sky130_fd_sc_hd__or2b_1
X_13132_ clknet_leaf_3_clk _00457_ net46 VGND VGND VPWR VPWR genblk2\[5\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10344_ _01678_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11188__S _05042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ clknet_leaf_29_clk _00390_ net95 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10275_ genblk2\[4\].wave_shpr.div.b1\[2\] genblk2\[4\].wave_shpr.div.acc\[2\] VGND
+ VGND VPWR VPWR _04587_ sky130_fd_sc_hd__and2b_1
XANTENNA__07719__B1 _01209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12014_ _02171_ net1278 VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap4 net1354 VGND VGND VPWR VPWR net1353 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11217__A _05249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12916_ clknet_leaf_35_clk _00247_ net105 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ clknet_leaf_58_clk _00178_ net211 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ clknet_leaf_41_clk _00111_ net123 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11729_ _05617_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold905 genblk2\[2\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 PWM.final_in\[0\] VGND VGND VPWR VPWR net1134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 genblk1\[3\].osc.clkdiv_C.cnt\[9\] VGND VGND VPWR VPWR net1145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold938 sig_norm.quo\[9\] VGND VGND VPWR VPWR net1156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold949 genblk1\[2\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR net1167 sky130_fd_sc_hd__dlygate4sd3_1
X_08940_ _03632_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08871_ sig_norm.b1\[1\] sig_norm.acc\[1\] VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__or2b_1
X_07822_ net7 net150 _02312_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__and3_2
XFILLER_0_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07605__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09092__A _01367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07753_ _02458_ _02459_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__and2_1
XANTENNA__13596__RESET_B net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06704_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01592_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__or2_1
X_07684_ _01179_ _01575_ genblk1\[10\].osc.clkdiv_C.cnt\[15\] VGND VGND VPWR VPWR
+ _02391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08139__C _02365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09423_ _03963_ _03985_ _03986_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__a21o_1
XANTENNA__06697__B1 _01304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06635_ _01523_ _01535_ _01536_ VGND VGND VPWR VPWR genblk1\[3\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__10966__A _04676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09354_ genblk2\[0\].wave_shpr.div.acc\[20\] _03927_ VGND VGND VPWR VPWR _03929_
+ sky130_fd_sc_hd__xor2_1
X_06566_ net1207 _01474_ _01477_ VGND VGND VPWR VPWR genblk1\[2\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08305_ _02977_ _02983_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11442__A0 genblk2\[8\].wave_shpr.div.fin_quo\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09285_ net1033 _03870_ _03840_ _03876_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__a22o_1
XANTENNA__10177__S _04507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07110__A1 genblk1\[8\].osc.clkdiv_C.cnt\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06497_ _01173_ _01191_ _01175_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_34_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10796__A2 _04858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08236_ net9 _02744_ _02365_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07661__A2 _01190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08167_ genblk1\[3\].osc.clkdiv_C.cnt\[9\] _01231_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12478__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11745__B2 _05613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07118_ net691 _01917_ VGND VGND VPWR VPWR genblk1\[8\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__09267__A _03838_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08098_ _01440_ _01576_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__nand2_2
XANTENNA__08602__C _02885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07049_ genblk1\[8\].osc.clkdiv_C.cnt\[4\] _01866_ _01865_ genblk1\[8\].osc.clkdiv_C.cnt\[9\]
+ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06403__B _01327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10060_ _04439_ VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11736__S _00023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10962_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[5\] VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__and2_1
XANTENNA__07234__B _01359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13750_ clknet_leaf_75_clk _01061_ net211 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13266__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12701_ clknet_leaf_89_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[14\] net172 VGND VGND
+ VPWR VPWR genblk1\[8\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
X_13681_ clknet_leaf_63_clk _00994_ net125 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10893_ _05030_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12632_ clknet_leaf_18_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[17\] net112 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_155_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12563_ clknet_leaf_30_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[2\] net96 VGND VGND
+ VPWR VPWR genblk1\[1\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__07101__A1 genblk1\[8\].osc.clkdiv_C.cnt\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11984__A1 _03813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11514_ _04676_ _01879_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12494_ clknet_leaf_106_clk _00056_ net153 VGND VGND VPWR VPWR sig_norm.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11445_ _05419_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11376_ _05248_ _05352_ _05354_ _05251_ net801 VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10327_ net1264 VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__clkbuf_1
X_13115_ clknet_leaf_115_clk _00440_ net135 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07409__B _02153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ clknet_leaf_112_clk _00373_ net128 VGND VGND VPWR VPWR genblk2\[4\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10258_ genblk2\[4\].wave_shpr.div.acc\[12\] genblk2\[4\].wave_shpr.div.b1\[12\]
+ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__or2b_1
X_10189_ _04402_ _04519_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09865__B1 _04252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__06679__B1 _01242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06983__B _01334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06420_ genblk1\[1\].osc.clkdiv_C.cnt\[16\] _01363_ _01341_ VGND VGND VPWR VPWR _01364_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07798__C _01209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07160__A genblk1\[9\].osc.clkdiv_C.cnt\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06351_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] _01295_ _01297_ VGND VGND VPWR VPWR genblk1\[0\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09093__A1 _01367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09093__B2 _01342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09070_ _03702_ _01996_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__nand2_4
X_06282_ genblk1\[0\].osc.clkdiv_C.cnt\[16\] _01242_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08021_ genblk1\[6\].osc.clkdiv_C.cnt\[15\] _01577_ _02704_ VGND VGND VPWR VPWR _02728_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold702 genblk2\[0\].wave_shpr.div.acc\[13\] VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 genblk2\[11\].wave_shpr.div.acc\[21\] VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 genblk2\[3\].wave_shpr.div.acc\[12\] VGND VGND VPWR VPWR net942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold735 genblk2\[2\].wave_shpr.div.acc\[13\] VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06504__A _01224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold746 genblk2\[0\].wave_shpr.div.acc\[7\] VGND VGND VPWR VPWR net964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold757 genblk2\[2\].wave_shpr.div.acc\[4\] VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 genblk2\[6\].wave_shpr.div.acc\[4\] VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ genblk2\[3\].wave_shpr.div.acc\[10\] genblk2\[3\].wave_shpr.div.b1\[10\]
+ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__or2b_1
XANTENNA__10026__A _04421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold779 genblk2\[11\].wave_shpr.div.acc\[7\] VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10950__A2 _05057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08923_ _03589_ _03602_ _03620_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09815__A _04247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08854_ _03500_ _03503_ _03501_ _03502_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__o211ai_1
XANTENNA__06906__A1 _01675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10702__A2 _02183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07805_ genblk2\[0\].wave_shpr.div.fin_quo\[3\] _02511_ VGND VGND VPWR VPWR _02512_
+ sky130_fd_sc_hd__or2_1
X_08785_ genblk2\[2\].wave_shpr.div.fin_quo\[0\] _03113_ genblk2\[2\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07736_ _02441_ _02437_ _02439_ _02442_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__o22a_1
XANTENNA__09856__B1 _04253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08123__A3 _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07667_ _01308_ _01187_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__nor2_4
XFILLER_0_79_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06893__B _01577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06618_ genblk1\[3\].osc.clkdiv_C.cnt\[1\] genblk1\[3\].osc.clkdiv_C.cnt\[0\] VGND
+ VGND VPWR VPWR _01525_ sky130_fd_sc_hd__nand2_1
X_09406_ genblk2\[1\].wave_shpr.div.acc\[1\] genblk2\[1\].wave_shpr.div.b1\[1\] VGND
+ VGND VPWR VPWR _03970_ sky130_fd_sc_hd__xnor2_1
X_07598_ genblk2\[9\].wave_shpr.div.fin_quo\[6\] _02304_ VGND VGND VPWR VPWR _02305_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09337_ net1050 _03903_ _03910_ _03916_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__a22o_1
X_06549_ genblk1\[2\].osc.clkdiv_C.cnt\[9\] _01464_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__and2_1
XANTENNA__11966__A1 _05787_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09268_ _02171_ genblk1\[0\].osc.clkdiv_C.cnt\[17\] VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__or2_1
XANTENNA__07634__A2 _01190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08219_ _02602_ _02924_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__xor2_1
XFILLER_0_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09199_ net1292 _03827_ _03822_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__mux2_1
XANTENNA__10635__S _04834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11230_ genblk2\[7\].wave_shpr.div.quo\[10\] _05251_ _05248_ net302 _05253_ VGND
+ VGND VPWR VPWR _00721_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11161_ _05219_ _05220_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06133__B net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10941__A2 _05052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10112_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[6\] VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11092_ genblk2\[6\].wave_shpr.div.i\[1\] genblk2\[6\].wave_shpr.div.i\[0\] VGND
+ VGND VPWR VPWR _05156_ sky130_fd_sc_hd__or2_1
X_10043_ _03732_ net1071 _03733_ VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__o21a_1
Xhold40 _00228_ VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 genblk2\[0\].wave_shpr.div.quo\[6\] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__buf_1
Xhold62 genblk2\[6\].wave_shpr.div.i\[4\] VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 _00875_ VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 genblk2\[7\].wave_shpr.div.quo\[9\] VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 genblk2\[6\].wave_shpr.div.quo\[19\] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11994_ _03707_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__clkbuf_8
X_13733_ clknet_leaf_45_clk net468 net121 VGND VGND VPWR VPWR genblk2\[11\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10945_ net241 _05052_ _05056_ net742 VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13664_ clknet_leaf_43_clk _00977_ net124 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10876_ genblk2\[6\].wave_shpr.div.acc\[22\] genblk2\[6\].wave_shpr.div.acc\[21\]
+ genblk2\[6\].wave_shpr.div.acc\[20\] _05019_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__or4_1
XFILLER_0_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12615_ clknet_leaf_121_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[0\] net81 VGND VGND
+ VPWR VPWR genblk1\[4\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13595_ clknet_leaf_72_clk _00910_ net216 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07625__A2 _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12546_ clknet_leaf_61_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[3\] net188 VGND VGND
+ VPWR VPWR genblk1\[0\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12477_ clknet_leaf_107_clk _00039_ net152 VGND VGND VPWR VPWR sig_norm.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12326__A _03689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 _04242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11428_ genblk2\[8\].wave_shpr.div.b1\[15\] genblk2\[8\].wave_shpr.div.acc\[15\]
+ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_880 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11359_ genblk2\[7\].wave_shpr.div.acc\[23\] _05219_ VGND VGND VPWR VPWR _05343_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_67_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ clknet_leaf_113_clk _00356_ net131 VGND VGND VPWR VPWR genblk2\[3\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12061__A _02155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08570_ genblk2\[9\].wave_shpr.div.fin_quo\[0\] _02303_ genblk2\[9\].wave_shpr.div.fin_quo\[1\]
+ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07521_ _02228_ PWM.final_sample_in\[6\] _02231_ _02240_ VGND VGND VPWR VPWR _02241_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07452_ genblk2\[6\].wave_shpr.div.i\[1\] _02185_ genblk2\[6\].wave_shpr.div.i\[4\]
+ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__or3b_1
XANTENNA__12000__S _05802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06403_ genblk1\[1\].osc.clkdiv_C.cnt\[14\] _01327_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07383_ _02134_ VGND VGND VPWR VPWR genblk1\[11\].osc.clkdiv_C.next_cnt\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09122_ _03760_ _03768_ _03769_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06334_ genblk1\[0\].osc.clkdiv_C.cnt\[9\] _01284_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09053_ _03716_ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__buf_8
X_06265_ _01224_ _01226_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__nor2_8
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout212_A net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08004_ genblk1\[6\].osc.clkdiv_C.cnt\[11\] _01519_ _02708_ _02710_ VGND VGND VPWR
+ VPWR _02711_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_5_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold510 genblk2\[0\].wave_shpr.div.quo\[3\] VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06196_ _01161_ _01162_ VGND VGND VPWR VPWR PWM.next_counter\[3\] sky130_fd_sc_hd__nor2_1
XFILLER_0_13_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold521 genblk2\[6\].wave_shpr.div.i\[2\] VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 _00464_ VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 genblk2\[2\].wave_shpr.div.b1\[17\] VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 genblk2\[5\].wave_shpr.div.acc\[9\] VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 genblk2\[5\].wave_shpr.div.i\[3\] VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10384__B1 _04655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold576 genblk2\[3\].wave_shpr.div.quo\[0\] VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold587 genblk2\[7\].wave_shpr.div.acc\[14\] VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 genblk2\[11\].wave_shpr.div.acc\[10\] VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ _04251_ _04353_ _04354_ _04253_ net1110 VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__a32o_1
XANTENNA__06888__B _01675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10190__S _04507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08906_ sig_norm.acc\[3\] _03596_ _03608_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__o21a_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ genblk2\[2\].wave_shpr.div.acc\[8\] _04304_ _04301_ VGND VGND VPWR VPWR _04305_
+ sky130_fd_sc_hd__mux2_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08349__A_N _02789_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08837_ _02574_ _03543_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11884__B1 _03694_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _03455_ _03456_ _03459_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__o21ba_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11636__B1 _05448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07719_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] _01309_ _01209_ genblk1\[1\].osc.clkdiv_C.cnt\[14\]
+ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__o22ai_2
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ _03401_ _03404_ _03405_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__nand3b_2
X_10730_ _04792_ _04774_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__or2b_1
XFILLER_0_137_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10661_ net253 _04853_ _04857_ net729 VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__12493__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06128__B net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12400_ _03942_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__clkbuf_4
X_13380_ clknet_leaf_80_clk _00699_ net200 VGND VGND VPWR VPWR genblk2\[8\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10592_ _04818_ _04819_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12331_ net483 _06014_ _06015_ net509 _06023_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12262_ _05991_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__clkbuf_1
X_11213_ _02170_ genblk2\[7\].wave_shpr.div.busy _02191_ VGND VGND VPWR VPWR _05247_
+ sky130_fd_sc_hd__and3_1
X_12193_ genblk2\[11\].wave_shpr.div.acc\[11\] genblk2\[11\].wave_shpr.div.b1\[11\]
+ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__or2b_1
XFILLER_0_102_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11144_ _05170_ _05202_ _05203_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11075_ genblk2\[6\].wave_shpr.div.acc\[20\] _05019_ net1350 VGND VGND VPWR VPWR
+ _05145_ sky130_fd_sc_hd__or3_1
XANTENNA__10127__B1 _04455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10026_ _04421_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08099__A2 _01498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11977_ _05793_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__clkbuf_1
X_13716_ clknet_leaf_36_clk _01027_ net103 VGND VGND VPWR VPWR genblk2\[1\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10928_ _05048_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09048__A1 _03712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13647_ clknet_leaf_47_clk _00960_ net114 VGND VGND VPWR VPWR genblk2\[10\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10859_ _04973_ _05001_ _05002_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07059__B1 _01869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13578_ clknet_leaf_78_clk _00893_ net207 VGND VGND VPWR VPWR genblk2\[9\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12529_ clknet_leaf_59_clk _00081_ net187 VGND VGND VPWR VPWR genblk2\[0\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09220__B2 net804 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08574__A3 _02350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07782__A1 genblk1\[0\].osc.clkdiv_C.cnt\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09740_ _04217_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__clkbuf_1
X_06952_ genblk1\[6\].osc.clkdiv_C.cnt\[16\] _01787_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__nand2_1
.ends

