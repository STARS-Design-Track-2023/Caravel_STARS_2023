* NGSPICE file created from Eighty_Twos.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt Eighty_Twos VGND VPWR clk cs gpi[0] gpi[10] gpi[11] gpi[12] gpi[13] gpi[14]
+ gpi[15] gpi[16] gpi[17] gpi[18] gpi[19] gpi[1] gpi[20] gpi[21] gpi[22] gpi[23] gpi[24]
+ gpi[25] gpi[26] gpi[27] gpi[28] gpi[29] gpi[2] gpi[30] gpi[31] gpi[32] gpi[33] gpi[3]
+ gpi[4] gpi[5] gpi[6] gpi[7] gpi[8] gpi[9] gpo[0] gpo[10] gpo[11] gpo[12] gpo[13]
+ gpo[14] gpo[15] gpo[16] gpo[17] gpo[18] gpo[19] gpo[1] gpo[20] gpo[21] gpo[22] gpo[23]
+ gpo[24] gpo[25] gpo[26] gpo[27] gpo[28] gpo[29] gpo[2] gpo[30] gpo[31] gpo[32] gpo[33]
+ gpo[3] gpo[4] gpo[5] gpo[6] gpo[7] gpo[8] gpo[9] nrst
X_2037_ ByteBuffer.instr\[19\] _0260_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__nand2_4
X_2409__9 clknet_1_1__leaf__0515_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__inv_2
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2106_ _0630_ _0285_ _1202_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2655_ net109 _0131_ net58 VGND VGND VPWR VPWR RegFile.D\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1606_ RegFile.A\[7\] _0792_ _0704_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__or3_1
X_2586_ PC.i_mem_addr\[15\] _0611_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__xnor2_1
X_1537_ ALU.flags_to_alu\[1\] _0711_ _0878_ _0654_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__a211oi_1
X_1399_ RegFile.A\[1\] _0704_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__nor2_1
X_1468_ ALU.flags_to_alu\[2\] _0765_ _0763_ RegFile.H\[2\] VGND VGND VPWR VPWR _0810_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2371_ _0495_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
X_1322_ _0626_ _0657_ _0635_ _0659_ _0663_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__o311a_4
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2569_ _0601_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__clkbuf_1
X_2638_ net92 _0114_ net58 VGND VGND VPWR VPWR RegFile.H\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1871_ _1156_ _1211_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__or2_1
X_1940_ _0922_ _1253_ _0175_ _1093_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2354_ _0486_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
X_1305_ _0624_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__inv_2
X_2285_ _0448_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2445__44 clknet_1_0__leaf__0516_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__inv_2
X_2460__58 clknet_1_0__leaf__0517_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__inv_2
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2070_ _0655_ _0285_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1785_ _0937_ _1056_ _1063_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__or3_2
X_1923_ _0937_ _1210_ _1259_ _1261_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__o211a_1
X_1854_ _1194_ _1195_ _0626_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2406_ clknet_2_0__leaf_clk VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__buf_1
XFILLER_0_12_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2199_ _0376_ _0374_ _0375_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2268_ _0260_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__inv_2
X_2337_ _0732_ _0476_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1570_ _0882_ _0910_ _0911_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__a21oi_2
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2122_ _0248_ RegFile.H\[0\] _0307_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__mux2_1
X_2053_ _0274_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1906_ _1244_ _1245_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__nor2_2
X_1837_ _0960_ _1162_ _1170_ _1178_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__a211o_1
X_1768_ _0908_ _0885_ _0896_ _1109_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__a31o_1
X_1699_ _0622_ _0624_ _0621_ _1040_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2471__5 clknet_1_0__leaf__0514_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__inv_2
Xoutput42 net42 VGND VGND VPWR VPWR gpo[6] sky130_fd_sc_hd__clkbuf_4
Xoutput20 net20 VGND VGND VPWR VPWR gpo[17] sky130_fd_sc_hd__clkbuf_4
Xoutput31 net31 VGND VGND VPWR VPWR gpo[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2671_ net125 _0147_ net59 VGND VGND VPWR VPWR RegFile.B\[5\] sky130_fd_sc_hd__dfrtp_4
X_1622_ RegFile.L\[6\] _0770_ _0763_ RegFile.H\[6\] net143 VGND VGND VPWR VPWR _0964_
+ sky130_fd_sc_hd__a221oi_1
X_1553_ _0893_ _0894_ _0693_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__o21a_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1484_ RegFile.C\[2\] _0705_ _0707_ RegFile.L\[2\] _0825_ VGND VGND VPWR VPWR _0826_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2036_ _0621_ _0628_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__nor2_2
X_2105_ _0305_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2585_ _0614_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__clkbuf_1
X_1605_ _0780_ _0946_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__nand2_4
X_2654_ net108 _0130_ net58 VGND VGND VPWR VPWR RegFile.D\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1536_ RegFile.C\[1\] _0705_ _0707_ RegFile.L\[1\] _0877_ VGND VGND VPWR VPWR _0878_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1398_ RegFile.A\[1\] _0652_ _0676_ _0739_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__o211ai_4
X_1467_ RegFile.D\[2\] _0767_ _0807_ _0808_ net50 VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__a2111o_1
X_2019_ _0250_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__buf_4
XFILLER_0_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2370_ _0417_ ALU.immediate\[15\] _0406_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__mux2_1
X_1321_ _0645_ _0662_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__nor2_1
X_2466__64 clknet_1_1__leaf__0517_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__inv_2
XFILLER_0_24_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2499_ PC.i_mem_addr\[0\] _0541_ _0542_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__mux2_1
X_2568_ PC.i_mem_addr\[11\] _0600_ _0542_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__mux2_1
X_1519_ ALU.flags_to_alu\[1\] _0765_ _0761_ RegFile.E\[1\] VGND VGND VPWR VPWR _0861_
+ sky130_fd_sc_hd__a22o_1
X_2637_ net91 _0113_ net58 VGND VGND VPWR VPWR RegFile.H\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1870_ _0983_ _1155_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2353_ net129 _0437_ _0430_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2284_ RegFile.A\[6\] net1 VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__and2_1
X_1304_ _0619_ _0640_ _0644_ _0632_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1999_ _0885_ _0896_ _1172_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1922_ _1072_ _1172_ _1260_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__o21ba_1
X_1784_ _1121_ _1124_ _1125_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__and3_1
X_1853_ _0647_ _0656_ _0660_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__or3b_1
XFILLER_0_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2336_ _0478_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
X_2405_ _0513_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
X_2198_ _0374_ _0375_ _0376_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2267_ net134 _0410_ _0409_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2121_ _0314_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2052_ RegFile.C\[5\] _0273_ _0269_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__mux2_1
X_1905_ _1011_ _1241_ _1243_ _1049_ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1836_ _0908_ net49 _1165_ _1177_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__a31o_1
X_1698_ _0619_ _0620_ _0647_ ByteBuffer.instr\[19\] _1039_ VGND VGND VPWR VPWR _1040_
+ sky130_fd_sc_hd__a221o_1
X_1767_ ALU.flags_to_alu\[0\] VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2319_ PC.i_mem_addr\[10\] _0451_ _0468_ _0441_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__o211a_1
X_2415__15 clknet_1_0__leaf__0515_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__inv_2
XFILLER_0_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2430__29 clknet_1_0__leaf__0516_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__inv_2
Xoutput21 net21 VGND VGND VPWR VPWR gpo[18] sky130_fd_sc_hd__clkbuf_4
Xoutput43 net43 VGND VGND VPWR VPWR gpo[7] sky130_fd_sc_hd__clkbuf_4
Xoutput32 net32 VGND VGND VPWR VPWR gpo[28] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1552_ ALU.flags_to_alu\[0\] _0711_ _0707_ RegFile.L\[0\] _0654_ VGND VGND VPWR VPWR
+ _0894_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2670_ net124 _0146_ net59 VGND VGND VPWR VPWR RegFile.B\[4\] sky130_fd_sc_hd__dfrtp_4
X_1621_ ALU.flags_to_alu\[6\] _0765_ _0767_ RegFile.D\[6\] _0962_ VGND VGND VPWR VPWR
+ _0963_ sky130_fd_sc_hd__a221oi_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1483_ RegFile.E\[2\] _0703_ _0699_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__o21a_1
X_2104_ RegFile.E\[0\] _0283_ _0297_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2035_ _0259_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1819_ _1092_ _1160_ _1151_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2584_ PC.i_mem_addr\[14\] _0613_ _0542_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1604_ _0629_ _0943_ _0944_ _0945_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__o22a_2
X_1535_ RegFile.E\[1\] _0699_ net56 VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__and3_1
X_2653_ net107 _0129_ net58 VGND VGND VPWR VPWR RegFile.D\[3\] sky130_fd_sc_hd__dfrtp_1
X_1397_ RegFile.H\[1\] net53 _0738_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__a21o_1
X_1466_ RegFile.L\[2\] _0638_ _0681_ _0762_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__and4_1
XFILLER_0_49_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2018_ _1188_ _1191_ _1201_ _1193_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1320_ ByteBuffer.instr\[22\] _0618_ _0660_ _0661_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__and4_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2636_ net90 _0112_ net58 VGND VGND VPWR VPWR RegFile.H\[2\] sky130_fd_sc_hd__dfrtp_2
X_2567_ net46 _0598_ _0599_ _0585_ ALU.immediate\[11\] VGND VGND VPWR VPWR _0600_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2498_ _0659_ _0411_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__nor2_8
X_1518_ RegFile.B\[1\] _0771_ _0763_ RegFile.H\[1\] VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1449_ ALU.flags_to_alu\[5\] _0788_ _0790_ _0711_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2352_ net131 _0415_ _0438_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1303_ ByteBuffer.instr\[23\] VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__buf_8
X_2283_ _0447_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1998_ _1059_ _1140_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2619_ net73 _0095_ net60 VGND VGND VPWR VPWR ALU.flags_to_alu\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1921_ _0934_ _1255_ _1164_ _0855_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__a22o_1
X_1852_ _0622_ ByteBuffer.instr\[19\] _0624_ _0619_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__a211o_1
X_2451__49 clknet_1_1__leaf__0517_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__inv_2
X_2436__35 clknet_1_0__leaf__0516_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__inv_2
X_1783_ _1101_ _1120_ _1098_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2335_ _0744_ _0476_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__and2_1
X_2266_ net140 _0412_ _0415_ _0627_ _0438_ VGND VGND VPWR VPWR FSM.next_state\[1\]
+ sky130_fd_sc_hd__a221o_1
X_2404_ _0417_ ALU.immediate\[7\] _0408_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__mux2_1
X_2197_ _0855_ _1092_ _0346_ _0174_ _0181_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_46_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold10 ALU.flags_to_alu\[4\] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2120_ _0229_ RegFile.H\[1\] net48 VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2051_ _1239_ _0261_ _0262_ net8 VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__a22o_2
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1904_ _1241_ _1243_ _1011_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1835_ _1172_ _1067_ _1176_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1697_ ByteBuffer.instr\[20\] _0622_ _0624_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__and3_1
X_1766_ _0885_ _0896_ _0908_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2318_ _0207_ _0451_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__nand2_1
X_2249_ net3 net5 VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__or2b_1
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput22 net22 VGND VGND VPWR VPWR gpo[19] sky130_fd_sc_hd__clkbuf_4
Xoutput33 net33 VGND VGND VPWR VPWR gpo[29] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput44 net44 VGND VGND VPWR VPWR gpo[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1551_ RegFile.C\[0\] _0705_ _0709_ RegFile.E\[0\] VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__a22o_1
X_1482_ RegFile.A\[2\] _0792_ _0704_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__or3_1
X_1620_ RegFile.C\[6\] _0638_ _0681_ _0760_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__and4_1
XFILLER_0_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2103_ _0304_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2034_ _0248_ RegFile.B\[0\] _0251_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1818_ _1122_ _1159_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__and2_2
XFILLER_0_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1749_ _1047_ _1048_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2652_ net106 _0128_ net58 VGND VGND VPWR VPWR RegFile.D\[2\] sky130_fd_sc_hd__dfrtp_2
X_2583_ _0540_ _0611_ _0612_ _0585_ ALU.immediate\[14\] VGND VGND VPWR VPWR _0613_
+ sky130_fd_sc_hd__a32o_1
X_1603_ RegFile.L\[7\] net53 net52 RegFile.C\[7\] VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__a22o_1
X_1534_ _0870_ _0871_ _0875_ _0741_ _0789_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__a32o_1
X_1465_ RegFile.C\[2\] _0638_ _0681_ _0760_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2017_ _0249_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__clkbuf_1
X_1396_ RegFile.D\[1\] _0683_ net52 RegFile.B\[1\] _0687_ VGND VGND VPWR VPWR _0738_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2635_ net89 _0111_ net60 VGND VGND VPWR VPWR RegFile.H\[1\] sky130_fd_sc_hd__dfrtp_2
X_2497_ _0522_ _0455_ net46 VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__mux2_1
X_2566_ PC.i_mem_addr\[9\] PC.i_mem_addr\[10\] _0582_ PC.i_mem_addr\[11\] VGND VGND
+ VPWR VPWR _0599_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1517_ RegFile.D\[1\] _0767_ _0857_ _0858_ net51 VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1448_ RegFile.E\[5\] _0789_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2457__55 clknet_1_1__leaf__0517_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__inv_2
X_1379_ RegFile.A\[3\] _0652_ _0676_ _0720_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__o211a_2
XFILLER_0_52_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2351_ net133 _0430_ _0431_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__o21a_1
X_1302_ _0618_ _0641_ _0635_ _0642_ _0643_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__o221ai_4
X_2282_ RegFile.A\[5\] net1 VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1997_ _0230_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2549_ _0534_ _0537_ _0520_ _0539_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__o211a_2
X_2618_ net72 _0094_ net60 VGND VGND VPWR VPWR ALU.flags_to_alu\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_30_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1920_ _0781_ _1253_ _1256_ _0922_ _1258_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__o221a_1
X_1851_ _0700_ _1185_ _1187_ ByteBuffer.instr\[21\] _0645_ VGND VGND VPWR VPWR _1193_
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_21_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1782_ net49 _1123_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__nor2_2
X_2403_ _0512_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2265_ _0431_ _0437_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__nor2_1
X_2196_ _0372_ _0373_ _0360_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__o21ai_1
X_2334_ _0477_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold11 ALU.flags_to_alu\[5\] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2050_ _0272_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__clkbuf_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1903_ _1000_ _1020_ _1242_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__a21o_1
X_1834_ _1174_ _1175_ _0947_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__mux2_1
X_1765_ _0868_ _0881_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1696_ _0715_ _1026_ _1037_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2179_ _0356_ _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__xnor2_2
X_2317_ _0467_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
X_2248_ net7 _0416_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput23 net23 VGND VGND VPWR VPWR gpo[1] sky130_fd_sc_hd__buf_2
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput12 net12 VGND VGND VPWR VPWR gpo[0] sky130_fd_sc_hd__clkbuf_4
Xoutput34 net34 VGND VGND VPWR VPWR gpo[2] sky130_fd_sc_hd__clkbuf_4
Xoutput45 net45 VGND VGND VPWR VPWR gpo[9] sky130_fd_sc_hd__clkbuf_4
X_1550_ _0886_ _0888_ _0890_ _0891_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__o31a_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1481_ _0819_ _0821_ _0822_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2102_ RegFile.E\[1\] _0281_ _0297_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__mux2_1
X_2033_ _0258_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__clkbuf_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1748_ _1037_ _1089_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1817_ ByteBuffer.instr\[21\] _0645_ _1045_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2420__20 clknet_1_1__leaf__0515_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__inv_2
X_1679_ _1014_ _1018_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2582_ PC.i_mem_addr\[14\] _0606_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__or2_1
X_2651_ net105 _0127_ net60 VGND VGND VPWR VPWR RegFile.D\[1\] sky130_fd_sc_hd__dfrtp_1
X_1602_ ALU.flags_to_alu\[7\] _0687_ _0683_ RegFile.E\[7\] _0654_ VGND VGND VPWR VPWR
+ _0944_ sky130_fd_sc_hd__a221o_1
X_1395_ _0736_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__inv_2
X_1464_ _0804_ _0805_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__nor2_2
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1533_ RegFile.L\[1\] _0817_ _0872_ _0873_ _0874_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__a2111oi_1
X_2016_ RegFile.A\[0\] _0248_ _1203_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2565_ _0597_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__inv_2
X_2703_ clknet_2_1__leaf_clk ByteBuffer.next_counter\[1\] net62 VGND VGND VPWR VPWR
+ ByteBuffer.counter\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2634_ net88 _0110_ net61 VGND VGND VPWR VPWR RegFile.H\[0\] sky130_fd_sc_hd__dfrtp_2
X_1516_ RegFile.C\[1\] _0638_ _0681_ _0760_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__and4_1
X_2496_ _0534_ _0537_ _0539_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__o21ai_4
X_1447_ _0678_ _0785_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__nand2_4
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1378_ RegFile.H\[3\] net53 _0719_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2350_ _0485_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
X_1301_ ByteBuffer.instr\[21\] _0624_ ByteBuffer.instr\[17\] ByteBuffer.instr\[20\]
+ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__or4bb_1
X_2281_ _0446_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1996_ RegFile.A\[1\] _0229_ _1203_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2548_ PC.i_mem_addr\[6\] PC.i_mem_addr\[7\] _0567_ PC.i_mem_addr\[8\] VGND VGND
+ VPWR VPWR _0584_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2617_ clknet_2_0__leaf_clk _0093_ net62 VGND VGND VPWR VPWR ALU.immediate\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2479_ _0678_ _0636_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1781_ _1047_ _1122_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__nand2_4
X_1850_ _1188_ _1191_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__nand2_4
XFILLER_0_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2402_ _0428_ ALU.immediate\[6\] _0408_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__mux2_1
X_2333_ _0752_ _0476_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2195_ _0360_ _0372_ _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__or3_1
X_2264_ net9 _0417_ _0432_ _0436_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1979_ _1108_ _1110_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__nand2_1
Xhold12 ByteDecoder.state\[1\] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2441__40 clknet_1_1__leaf__0516_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__inv_2
XFILLER_0_67_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1902_ _1151_ _1021_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1764_ _0816_ _0831_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__nand2_1
X_1833_ net49 _1173_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__nand2_2
XFILLER_0_32_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2316_ _0441_ _0466_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__and2_1
X_1695_ _1034_ _1036_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__nand2_1
X_2247_ net8 _0416_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__and2_1
X_2178_ _0908_ _0231_ _1092_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput24 net24 VGND VGND VPWR VPWR gpo[20] sky130_fd_sc_hd__buf_2
XFILLER_0_43_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput35 net35 VGND VGND VPWR VPWR gpo[30] sky130_fd_sc_hd__clkbuf_4
Xoutput13 net13 VGND VGND VPWR VPWR gpo[10] sky130_fd_sc_hd__buf_2
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1480_ RegFile.C\[2\] _0793_ _0786_ RegFile.D\[2\] VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__a22o_1
X_2032_ _0229_ RegFile.B\[1\] _0251_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__mux2_1
X_2101_ _0303_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__clkbuf_1
X_1678_ _1019_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__inv_2
X_1816_ _0960_ _1157_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__xnor2_1
X_1747_ _0718_ _1088_ _0716_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2581_ PC.i_mem_addr\[14\] _0606_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__nand2_1
X_1601_ _0939_ _0941_ _0942_ _0774_ RegFile.A\[7\] VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__o32a_1
X_1532_ RegFile.E\[1\] _0789_ _0699_ _0703_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2650_ net104 _0126_ net61 VGND VGND VPWR VPWR RegFile.D\[0\] sky130_fd_sc_hd__dfrtp_1
X_1394_ _0734_ _0735_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__and2_1
X_1463_ _0781_ _0803_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2015_ _0655_ _0242_ _0247_ _0631_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2702_ clknet_2_1__leaf_clk ByteBuffer.next_counter\[0\] net62 VGND VGND VPWR VPWR
+ ByteBuffer.counter\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2564_ PC.i_mem_addr\[10\] PC.i_mem_addr\[11\] _0588_ VGND VGND VPWR VPWR _0597_
+ sky130_fd_sc_hd__and3_1
X_2495_ _0525_ _0527_ _0538_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__or3_2
X_2633_ net87 _0109_ net60 VGND VGND VPWR VPWR RegFile.L\[7\] sky130_fd_sc_hd__dfrtp_2
X_1515_ RegFile.L\[1\] _0638_ _0681_ _0762_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__and4_1
X_1446_ _0783_ _0708_ _0703_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__and3_4
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1377_ RegFile.D\[3\] _0683_ net52 RegFile.B\[3\] _0687_ VGND VGND VPWR VPWR _0719_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2448__46 clknet_1_0__leaf__0517_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__inv_2
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1300_ ByteBuffer.instr\[17\] _0624_ ByteBuffer.instr\[19\] _0619_ VGND VGND VPWR
+ VPWR _0642_ sky130_fd_sc_hd__and4bb_4
X_2280_ RegFile.A\[4\] net1 VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1995_ _0655_ _0223_ _0228_ _0631_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a22o_2
X_2616_ clknet_2_0__leaf_clk _0092_ net59 VGND VGND VPWR VPWR ALU.immediate\[6\] sky130_fd_sc_hd__dfrtp_2
X_2462__60 clknet_1_0__leaf__0517_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__inv_2
XFILLER_0_15_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2547_ _0582_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2478_ ALU.immediate\[0\] _0520_ _0521_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1429_ net57 _0650_ _0766_ _0638_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__o211a_4
XFILLER_0_2_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1780_ _0645_ _1044_ _1045_ ByteBuffer.instr\[19\] VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__o211a_2
XFILLER_0_24_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2401_ _0511_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
X_2332_ _0475_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__inv_2
X_2194_ _0364_ _0365_ _0371_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__and3_1
X_2263_ net2 _0433_ _0434_ _0435_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__and4b_1
XFILLER_0_46_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1978_ _1141_ _0211_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold13 ALU.flags_to_alu\[3\] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1901_ _1022_ _1085_ _1240_ _1151_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1832_ _1151_ _1173_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1763_ _0937_ _1104_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1694_ _1035_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__inv_2
X_2315_ PC.i_mem_addr\[9\] _0228_ _0451_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__mux2_1
X_2246_ net5 net3 VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__or2b_1
XFILLER_0_67_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2177_ _0781_ _1049_ _0355_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput36 net36 VGND VGND VPWR VPWR gpo[31] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput25 net25 VGND VGND VPWR VPWR gpo[21] sky130_fd_sc_hd__clkbuf_4
Xoutput14 net14 VGND VGND VPWR VPWR gpo[11] sky130_fd_sc_hd__clkbuf_4
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2100_ RegFile.E\[2\] _0279_ _0297_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2031_ _0257_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__clkbuf_1
X_1815_ _1069_ _1153_ _1156_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1677_ _1014_ _1018_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__nor2_1
X_1746_ _1011_ _1022_ _1085_ _1087_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2229_ _0405_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2411__11 clknet_1_0__leaf__0515_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__inv_2
XFILLER_0_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2580_ _0610_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__clkbuf_1
X_1462_ _0781_ _0803_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1600_ RegFile.L\[7\] _0770_ _0763_ RegFile.H\[7\] net50 VGND VGND VPWR VPWR _0942_
+ sky130_fd_sc_hd__a221o_1
X_1531_ RegFile.D\[1\] _0785_ net54 _0703_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__and4_1
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1393_ _0729_ _0733_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2014_ _0245_ _0246_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__nor2_2
XFILLER_0_9_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1729_ _0782_ _0802_ _0781_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2701_ clknet_2_2__leaf_clk FSM.next_state\[1\] net63 VGND VGND VPWR VPWR ByteDecoder.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_42_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2632_ net86 _0108_ net59 VGND VGND VPWR VPWR RegFile.L\[6\] sky130_fd_sc_hd__dfrtp_2
X_2563_ _0596_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1514_ _0844_ _0855_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__and2b_1
X_2494_ ByteBuffer.instr\[21\] _0621_ _0648_ _0647_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__o211a_1
X_1445_ RegFile.H\[5\] _0784_ _0786_ RegFile.D\[5\] VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__a22o_1
X_1376_ _0716_ _0717_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout60 net64 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_8
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1994_ _0227_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2615_ clknet_2_1__leaf_clk _0091_ net62 VGND VGND VPWR VPWR ALU.immediate\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2546_ PC.i_mem_addr\[7\] PC.i_mem_addr\[8\] _0573_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2477_ _0903_ _0906_ _0519_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__and3_1
X_1428_ _0638_ _0681_ _0762_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__and3_2
X_1359_ _0645_ _0700_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2400_ _0420_ ALU.immediate\[5\] _0408_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2262_ net3 _0416_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__and2_1
X_2331_ net1 net4 _0451_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__nand3_1
XFILLER_0_62_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2193_ _0364_ _0365_ _0371_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1977_ _1139_ _1059_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2529_ PC.i_mem_addr\[4\] _0556_ PC.i_mem_addr\[5\] VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold14 ALU.flags_to_alu\[6\] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1900_ _1086_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__inv_2
X_1831_ ByteBuffer.instr\[21\] _0670_ _1044_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2432__31 clknet_1_1__leaf__0516_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__inv_2
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1762_ _0855_ _0844_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__and2b_1
X_1693_ _1029_ _1033_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2176_ net49 _1229_ _1235_ _1092_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__o211a_1
X_2245_ net9 _0417_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__nand2_1
X_2314_ _0465_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput37 net37 VGND VGND VPWR VPWR gpo[32] sky130_fd_sc_hd__buf_2
Xoutput26 net26 VGND VGND VPWR VPWR gpo[22] sky130_fd_sc_hd__clkbuf_4
Xoutput15 net15 VGND VGND VPWR VPWR gpo[12] sky130_fd_sc_hd__buf_2
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2030_ _0209_ RegFile.B\[2\] _0251_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1745_ _1008_ _1086_ _1010_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__a21oi_1
X_1814_ _0983_ _1155_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1676_ ALU.immediate\[12\] _0675_ _0693_ _1017_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2159_ _1182_ _0338_ _0339_ _0341_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__or4_1
X_2228_ ALU.flags_to_alu\[0\] _0404_ _0334_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1392_ _0729_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__nand2_1
X_1461_ _0782_ _0802_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__nand2_1
X_1530_ RegFile.B\[1\] _0785_ net54 net56 VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__and4_1
XFILLER_0_22_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2013_ _0756_ _0243_ _0244_ _1049_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1728_ _1069_ _0982_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__nand2_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1659_ RegFile.D\[5\] _0683_ net52 RegFile.B\[5\] _0687_ VGND VGND VPWR VPWR _1001_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2562_ PC.i_mem_addr\[10\] _0595_ _0542_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2700_ clknet_2_2__leaf_clk net130 net63 VGND VGND VPWR VPWR ByteDecoder.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2631_ net85 _0107_ net61 VGND VGND VPWR VPWR RegFile.L\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1375_ _0690_ _0714_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__nor2_1
X_2493_ _0535_ _0536_ _0387_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__mux2_1
X_1513_ _0854_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__clkbuf_4
X_1444_ _0785_ net54 _0703_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__and3_2
XFILLER_0_65_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout61 net64 VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_4
XFILLER_0_24_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1993_ _1054_ _0225_ _0226_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2545_ _0581_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__clkbuf_1
X_2614_ clknet_2_1__leaf_clk _0090_ net62 VGND VGND VPWR VPWR ALU.immediate\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2476_ _0519_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__inv_2
X_1358_ ByteBuffer.instr\[22\] VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__inv_2
X_1427_ ALU.flags_to_alu\[5\] _0765_ _0767_ RegFile.D\[5\] _0768_ VGND VGND VPWR VPWR
+ _0769_ sky130_fd_sc_hd__a221o_1
X_1289_ _0618_ _0621_ _0630_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__o21a_2
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2453__51 clknet_1_0__leaf__0517_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__inv_2
XFILLER_0_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2330_ _0474_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
X_2192_ _0207_ _0370_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2261_ net5 _0416_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1976_ _0210_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__clkbuf_1
X_2528_ PC.i_mem_addr\[4\] PC.i_mem_addr\[5\] _0556_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2418__18 clknet_1_0__leaf__0515_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__inv_2
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1761_ _1101_ _1102_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1830_ _1171_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__buf_2
X_1692_ _1029_ _1033_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__nand2_1
X_2313_ _0441_ _0464_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__and2_1
X_2175_ _0348_ _0353_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__xnor2_1
X_2244_ net10 _0416_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__and2_2
XFILLER_0_43_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1959_ _0912_ _0193_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput16 net16 VGND VGND VPWR VPWR gpo[13] sky130_fd_sc_hd__buf_2
Xoutput27 net27 VGND VGND VPWR VPWR gpo[23] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput38 net38 VGND VGND VPWR VPWR gpo[33] sky130_fd_sc_hd__clkbuf_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1744_ _1014_ _1018_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__or2b_1
X_1813_ _1132_ _1154_ _0804_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_25_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1675_ RegFile.A\[4\] _0704_ _1016_ _0630_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__o211a_2
X_2158_ _1221_ _1239_ _1265_ _0340_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__or4_1
X_2227_ _0283_ _0403_ _1201_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__mux2_1
X_2089_ _1192_ _0655_ _0287_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1391_ ALU.immediate\[10\] _0675_ _0693_ _0732_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1460_ _0630_ _0798_ _0801_ _0693_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_22_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2012_ _0243_ _0244_ _0756_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__a21oi_1
X_1658_ _0726_ _0997_ _0999_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__a21oi_1
X_1727_ _1068_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1589_ RegFile.C\[4\] _0705_ _0707_ RegFile.L\[4\] VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2561_ net46 _0593_ _0594_ _0585_ ALU.immediate\[10\] VGND VGND VPWR VPWR _0595_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2492_ _0636_ _0525_ _0697_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__and3b_1
X_1512_ _0780_ _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__and2_1
X_2630_ net84 _0106_ net60 VGND VGND VPWR VPWR RegFile.L\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_65_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1374_ _0690_ _0714_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__and2_1
X_1443_ _0645_ _0647_ _0642_ _0672_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__a22o_2
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout62 net64 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_6
XFILLER_0_36_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2439__38 clknet_1_1__leaf__0516_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__inv_2
X_1992_ _1054_ _0225_ _1049_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__a21oi_1
X_2544_ PC.i_mem_addr\[7\] _0580_ _0542_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__mux2_1
X_2613_ clknet_2_0__leaf_clk _0089_ net62 VGND VGND VPWR VPWR ALU.immediate\[3\] sky130_fd_sc_hd__dfrtp_1
X_2475_ _0518_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1288_ _0629_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__buf_8
X_1357_ _0694_ _0698_ _0648_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__a21o_4
X_1426_ RegFile.C\[5\] _0638_ _0681_ _0760_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__and4_1
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2191_ _0366_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__xnor2_1
X_2260_ _0417_ _0428_ _0418_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1975_ RegFile.A\[2\] _0209_ _1203_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2527_ ALU.immediate\[5\] _0565_ _0519_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1409_ RegFile.B\[0\] _0705_ _0750_ _0711_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__a211o_1
X_2389_ _0505_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1760_ _1100_ _0805_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1691_ ALU.immediate\[15\] _0675_ _0693_ _1032_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2312_ PC.i_mem_addr\[8\] _0247_ _0451_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__mux2_1
X_2243_ net4 net1 VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__and2b_1
X_2174_ _0350_ _0352_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput28 net28 VGND VGND VPWR VPWR gpo[24] sky130_fd_sc_hd__buf_2
Xoutput17 net17 VGND VGND VPWR VPWR gpo[14] sky130_fd_sc_hd__clkbuf_4
X_1889_ _1132_ _1154_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1958_ _0911_ _0882_ _0910_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__and3_1
Xoutput39 net39 VGND VGND VPWR VPWR gpo[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1743_ _1052_ _0736_ _1082_ _1084_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__a31o_1
X_1812_ _0935_ _0938_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1674_ RegFile.B\[4\] _0705_ _1015_ _0711_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__a211o_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _0392_ _0398_ _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2157_ _0182_ _0203_ _0223_ _0242_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2088_ _0296_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1390_ RegFile.A\[2\] _0704_ _0731_ _0630_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__o211a_1
X_2011_ _1043_ _0990_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1657_ _0998_ _0725_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__nor2_1
X_1726_ _0780_ _0969_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1588_ ALU.flags_to_alu\[4\] _0699_ _0703_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__and3_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2209_ _0279_ _0387_ _1201_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2467__1 clknet_1_1__leaf__0514_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__inv_2
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2560_ PC.i_mem_addr\[10\] _0588_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2491_ _0678_ _0526_ _0531_ _0523_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__o211a_1
X_1511_ _0629_ _0850_ _0851_ _0852_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__o22a_1
X_1442_ _0783_ _0708_ net56 VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__and3_4
XFILLER_0_65_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1373_ _0691_ _0714_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2689_ clknet_2_3__leaf_clk _0165_ net63 VGND VGND VPWR VPWR PC.i_mem_addr\[7\] sky130_fd_sc_hd__dfrtp_1
X_1709_ _1037_ _0715_ _1026_ _1050_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__o31ai_2
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout63 net64 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1991_ _0224_ _1080_ _1043_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2612_ clknet_2_0__leaf_clk _0088_ net59 VGND VGND VPWR VPWR ALU.immediate\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2543_ _0578_ _0579_ net46 VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2474_ _0659_ _0669_ _0648_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__and3_1
X_1425_ net57 _0650_ _0766_ _0684_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__o211a_2
X_1287_ _0623_ _0628_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__nor2_8
X_1356_ _0695_ _0696_ _0672_ _0642_ _0697_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_65_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2190_ _0247_ _0368_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1974_ _0655_ _0203_ _0208_ _0631_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__a22o_2
XFILLER_0_1_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2388_ _0417_ _0645_ _0497_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__mux2_1
X_2526_ _0630_ _0775_ _0778_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1408_ RegFile.H\[0\] _0707_ _0709_ RegFile.D\[0\] VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1339_ _0619_ _0640_ _0644_ _0632_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__a22o_4
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1690_ RegFile.A\[7\] _0704_ _1031_ _0630_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__o211a_1
X_2311_ _1182_ _0454_ _0463_ _0441_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__o211a_1
X_2242_ ByteDecoder.state\[1\] ByteDecoder.state\[0\] VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2173_ _0196_ _1092_ _1093_ _0211_ _0351_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__o221a_1
X_1957_ _1057_ _1107_ _1111_ _1236_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__a31o_1
X_2423__23 clknet_1_1__leaf__0515_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__inv_2
Xoutput18 net18 VGND VGND VPWR VPWR gpo[15] sky130_fd_sc_hd__clkbuf_4
X_2509_ PC.i_mem_addr\[1\] PC.i_mem_addr\[0\] PC.i_mem_addr\[2\] VGND VGND VPWR VPWR
+ _0551_ sky130_fd_sc_hd__and3_1
X_1888_ _1134_ _1227_ _1207_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput29 net29 VGND VGND VPWR VPWR gpo[25] sky130_fd_sc_hd__clkbuf_4
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1811_ _0982_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__inv_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1742_ _0721_ _0725_ _1083_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1673_ RegFile.H\[4\] _0707_ _0709_ RegFile.D\[4\] VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__a22o_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _0346_ _1038_ _0400_ _0401_ _0630_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__o311a_1
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2156_ _0228_ _0247_ _0630_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2087_ RegFile.D\[0\] _0248_ _0288_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2010_ _1043_ _1079_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1725_ _1066_ _0959_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__nand2_1
X_1656_ _0721_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__inv_2
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1587_ _0923_ _0928_ _0629_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__a21o_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2208_ _0655_ _0377_ _0378_ _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__o31ai_2
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2139_ _0283_ RegFile.L\[0\] _0316_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2490_ _0523_ _0529_ _0533_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__o21ai_2
X_1441_ _0672_ _0642_ _0624_ _0670_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__o2bb2a_1
X_1510_ RegFile.L\[3\] net53 net52 RegFile.C\[3\] VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1372_ ALU.immediate\[14\] _0675_ _0693_ _0713_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2688_ clknet_2_3__leaf_clk _0164_ net64 VGND VGND VPWR VPWR PC.i_mem_addr\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1708_ _1043_ _1049_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__nor2_2
XFILLER_0_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1639_ _0654_ _0980_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__or2_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout64 net11 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1990_ _0756_ _0990_ _0993_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2542_ PC.i_mem_addr\[7\] _0573_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2611_ clknet_2_0__leaf_clk _0087_ net59 VGND VGND VPWR VPWR ALU.immediate\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_50_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1355_ ByteBuffer.instr\[20\] VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__inv_2
X_1424_ _0670_ _0757_ _0759_ _0650_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1286_ _0624_ _0626_ _0627_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__or3_4
XFILLER_0_46_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2444__43 clknet_1_0__leaf__0516_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__inv_2
XFILLER_0_64_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1973_ _0207_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2525_ _0564_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1407_ RegFile.A\[0\] _0652_ _0676_ _0748_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__o211a_1
X_2387_ _0504_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
X_1338_ _0677_ _0679_ _0638_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2310_ PC.i_mem_addr\[7\] _0451_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2241_ ByteDecoder.state\[1\] _0412_ _0413_ net129 _0414_ VGND VGND VPWR VPWR FSM.next_state\[0\]
+ sky130_fd_sc_hd__a221o_1
X_2172_ _1050_ _0217_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1887_ _1136_ _1146_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__or2_1
X_1956_ _1107_ _1111_ _1057_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2508_ PC.i_mem_addr\[1\] PC.i_mem_addr\[0\] PC.i_mem_addr\[2\] VGND VGND VPWR VPWR
+ _0550_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput19 net19 VGND VGND VPWR VPWR gpo[16] sky130_fd_sc_hd__clkbuf_4
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap50 net143 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1810_ _1130_ _1148_ _1149_ _1151_ _1123_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__a2111oi_1
X_1741_ _0721_ _0725_ _0729_ _0733_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1672_ RegFile.A\[4\] _0652_ _0676_ _1013_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__o211ai_4
X_2224_ _1034_ _1089_ _1035_ _1093_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__a211o_1
X_2155_ _1094_ _0186_ _0337_ _0630_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__o31a_1
XFILLER_0_0_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2086_ _0295_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__clkbuf_1
X_1939_ _0855_ _1175_ _1214_ _0816_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1724_ _0780_ _0946_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1655_ _0737_ _0746_ _0994_ _0996_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__a31o_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1586_ RegFile.L\[4\] _0817_ _0924_ _0925_ _0927_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__a2111o_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _0655_ _0385_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__nand2_1
X_2138_ _0323_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
X_2069_ _0265_ _1191_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1440_ ALU.immediate\[5\] _0675_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__nand2_1
X_1371_ RegFile.A\[6\] _0704_ _0712_ _0630_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2465__63 clknet_1_0__leaf__0517_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__inv_2
XFILLER_0_14_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2687_ clknet_2_3__leaf_clk _0163_ net64 VGND VGND VPWR VPWR PC.i_mem_addr\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1707_ _1047_ _1048_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__nand2_8
XFILLER_0_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1638_ ALU.flags_to_alu\[6\] _0711_ _0709_ RegFile.E\[6\] _0979_ VGND VGND VPWR VPWR
+ _0980_ sky130_fd_sc_hd__a221o_1
X_1569_ _0816_ _0831_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__xnor2_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2541_ ALU.immediate\[7\] _0946_ _0519_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__mux2_1
X_2610_ clknet_2_0__leaf_clk _0086_ net62 VGND VGND VPWR VPWR ALU.immediate\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1285_ ByteDecoder.state\[1\] ByteDecoder.state\[0\] VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__nand2_1
X_1354_ _0619_ _0624_ _0622_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__or3b_2
X_1423_ net57 _0650_ _0762_ _0684_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__o211a_2
XFILLER_0_25_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1972_ _0736_ _0205_ _0206_ _1049_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__a211o_2
XFILLER_0_7_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2524_ PC.i_mem_addr\[4\] _0563_ _0542_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2386_ _0428_ ByteBuffer.instr\[22\] _0497_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__mux2_1
X_1406_ RegFile.B\[0\] _0685_ _0747_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__a21o_1
X_1337_ _0622_ _0624_ _0678_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__or3_4
XFILLER_0_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2240_ ByteDecoder.state\[0\] VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__inv_2
X_2171_ _1050_ _0194_ _0349_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1955_ _1143_ _0189_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1886_ _1226_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2507_ ALU.immediate\[2\] _0815_ _0519_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2369_ _0494_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2414__14 clknet_1_0__leaf__0515_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__inv_2
XFILLER_0_19_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap51 _0772_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1740_ _1054_ _1080_ _1081_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1671_ RegFile.H\[4\] net53 _1012_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__a21o_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2223_ _0399_ _1033_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__nor2_1
X_2154_ _1224_ _1246_ _1268_ _0208_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__or4_1
X_2085_ RegFile.D\[1\] _0229_ _0288_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1938_ _1113_ _1275_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__xnor2_2
X_1869_ net49 _1160_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__nand2_2
XFILLER_0_31_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1654_ _0995_ _0733_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__nor2_1
X_1723_ _0806_ _0937_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__nor2_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ _0182_ _0384_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__xnor2_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1585_ ALU.flags_to_alu\[4\] _0788_ _0926_ _0711_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2068_ _0284_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__clkbuf_1
X_2137_ _0281_ RegFile.L\[1\] _0316_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1370_ RegFile.B\[6\] _0705_ _0710_ _0711_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2686_ clknet_2_3__leaf_clk _0162_ net64 VGND VGND VPWR VPWR PC.i_mem_addr\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1706_ _0645_ _1044_ _1045_ ByteBuffer.instr\[19\] VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_30_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1637_ RegFile.C\[6\] _0705_ _0707_ RegFile.L\[6\] VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1568_ _0883_ _0884_ _0909_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__a21o_1
X_1499_ RegFile.C\[3\] _0705_ _0707_ RegFile.L\[3\] _0840_ VGND VGND VPWR VPWR _0841_
+ sky130_fd_sc_hd__a221o_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__0517_ clknet_0__0517_ VGND VGND VPWR VPWR clknet_1_1__leaf__0517_
+ sky130_fd_sc_hd__clkbuf_16
X_2540_ _0577_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__clkbuf_1
X_1422_ RegFile.E\[5\] _0761_ _0763_ RegFile.H\[5\] VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__a22o_1
X_1284_ _0625_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__clkbuf_4
X_1353_ ByteBuffer.instr\[21\] VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2669_ net123 _0145_ net58 VGND VGND VPWR VPWR RegFile.B\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2435__34 clknet_1_0__leaf__0516_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__inv_2
X_1971_ _0736_ _0205_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__nor2_1
X_2450__48 clknet_1_1__leaf__0517_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__inv_2
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2523_ _0561_ _0562_ net46 VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__mux2_1
X_2385_ _0503_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkbuf_1
X_1405_ RegFile.H\[0\] _0680_ _0683_ RegFile.D\[0\] _0687_ VGND VGND VPWR VPWR _0747_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1336_ _0645_ ByteBuffer.instr\[22\] VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__nand2_4
Xinput1 cs VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_4
XFILLER_0_46_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2170_ _0816_ _1049_ _1166_ _1137_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__a22o_1
X_1954_ _1137_ _1142_ _1207_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1885_ RegFile.A\[6\] _1225_ _1203_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__mux2_1
X_2506_ _0548_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__clkbuf_1
X_2368_ _0428_ ALU.immediate\[14\] _0406_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2299_ _0223_ _0454_ _0457_ _0441_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__o211a_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1319_ _0619_ _0622_ _0624_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__and3b_1
XFILLER_0_2_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap52 _0685_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1670_ RegFile.D\[4\] _0683_ net52 RegFile.B\[4\] _0687_ VGND VGND VPWR VPWR _1012_
+ sky130_fd_sc_hd__a221o_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _1029_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2153_ _0334_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__inv_2
X_2084_ _0294_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__clkbuf_1
X_1937_ _0832_ _0912_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1868_ _1148_ _1207_ _1208_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__and3_1
X_1799_ ALU.flags_to_alu\[0\] _1059_ _1140_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1653_ _0729_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__inv_2
X_1722_ _1056_ _1063_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__nor2_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1584_ RegFile.E\[4\] _0789_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__or2_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _0382_ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__xnor2_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2136_ _0322_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
X_2067_ RegFile.C\[0\] _0283_ _0269_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1705_ _0670_ _1044_ _1046_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_5_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2685_ clknet_2_3__leaf_clk _0161_ net64 VGND VGND VPWR VPWR PC.i_mem_addr\[3\] sky130_fd_sc_hd__dfrtp_1
X_1567_ _0885_ _0896_ _0908_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__a21oi_1
X_1636_ _0971_ _0977_ _0629_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__a21o_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ RegFile.E\[3\] _0703_ _0699_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__o21a_1
X_2119_ _0313_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2456__54 clknet_1_0__leaf__0517_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__inv_2
XFILLER_0_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__0516_ clknet_0__0516_ VGND VGND VPWR VPWR clknet_1_1__leaf__0516_
+ sky130_fd_sc_hd__clkbuf_16
X_1421_ net57 _0650_ _0762_ _0638_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__o211a_2
X_1283_ ByteBuffer.instr\[23\] ByteBuffer.instr\[22\] VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__or2_1
X_1352_ _0670_ _0619_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2668_ net122 _0144_ net58 VGND VGND VPWR VPWR RegFile.B\[2\] sky130_fd_sc_hd__dfrtp_2
X_2599_ clknet_2_2__leaf_clk _0075_ net63 VGND VGND VPWR VPWR ALU.immediate\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1619_ RegFile.E\[6\] _0761_ _0771_ RegFile.B\[6\] VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_24_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1970_ _0204_ _1082_ _1043_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__mux2_1
X_2522_ PC.i_mem_addr\[4\] _0556_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1404_ _0740_ _0745_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__nand2_1
X_2384_ _0420_ ByteBuffer.instr\[21\] _0497_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__mux2_1
X_1335_ _0619_ _0640_ _0644_ _0632_ _0645_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__a221o_2
XFILLER_0_11_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput2 gpi[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1884_ _0655_ _1221_ _1224_ _0631_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__a22o_1
X_1953_ _0188_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2505_ PC.i_mem_addr\[1\] _0547_ _0542_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2298_ PC.i_mem_addr\[1\] _0451_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__or2_1
X_2367_ _0493_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1318_ ByteBuffer.instr\[20\] ByteBuffer.instr\[21\] VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap53 _0680_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_4
XFILLER_0_65_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _1049_ _0243_ _0397_ _0655_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__o211a_1
X_2152_ _0335_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2083_ RegFile.D\[2\] _0209_ _0288_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1867_ _1131_ _1147_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__or2_1
X_1936_ _1143_ _1145_ _1207_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1798_ _0908_ _0885_ _0896_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2472__6 clknet_1_0__leaf__0514_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__inv_2
XFILLER_0_30_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1721_ _1057_ _1060_ _1061_ _1062_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1652_ _0756_ _0990_ _0991_ _0993_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1583_ RegFile.C\[4\] _0793_ _0794_ RegFile.B\[4\] VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__a22o_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ _1239_ _0223_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__xnor2_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ _0279_ RegFile.L\[2\] _0316_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2066_ _0242_ _0261_ _0262_ net2 VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__a22o_1
X_1919_ _1257_ _1175_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2684_ clknet_2_3__leaf_clk _0160_ net64 VGND VGND VPWR VPWR PC.i_mem_addr\[2\] sky130_fd_sc_hd__dfrtp_1
X_1704_ _0645_ _1044_ _1045_ ByteBuffer.instr\[21\] VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1566_ _0907_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__buf_2
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1497_ RegFile.A\[3\] _0792_ _0704_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__or3_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1635_ _0972_ _0973_ _0975_ _0976_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__or4_1
X_2118_ _0209_ RegFile.H\[2\] net48 VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__mux2_1
X_2049_ RegFile.C\[6\] _0271_ _0269_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__mux2_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__0515_ clknet_0__0515_ VGND VGND VPWR VPWR clknet_1_1__leaf__0515_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1351_ _0664_ _0692_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__nor2_8
X_1420_ _0670_ _0757_ _0759_ _0650_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__a31oi_4
X_1282_ ByteBuffer.instr\[18\] VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1618_ _0947_ _0959_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_41_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2667_ net121 _0143_ net60 VGND VGND VPWR VPWR RegFile.B\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2598_ clknet_2_2__leaf_clk _0074_ net63 VGND VGND VPWR VPWR ALU.immediate\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1549_ RegFile.A\[0\] _0792_ _0704_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2521_ ALU.immediate\[4\] _0921_ _0519_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1403_ ALU.immediate\[9\] _0675_ _0693_ _0744_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__a22o_1
X_2383_ _0502_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
X_1334_ _0655_ _0675_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__nor2_4
XFILLER_0_11_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput3 gpi[1] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
XFILLER_0_61_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0__0517_ _0517_ VGND VGND VPWR VPWR clknet_0__0517_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1883_ _1092_ _1223_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1952_ RegFile.A\[3\] _0187_ _1203_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__mux2_1
X_2504_ _0545_ _0546_ net46 VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2366_ _0420_ ALU.immediate\[13\] _0406_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1317_ _0658_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__clkbuf_4
X_2297_ _0242_ _0454_ _0456_ _0441_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__o211a_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap54 _0708_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_4
XFILLER_0_65_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2220_ _1213_ _0990_ _0393_ _0395_ _0396_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__o2111a_1
X_2151_ ALU.flags_to_alu\[7\] _0327_ _0334_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__mux2_1
X_2082_ _0293_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1866_ _1151_ _1123_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__nor2_2
X_1935_ _1114_ _1272_ _1236_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__a21oi_1
X_1797_ _1138_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_31_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2349_ net134 MemControl.state\[1\] _0410_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1651_ _0992_ _0753_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__nor2_1
X_1720_ _0816_ _0831_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__or2b_1
XFILLER_0_38_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1582_ RegFile.H\[4\] _0784_ _0786_ RegFile.D\[4\] VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _0380_ _0381_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2065_ _0282_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__clkbuf_1
X_2134_ _0321_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1918_ _0780_ _0921_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__and2_1
X_1849_ ByteBuffer.instr\[20\] _1187_ _1190_ _0700_ _0645_ VGND VGND VPWR VPWR _1191_
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_39_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2683_ clknet_2_3__leaf_clk _0159_ net64 VGND VGND VPWR VPWR PC.i_mem_addr\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1703_ _0622_ _0624_ _0678_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__a21o_2
XFILLER_0_30_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1634_ RegFile.H\[6\] _0784_ _0817_ RegFile.L\[6\] VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__a22o_1
X_1565_ _0780_ _0903_ _0906_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__and3_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1496_ _0834_ _0836_ _0837_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__or3_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2048_ _1221_ _0261_ _0262_ net9 VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__a22o_1
X_2117_ _0312_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout58 net59 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_8
Xclkbuf_1_1__f__0514_ clknet_0__0514_ VGND VGND VPWR VPWR clknet_1_1__leaf__0514_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1281_ _0619_ _0622_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__nor2_2
X_1350_ _0666_ _0626_ _0673_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__o21a_2
XFILLER_0_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2597_ clknet_2_2__leaf_clk _0073_ net63 VGND VGND VPWR VPWR ALU.immediate\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1617_ _0955_ _0693_ _0958_ _0675_ ALU.immediate\[7\] VGND VGND VPWR VPWR _0959_
+ sky130_fd_sc_hd__a32o_2
X_2666_ net120 _0142_ net61 VGND VGND VPWR VPWR RegFile.B\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1479_ RegFile.H\[2\] _0784_ _0820_ _0711_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__a22o_1
X_1548_ RegFile.L\[0\] _0817_ _0889_ _0711_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2520_ _0560_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__clkbuf_1
X_1402_ _0741_ _0743_ _0630_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__and3b_2
X_2382_ _0421_ ByteBuffer.instr\[20\] _0497_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__mux2_1
X_1333_ _0664_ _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__nor2_8
Xinput4 gpi[23] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_2426__26 clknet_1_0__leaf__0515_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__inv_2
XFILLER_0_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2649_ net103 _0125_ net60 VGND VGND VPWR VPWR RegFile.E\[7\] sky130_fd_sc_hd__dfrtp_2
Xclkbuf_0__0516_ _0516_ VGND VGND VPWR VPWR clknet_0__0516_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1882_ _0718_ _1222_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__xor2_1
X_1951_ _0655_ _0182_ _0186_ _0631_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__a22o_2
XFILLER_0_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2503_ PC.i_mem_addr\[1\] PC.i_mem_addr\[0\] VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__xor2_1
X_2365_ _0492_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2296_ _0455_ _0454_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__nand2_1
X_1316_ ByteDecoder.state\[1\] ByteDecoder.state\[0\] VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap55 net56 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_4
XFILLER_0_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2150_ _0659_ _1201_ _0332_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__a31o_2
X_2081_ RegFile.D\[3\] _0187_ _0288_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1934_ _1113_ _1271_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__or2_1
X_1865_ _1120_ _1205_ _1131_ _1166_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_56_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1796_ _0883_ _0884_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2348_ _0484_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2279_ _0445_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2410__10 clknet_1_0__leaf__0515_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__inv_2
XFILLER_0_30_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1650_ _0749_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__inv_2
X_1581_ RegFile.A\[4\] _0792_ _0704_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__or3_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _1182_ _0203_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__xor2_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2064_ RegFile.C\[1\] _0281_ _0269_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__mux2_1
X_2133_ _0277_ RegFile.L\[3\] _0316_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1917_ _1254_ _1255_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1779_ _1098_ _1101_ _1120_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__or3_1
X_1848_ _1189_ _0666_ _0665_ ByteBuffer.instr\[21\] VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2682_ clknet_2_3__leaf_clk _0158_ net64 VGND VGND VPWR VPWR PC.i_mem_addr\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1702_ _0656_ _0700_ _0624_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__and3b_4
XFILLER_0_26_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1564_ _0904_ _0905_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__or2_1
X_1633_ RegFile.B\[6\] _0794_ _0974_ _0711_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ RegFile.C\[3\] _0793_ _0786_ RegFile.D\[3\] VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__a22o_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2047_ _0270_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__clkbuf_1
X_2116_ _0187_ RegFile.H\[3\] net48 VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout59 net64 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_8
XFILLER_0_67_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1280_ ByteBuffer.instr\[17\] VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2596_ clknet_2_2__leaf_clk _0072_ net63 VGND VGND VPWR VPWR ALU.immediate\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2665_ net119 _0141_ net60 VGND VGND VPWR VPWR RegFile.C\[7\] sky130_fd_sc_hd__dfrtp_1
X_1616_ RegFile.E\[7\] _0709_ _0957_ _0654_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__a211o_1
X_1547_ RegFile.E\[0\] _0789_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1478_ RegFile.E\[2\] _0789_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2381_ _0501_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
X_1401_ RegFile.B\[1\] _0705_ _0742_ _0711_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__a211o_1
Xinput5 gpi[2] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
X_1332_ _0666_ _0626_ _0673_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_52_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0__0515_ _0515_ VGND VGND VPWR VPWR clknet_0__0515_ sky130_fd_sc_hd__clkbuf_16
X_2579_ PC.i_mem_addr\[13\] _0609_ _0542_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2648_ net102 _0124_ net61 VGND VGND VPWR VPWR RegFile.E\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1950_ _0726_ _0184_ _0185_ _1092_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__o211a_2
X_1881_ _1025_ _1088_ _1043_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__mux2_1
X_2502_ _0867_ _0519_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__a21oi_1
X_2431__30 clknet_1_0__leaf__0516_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__inv_2
X_2364_ _0421_ ALU.immediate\[12\] _0406_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__mux2_1
X_1315_ ByteBuffer.instr\[21\] _0656_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2295_ PC.i_mem_addr\[0\] VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2080_ _0292_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__clkbuf_1
X_1933_ _1106_ _1112_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__nand2_1
X_1864_ _1103_ _1119_ _1124_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__o21ai_1
X_1795_ _1057_ _1060_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2347_ _1032_ _0476_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__and2_1
X_2278_ RegFile.A\[3\] net1 VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1580_ _0780_ _0921_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__nand2_2
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _0242_ _0379_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__xnor2_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2132_ _0320_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2063_ _0223_ _0261_ _0262_ net3 VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__a22o_2
XFILLER_0_21_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1916_ _1151_ _1048_ _1159_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1847_ _0668_ _0696_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__nor2_1
X_1778_ _1103_ _1119_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1701_ _0678_ _1039_ _1042_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_26_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2681_ net71 _0157_ net59 VGND VGND VPWR VPWR RegFile.A\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1563_ RegFile.L\[0\] _0680_ _0687_ ALU.flags_to_alu\[0\] VGND VGND VPWR VPWR _0905_
+ sky130_fd_sc_hd__a22o_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1494_ RegFile.H\[3\] _0784_ _0835_ _0711_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__a22o_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1632_ RegFile.E\[6\] _0789_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__or2_1
X_2115_ _0311_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2046_ RegFile.C\[7\] _0263_ _0269_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2664_ net118 _0140_ net59 VGND VGND VPWR VPWR RegFile.C\[6\] sky130_fd_sc_hd__dfrtp_1
X_2595_ clknet_2_2__leaf_clk _0071_ net63 VGND VGND VPWR VPWR ALU.immediate\[9\] sky130_fd_sc_hd__dfrtp_1
X_1546_ RegFile.H\[0\] _0784_ _0788_ ALU.flags_to_alu\[0\] _0887_ VGND VGND VPWR VPWR
+ _0888_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1615_ ALU.flags_to_alu\[7\] _0711_ _0707_ RegFile.L\[7\] _0956_ VGND VGND VPWR VPWR
+ _0957_ sky130_fd_sc_hd__a221o_1
X_1477_ ALU.flags_to_alu\[2\] _0788_ _0817_ RegFile.L\[2\] _0818_ VGND VGND VPWR VPWR
+ _0819_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2029_ _0256_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__clkbuf_1
X_2452__50 clknet_1_0__leaf__0517_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__inv_2
XFILLER_0_13_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2380_ _0490_ ByteBuffer.instr\[19\] _0497_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__mux2_1
X_1331_ _0669_ _0671_ _0672_ _0659_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__o211a_1
X_1400_ RegFile.H\[1\] _0707_ _0709_ RegFile.D\[1\] VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput6 gpi[3] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0__0514_ _0514_ VGND VGND VPWR VPWR clknet_0__0514_ sky130_fd_sc_hd__clkbuf_16
X_2647_ net101 _0123_ net61 VGND VGND VPWR VPWR RegFile.E\[5\] sky130_fd_sc_hd__dfrtp_1
X_2578_ _0540_ _0607_ _0608_ _0585_ ALU.immediate\[13\] VGND VGND VPWR VPWR _0609_
+ sky130_fd_sc_hd__a32o_1
X_1529_ RegFile.H\[1\] _0784_ _0788_ ALU.flags_to_alu\[1\] VGND VGND VPWR VPWR _0871_
+ sky130_fd_sc_hd__a22oi_1
X_2417__17 clknet_1_1__leaf__0515_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__inv_2
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1880_ _1220_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__buf_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2501_ ALU.immediate\[1\] _0519_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2363_ _0491_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
X_2294_ _0453_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__buf_4
X_1314_ _0619_ _0622_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap57 _0646_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_2
XFILLER_0_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1863_ _1204_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkbuf_1
X_1932_ _1270_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1794_ _1127_ _1135_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__nand2_2
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2346_ _0483_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2277_ _0444_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _1221_ _1265_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__xor2_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2062_ _0280_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__clkbuf_1
X_2131_ _0275_ RegFile.L\[4\] _0316_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1777_ _0806_ _0936_ _1118_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__o21bai_1
X_1915_ _1151_ _1173_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__and2_1
X_1846_ _0700_ _1186_ _1187_ ByteBuffer.instr\[19\] _0645_ VGND VGND VPWR VPWR _1188_
+ sky130_fd_sc_hd__a221o_2
X_2329_ _0441_ _0473_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1700_ ByteBuffer.instr\[20\] _0645_ _0672_ _1041_ _0648_ VGND VGND VPWR VPWR _1042_
+ sky130_fd_sc_hd__a221o_1
X_2680_ net70 _0156_ net59 VGND VGND VPWR VPWR RegFile.A\[6\] sky130_fd_sc_hd__dfrtp_4
X_1631_ RegFile.C\[6\] _0793_ _0786_ RegFile.D\[6\] VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1562_ RegFile.E\[0\] _0683_ _0685_ RegFile.C\[0\] _0654_ VGND VGND VPWR VPWR _0904_
+ sky130_fd_sc_hd__a221o_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ RegFile.E\[3\] _0789_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__or2_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2114_ _1269_ RegFile.H\[4\] net48 VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__mux2_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2045_ _0655_ _0264_ _0267_ _0268_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__o211a_4
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1829_ _1151_ _1122_ _1159_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__or3b_1
XFILLER_0_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2438__37 clknet_1_1__leaf__0516_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__inv_2
X_2594_ clknet_2_2__leaf_clk _0070_ net63 VGND VGND VPWR VPWR ALU.immediate\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1614_ RegFile.C\[7\] net54 net56 VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__and3_1
X_2663_ net117 _0139_ net61 VGND VGND VPWR VPWR RegFile.C\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_22_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1545_ RegFile.C\[0\] _0792_ _0699_ net55 VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1476_ RegFile.B\[2\] _0785_ _0708_ net56 VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__and4_1
XFILLER_0_49_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2028_ _0187_ RegFile.B\[3\] _0251_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1330_ _0645_ ByteBuffer.instr\[22\] VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_52_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 gpi[4] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_54_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2577_ PC.i_mem_addr\[12\] _0597_ PC.i_mem_addr\[13\] VGND VGND VPWR VPWR _0608_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2646_ net100 _0122_ net60 VGND VGND VPWR VPWR RegFile.E\[4\] sky130_fd_sc_hd__dfrtp_2
X_1528_ RegFile.C\[1\] _0793_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__nand2_1
X_1459_ ALU.flags_to_alu\[5\] _0711_ _0799_ _0800_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2500_ _0543_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2362_ _0490_ ALU.immediate\[11\] _0406_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__mux2_1
X_2293_ _0450_ _0655_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1313_ _0654_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2629_ net83 _0105_ net58 VGND VGND VPWR VPWR RegFile.L\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap47 _0333_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput10 gpi[7] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
X_1793_ _0935_ _0936_ _1064_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1862_ RegFile.A\[7\] _1184_ _1203_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__mux2_1
X_1931_ RegFile.A\[4\] _1269_ _1203_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2345_ _0713_ _0476_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__and2_1
X_2276_ RegFile.A\[2\] net1 VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2061_ RegFile.C\[2\] _0279_ _0269_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__mux2_1
X_2130_ _0319_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1914_ _1165_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1776_ _1105_ _1116_ _1117_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1845_ _0700_ _0641_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__nand2_1
X_2328_ _0450_ _0325_ _0454_ PC.i_mem_addr\[15\] VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2259_ net8 _0419_ _0425_ net7 VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__and4bb_1
X_2459__57 clknet_1_1__leaf__0517_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__inv_2
XFILLER_0_62_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1630_ ALU.flags_to_alu\[6\] _0788_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__and2_1
X_1561_ RegFile.A\[0\] net51 _0898_ _0902_ _0629_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__a2111o_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ ALU.flags_to_alu\[3\] _0788_ _0817_ RegFile.L\[3\] _0833_ VGND VGND VPWR VPWR
+ _0834_ sky130_fd_sc_hd__a221o_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2113_ _0310_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
X_2044_ _0655_ _1193_ _1201_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_44_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1759_ _1100_ _0805_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__nor2_1
X_1828_ _1069_ _1164_ _1167_ _1169_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2593_ clknet_2_1__leaf_clk _0069_ net62 VGND VGND VPWR VPWR ByteDecoder.num_bytes\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2662_ net116 _0138_ net60 VGND VGND VPWR VPWR RegFile.C\[4\] sky130_fd_sc_hd__dfrtp_2
X_1613_ _0948_ _0954_ _0629_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__a21o_1
X_1544_ RegFile.D\[0\] _0786_ _0794_ RegFile.B\[0\] VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1475_ _0789_ _0699_ net55 VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__and3_2
X_2027_ _0255_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 gpi[5] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_0_54_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2576_ _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__inv_2
X_1527_ ALU.immediate\[1\] _0675_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__nand2_1
X_2645_ net99 _0121_ net58 VGND VGND VPWR VPWR RegFile.E\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1389_ RegFile.B\[2\] _0705_ _0730_ _0711_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__a211o_1
X_1458_ RegFile.E\[5\] _0699_ net55 _0654_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2361_ net6 _0416_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1312_ _0653_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__clkbuf_8
X_2292_ _0452_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2422__22 clknet_1_0__leaf__0515_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__inv_2
X_2559_ PC.i_mem_addr\[10\] _0588_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__nand2_1
X_2628_ net82 _0104_ net58 VGND VGND VPWR VPWR RegFile.L\[2\] sky130_fd_sc_hd__dfrtp_2
Xmax_cap48 _0307_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_4
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1930_ _0655_ _1265_ _1268_ _0631_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__a22o_2
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1792_ _1132_ _1133_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__xnor2_2
Xinput11 nrst VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1861_ _1192_ _1202_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__nor2_8
X_2344_ _0482_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2275_ _0443_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2060_ _0203_ _0261_ _0262_ net5 VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1913_ _0938_ _1251_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1775_ _0806_ _0936_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1844_ ByteBuffer.instr\[20\] _0665_ _1185_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__a21o_1
X_2258_ _0418_ _0424_ _0429_ _0430_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__o211ai_1
X_2327_ _1224_ _0454_ _0472_ _0441_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__o211a_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2189_ _1069_ _1092_ _1093_ _1131_ _0367_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1560_ RegFile.E\[0\] _0761_ _0899_ _0900_ _0901_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__a2111o_1
X_2112_ _1247_ RegFile.H\[5\] net48 VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__mux2_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1491_ RegFile.B\[3\] _0785_ _0708_ net56 VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__and4_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2043_ _0630_ _0266_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__or2_2
X_1827_ _1075_ _1168_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1758_ _1099_ _1095_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__and2_1
X_1689_ RegFile.B\[7\] _0705_ _1030_ _0711_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2661_ net115 _0137_ net59 VGND VGND VPWR VPWR RegFile.C\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2592_ clknet_2_2__leaf_clk _0068_ net63 VGND VGND VPWR VPWR ByteDecoder.num_bytes\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1543_ ALU.immediate\[0\] _0664_ _0692_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__o21ai_4
X_1474_ _0780_ _0815_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__nand2_8
XFILLER_0_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1612_ _0949_ _0950_ _0952_ _0953_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2026_ _1269_ RegFile.B\[4\] _0251_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__mux2_1
X_2429__28 clknet_1_0__leaf__0516_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__inv_2
XFILLER_0_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2443__42 clknet_1_0__leaf__0516_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__inv_2
XFILLER_0_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput9 gpi[6] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2644_ net98 _0120_ net58 VGND VGND VPWR VPWR RegFile.E\[2\] sky130_fd_sc_hd__dfrtp_1
X_2575_ PC.i_mem_addr\[12\] PC.i_mem_addr\[13\] _0597_ VGND VGND VPWR VPWR _0606_
+ sky130_fd_sc_hd__and3_1
X_1526_ _0675_ _0867_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1457_ RegFile.C\[5\] _0705_ _0707_ RegFile.L\[5\] VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__a22o_1
X_1388_ RegFile.H\[2\] _0707_ _0709_ RegFile.D\[2\] VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2009_ _1166_ _0231_ _0235_ _0241_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__a211o_2
XFILLER_0_37_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2360_ _0489_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1311_ _0623_ _0628_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__or2_1
X_2291_ _0441_ _0451_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2627_ net81 _0103_ net60 VGND VGND VPWR VPWR RegFile.L\[1\] sky130_fd_sc_hd__dfrtp_2
X_2558_ _0592_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__clkbuf_1
X_2489_ _0678_ _0636_ _0526_ _0530_ _0532_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__o41a_1
X_1509_ ALU.flags_to_alu\[3\] _0687_ _0683_ RegFile.E\[3\] _0654_ VGND VGND VPWR VPWR
+ _0851_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap49 _1043_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_4
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1860_ _0630_ _1193_ _1201_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__o21bai_4
X_1791_ _1072_ _1127_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2343_ _1006_ _0476_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2274_ RegFile.A\[1\] _0441_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1989_ _1142_ _1207_ _0212_ _0222_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__a31o_2
XFILLER_0_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1912_ _0937_ _1250_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1843_ _0642_ _0666_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f__0517_ clknet_0__0517_ VGND VGND VPWR VPWR clknet_1_0__leaf__0517_
+ sky130_fd_sc_hd__clkbuf_16
X_1774_ _1114_ _1115_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2257_ ByteDecoder.state\[1\] ByteDecoder.state\[0\] VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__nor2_1
X_2326_ PC.i_mem_addr\[14\] _0451_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2188_ _1050_ _1212_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1490_ _0816_ _0831_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 ByteDecoder.num_bytes\[1\] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlygate4sd3_1
X_2111_ _0309_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2042_ _0265_ _1191_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2464__62 clknet_1_0__leaf__0517_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__inv_2
X_1826_ net49 _1122_ _1159_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__or3b_4
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1757_ _0970_ _0982_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1688_ RegFile.H\[7\] _0707_ _0709_ RegFile.D\[7\] VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__a22o_1
X_2309_ _1221_ _0454_ _0462_ _0441_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__o211a_1
XFILLER_0_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1611_ RegFile.H\[7\] _0784_ _0817_ RegFile.L\[7\] VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__a22o_1
X_2660_ net114 _0136_ net58 VGND VGND VPWR VPWR RegFile.C\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2591_ clknet_2_1__leaf_clk _0067_ net62 VGND VGND VPWR VPWR ByteDecoder.num_bytes\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1542_ _0675_ _0867_ _0869_ _0880_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_1_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1473_ _0629_ _0812_ _0813_ _0814_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__o22a_2
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2025_ _0254_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__clkbuf_1
X_1809_ _1150_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2574_ _0605_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__clkbuf_1
X_2643_ net97 _0119_ net60 VGND VGND VPWR VPWR RegFile.E\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1525_ _0629_ _0862_ _0863_ _0865_ _0866_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__o32a_4
X_1387_ RegFile.A\[2\] _0652_ _0676_ _0728_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__o211a_2
X_1456_ _0787_ _0791_ _0796_ _0797_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__o31a_1
X_2008_ _0236_ _0237_ _0240_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2290_ _0450_ _0655_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__nor2_8
X_1310_ _0651_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__buf_4
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2557_ PC.i_mem_addr\[9\] _0591_ _0542_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2626_ net80 _0102_ net61 VGND VGND VPWR VPWR RegFile.L\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2488_ ByteBuffer.instr\[20\] _0342_ _0531_ _0636_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__or4b_1
X_1439_ _0629_ _0775_ _0778_ _0780_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__o211ai_4
X_1508_ _0847_ _0848_ _0849_ _0774_ RegFile.A\[3\] VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__o32a_1
XFILLER_0_33_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2413__13 clknet_1_1__leaf__0515_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__inv_2
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1790_ _0806_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2342_ _0481_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
X_2273_ _0442_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
X_1988_ _1166_ _0211_ _0214_ _1124_ _0221_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__a221o_1
X_2609_ clknet_2_0__leaf_clk _0085_ net62 VGND VGND VPWR VPWR ByteBuffer.instr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1773_ _0937_ _0913_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__xnor2_1
X_1911_ _0832_ _0856_ _0912_ _0913_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__o31a_1
X_1842_ _0631_ _1094_ _1183_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_1_0__f__0516_ clknet_0__0516_ VGND VGND VPWR VPWR clknet_1_0__leaf__0516_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2325_ _1246_ _0454_ _0471_ _0441_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__o211a_1
X_2187_ _1066_ _1092_ _1158_ _0346_ _1181_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__o221a_1
X_2256_ _0426_ _0427_ _0417_ _0428_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2 FSM.next_state\[0\] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dlygate4sd3_1
X_2041_ _1188_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__inv_2
X_2110_ _1225_ RegFile.H\[6\] net48 VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__mux2_1
X_1756_ _1096_ _1097_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1825_ ALU.flags_to_alu\[0\] _1151_ _1165_ _1166_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2308_ PC.i_mem_addr\[6\] _0451_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__or2_1
X_1687_ RegFile.A\[7\] _0652_ _1028_ _0676_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2239_ ByteDecoder.state\[1\] ByteDecoder.num_bytes\[2\] ByteDecoder.num_bytes\[3\]
+ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__nor3_1
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2468__2 clknet_1_0__leaf__0514_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__inv_2
X_2590_ clknet_2_0__leaf_clk _0066_ net62 VGND VGND VPWR VPWR MemControl.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1610_ RegFile.B\[7\] _0794_ _0951_ _0711_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1541_ _0675_ _0867_ _0880_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__or3_1
X_1472_ RegFile.L\[2\] net53 net52 RegFile.C\[2\] VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2024_ _1247_ RegFile.B\[5\] _0251_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1739_ _0740_ _0745_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__and2b_1
X_1808_ _0678_ _1039_ _1042_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2434__33 clknet_1_1__leaf__0516_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__inv_2
X_2573_ PC.i_mem_addr\[12\] _0604_ _0542_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1524_ ALU.flags_to_alu\[1\] _0652_ _0629_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2642_ net96 _0118_ net61 VGND VGND VPWR VPWR RegFile.E\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1386_ RegFile.H\[2\] net53 _0727_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__a21o_1
X_1455_ RegFile.A\[5\] _0792_ _0704_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__or3_1
X_2007_ _1140_ _0238_ _0239_ net49 VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__a22o_1
X_2408__8 clknet_1_1__leaf__0515_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__inv_2
XFILLER_0_45_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2556_ net46 _0589_ _0590_ _0585_ ALU.immediate\[9\] VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__a32o_1
X_2487_ _0678_ _0524_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__or2_1
X_2625_ net79 _0101_ net61 VGND VGND VPWR VPWR ALU.flags_to_alu\[7\] sky130_fd_sc_hd__dfrtp_2
X_1507_ ALU.flags_to_alu\[3\] _0765_ _0763_ RegFile.H\[3\] VGND VGND VPWR VPWR _0849_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1438_ _0779_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1369_ net54 net55 VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__nor2_8
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2341_ _1017_ _0476_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__and2_1
X_2272_ RegFile.A\[0\] _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1987_ _0816_ _1253_ _0215_ _0220_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__o211ai_1
X_2539_ PC.i_mem_addr\[6\] _0576_ _0542_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__mux2_1
X_2608_ clknet_2_0__leaf_clk _0084_ net59 VGND VGND VPWR VPWR ByteBuffer.instr\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1910_ _1136_ _1146_ _1207_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_52_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1772_ _1106_ _1112_ _1113_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__a21bo_1
X_1841_ _0655_ _1182_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__0515_ clknet_0__0515_ VGND VGND VPWR VPWR clknet_1_0__leaf__0515_
+ sky130_fd_sc_hd__clkbuf_16
X_2324_ PC.i_mem_addr\[13\] _0451_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__or2_1
X_2186_ _0362_ _0363_ _0361_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__o21ai_1
X_2255_ net9 _0416_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3 ByteDecoder.num_bytes\[2\] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ _1188_ _1191_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__nor2_1
X_1824_ _1151_ _1049_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__nor2_2
X_1755_ _0960_ _1095_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1686_ RegFile.H\[7\] net53 _1027_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2307_ _1239_ _0454_ _0461_ _0441_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__o211a_1
X_2238_ _0409_ _0410_ _0411_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__or3_2
X_2169_ _1093_ _1136_ _0346_ _1252_ _0347_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__o221a_1
X_2455__53 clknet_1_1__leaf__0517_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__inv_2
XFILLER_0_50_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1540_ _0868_ _0881_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1471_ ALU.flags_to_alu\[2\] _0687_ _0683_ RegFile.E\[2\] _0654_ VGND VGND VPWR VPWR
+ _0813_ sky130_fd_sc_hd__a221o_1
X_2023_ _0253_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__clkbuf_1
X_1807_ _1130_ _1148_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1738_ _1055_ _1079_ _0754_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__a21bo_1
X_1669_ _1009_ _1010_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2470__4 clknet_1_1__leaf__0514_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__inv_2
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2572_ _0540_ _0602_ _0603_ _0585_ ALU.immediate\[12\] VGND VGND VPWR VPWR _0604_
+ sky130_fd_sc_hd__a32o_1
X_2641_ net95 _0117_ net60 VGND VGND VPWR VPWR RegFile.H\[7\] sky130_fd_sc_hd__dfrtp_2
X_1523_ RegFile.L\[1\] net53 _0864_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__a21oi_1
X_1454_ RegFile.C\[5\] _0793_ _0794_ RegFile.B\[5\] _0795_ VGND VGND VPWR VPWR _0796_
+ sky130_fd_sc_hd__a221o_1
X_1385_ RegFile.D\[2\] _0683_ net52 RegFile.B\[2\] _0687_ VGND VGND VPWR VPWR _0727_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2006_ _0947_ _1214_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__nor2_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2624_ net78 _0100_ net60 VGND VGND VPWR VPWR ALU.flags_to_alu\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2555_ PC.i_mem_addr\[9\] _0582_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2486_ _0326_ _0525_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__xnor2_1
X_1437_ _0664_ _0674_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1506_ RegFile.D\[3\] _0767_ _0771_ RegFile.B\[3\] VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__a22o_1
X_1299_ _0619_ _0622_ _0624_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__a21bo_1
X_1368_ RegFile.H\[6\] _0707_ _0709_ RegFile.D\[6\] VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2340_ _0480_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
X_2271_ net1 VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__buf_8
XFILLER_0_59_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1986_ _1213_ _0217_ _0219_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2607_ clknet_2_1__leaf_clk _0083_ net62 VGND VGND VPWR VPWR ByteBuffer.instr\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2538_ _0572_ _0575_ net46 VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1840_ _1126_ _1152_ _1180_ _1181_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__o31a_2
X_1771_ _1104_ _0856_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__nor2_2
XFILLER_0_37_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__0514_ clknet_0__0514_ VGND VGND VPWR VPWR clknet_1_0__leaf__0514_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2323_ _1268_ _0454_ _0470_ _0441_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__o211a_1
X_2254_ net2 _0419_ _0420_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__or3b_1
X_2185_ _0361_ _0362_ _0363_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1969_ _0746_ _0994_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold4 ByteBuffer.counter\[0\] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1823_ _1048_ _1163_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1754_ _0960_ _1095_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1685_ RegFile.D\[7\] _0683_ net52 RegFile.B\[7\] _0687_ VGND VGND VPWR VPWR _1027_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2306_ PC.i_mem_addr\[5\] _0451_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__or2_1
X_2237_ MemControl.state\[2\] MemControl.state\[1\] MemControl.state\[0\] VGND VGND
+ VPWR VPWR _0411_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2168_ _1257_ _1049_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2099_ _0302_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1470_ _0809_ _0810_ _0811_ _0774_ RegFile.A\[2\] VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__o32a_1
X_2022_ _1225_ RegFile.B\[6\] _0251_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__mux2_1
X_1806_ _1131_ _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1668_ _1003_ _1007_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__nor2_1
X_1737_ _0960_ _0983_ _1064_ _1065_ _1078_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__a41o_1
XFILLER_0_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1599_ ALU.flags_to_alu\[7\] _0765_ _0767_ RegFile.D\[7\] _0940_ VGND VGND VPWR VPWR
+ _0941_ sky130_fd_sc_hd__a221o_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2640_ net94 _0116_ net59 VGND VGND VPWR VPWR RegFile.H\[6\] sky130_fd_sc_hd__dfrtp_2
X_2571_ PC.i_mem_addr\[12\] _0597_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__or2_1
X_1522_ RegFile.E\[1\] _0683_ net52 RegFile.C\[1\] _0687_ VGND VGND VPWR VPWR _0864_
+ sky130_fd_sc_hd__a221o_1
X_1453_ RegFile.L\[5\] _0789_ _0699_ net55 VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__and4_1
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1384_ _0721_ _0725_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__xnor2_2
X_2005_ _1059_ _1161_ _1255_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2554_ _0588_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2623_ net77 _0099_ net60 VGND VGND VPWR VPWR ALU.flags_to_alu\[5\] sky130_fd_sc_hd__dfrtp_2
X_2485_ _0524_ _0525_ _0528_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1505_ RegFile.E\[3\] _0761_ _0845_ _0846_ net50 VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_10_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1436_ _0776_ _0777_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__or2_2
X_1367_ net54 _0703_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__nor2_4
XFILLER_0_37_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1298_ ByteBuffer.instr\[20\] _0639_ _0632_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_65_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2270_ MemControl.state\[0\] _0439_ _0440_ net135 VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1985_ _0196_ _1254_ _1164_ _0908_ _0218_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__a221o_1
X_2537_ _0573_ _0574_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__nor2_1
X_2606_ clknet_2_0__leaf_clk _0082_ net62 VGND VGND VPWR VPWR ByteBuffer.instr\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_30_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2399_ _0510_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
X_1419_ _0684_ _0677_ _0679_ _0760_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__and4_4
XFILLER_0_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1770_ _1107_ _1111_ _0832_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2322_ PC.i_mem_addr\[12\] _0451_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__or2_1
X_2184_ _1092_ _1223_ _0227_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__and3_1
X_2253_ net3 net5 net6 _0425_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__or4b_1
XFILLER_0_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1899_ _1147_ _1228_ _1234_ _1238_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1968_ _1166_ _1137_ _0190_ _0202_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold5 ByteDecoder.num_bytes\[3\] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1753_ _0970_ _0982_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1822_ _1122_ _1163_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__nor2_2
XFILLER_0_37_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1684_ _0718_ _1025_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2305_ _1265_ _0454_ _0460_ _0441_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__o211a_1
X_2167_ _1151_ _1092_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__nand2_2
X_2236_ _0670_ _0659_ _0662_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__and3_2
XFILLER_0_67_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2098_ RegFile.E\[3\] _0277_ _0297_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2021_ _0252_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1805_ _1134_ _1136_ _1146_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__nor3_2
X_1736_ _1067_ _1077_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__nand2_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1667_ _1008_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1598_ RegFile.C\[7\] _0638_ _0681_ _0760_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__and4_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ _0908_ _1165_ _0239_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2570_ PC.i_mem_addr\[12\] _0597_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1383_ ALU.immediate\[11\] _0675_ _0693_ _0724_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__a22o_2
X_1521_ RegFile.A\[1\] _0774_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__nor2_1
X_1452_ _0785_ net54 net55 VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__and3_2
XFILLER_0_22_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2004_ _0908_ _1175_ _1165_ _0196_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2425__25 clknet_1_1__leaf__0515_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__inv_2
X_2440__39 clknet_1_1__leaf__0516_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__inv_2
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1719_ _0855_ _0844_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__nand2_1
X_2699_ clknet_2_1__leaf_clk _0001_ net62 VGND VGND VPWR VPWR MemControl.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2553_ PC.i_mem_addr\[9\] _0582_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1504_ RegFile.L\[3\] _0638_ _0681_ _0762_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2622_ net76 _0098_ net60 VGND VGND VPWR VPWR ALU.flags_to_alu\[4\] sky130_fd_sc_hd__dfrtp_1
X_2484_ _0403_ _0527_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__nand2_1
X_1366_ _0694_ _0698_ _0648_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__a21oi_2
X_1435_ RegFile.L\[5\] _0680_ _0687_ ALU.flags_to_alu\[5\] VGND VGND VPWR VPWR _0777_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1297_ _0624_ ByteBuffer.instr\[17\] VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1984_ _0196_ _1175_ _1162_ _1139_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2536_ PC.i_mem_addr\[6\] _0567_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__nor2_1
X_2605_ clknet_2_0__leaf_clk _0081_ net62 VGND VGND VPWR VPWR ByteBuffer.instr\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1349_ _0690_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2398_ _0421_ ALU.immediate\[4\] _0408_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__mux2_1
X_1418_ _0670_ _0757_ _0759_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__and3_4
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2321_ _0186_ _0454_ _0469_ _0441_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__o211a_1
XFILLER_0_12_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2183_ _1092_ _1223_ _0227_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__a21oi_1
X_2252_ net2 _0416_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1898_ _1049_ _1235_ _1237_ _1118_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1967_ _0191_ _0192_ _0201_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2519_ PC.i_mem_addr\[3\] _0559_ _0542_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold6 MemControl.state\[2\] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1683_ _1000_ _1011_ _1022_ _1024_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__o31a_1
X_1752_ _1038_ _1051_ _1090_ _1093_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_44_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1821_ ByteBuffer.instr\[21\] _0645_ _1044_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__or3b_2
XFILLER_0_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2304_ PC.i_mem_addr\[4\] _0451_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__or2_1
X_2166_ _1094_ _0186_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__xor2_1
X_2235_ MemControl.state\[0\] _0260_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__and2_1
X_2097_ _0301_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2446__45 clknet_1_0__leaf__0516_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__inv_2
X_2461__59 clknet_1_0__leaf__0517_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__inv_2
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2020_ _1184_ RegFile.B\[7\] _0251_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1666_ _1003_ _1007_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__nand2_1
X_1804_ _1143_ _1145_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__nand2_2
X_1735_ _1070_ _1074_ _1075_ _1076_ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1597_ RegFile.E\[7\] _0761_ _0771_ RegFile.B\[7\] VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__a22o_1
X_2218_ ALU.flags_to_alu\[0\] _1151_ _1122_ _0394_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__a31o_1
X_2149_ _1192_ _0630_ _1202_ _0286_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1520_ _0859_ _0860_ _0861_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__nor3_1
XFILLER_0_10_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1382_ RegFile.A\[3\] _0704_ _0723_ _0630_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__o211a_1
X_1451_ _0792_ _0699_ net55 VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__and3_2
X_2003_ ALU.flags_to_alu\[0\] _1151_ _1164_ _1254_ _0908_ VGND VGND VPWR VPWR _0236_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_60_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1649_ _0740_ _0745_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__nor2_1
X_2698_ clknet_2_0__leaf_clk net136 net62 VGND VGND VPWR VPWR MemControl.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_1718_ _1058_ _1059_ _0883_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2552_ _0587_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2483_ _0678_ _0526_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1503_ RegFile.C\[3\] _0638_ _0681_ _0760_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__and4_1
X_2621_ net75 _0097_ net58 VGND VGND VPWR VPWR ALU.flags_to_alu\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1296_ _0622_ _0632_ _0634_ _0637_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__a2bb2o_4
X_1365_ _0699_ net56 VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__nor2_8
X_1434_ RegFile.E\[5\] _0683_ _0685_ RegFile.C\[5\] _0654_ VGND VGND VPWR VPWR _0776_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1983_ _0910_ _0216_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__nand2_1
X_2604_ clknet_2_0__leaf_clk _0080_ net59 VGND VGND VPWR VPWR ByteBuffer.instr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_2535_ PC.i_mem_addr\[6\] _0567_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__and2_1
X_1417_ _0700_ _0758_ _0647_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__a21o_1
X_1279_ _0619_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__or2_2
X_2397_ _0509_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
X_1348_ RegFile.A\[6\] _0652_ _0676_ _0689_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2320_ PC.i_mem_addr\[11\] _0451_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__or2_1
X_2251_ _0419_ _0420_ _0421_ _0423_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2182_ _1246_ _1268_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__xnor2_1
X_1966_ _1213_ _0194_ _0200_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1897_ _1117_ _1105_ _1116_ _1236_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__a31o_1
X_2518_ _0555_ _0558_ net46 VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2473__7 clknet_1_1__leaf__0514_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__inv_2
XFILLER_0_61_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold7 MemControl.state\[1\] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dlygate4sd3_1
X_1820_ net49 _1160_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1682_ _1023_ _1007_ _1011_ _1020_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__o22a_1
X_1751_ net49 _1092_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__nand2_4
XFILLER_0_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2303_ _0182_ _0454_ _0459_ _0441_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__o211a_1
X_2234_ _0406_ _0408_ VGND VGND VPWR VPWR ByteBuffer.next_counter\[1\] sky130_fd_sc_hd__nand2_1
XFILLER_0_29_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2165_ _0277_ net47 _0336_ net141 VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__a22o_1
X_2096_ RegFile.E\[4\] _0275_ _0297_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__mux2_1
X_1949_ _0726_ _0184_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1803_ _1144_ _1113_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1665_ ALU.immediate\[13\] _0675_ _0693_ _1006_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__a22o_1
X_1596_ _0832_ _0856_ _0912_ _0913_ _0937_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__o311a_1
X_1734_ _1069_ _0982_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ ALU.flags_to_alu\[0\] _1151_ _1173_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2148_ _0331_ _0626_ _0645_ _1197_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__a2bb2o_1
X_2079_ RegFile.D\[4\] _1269_ _0288_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1450_ _0648_ _0783_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__nor2_2
X_1381_ RegFile.B\[3\] _0705_ _0722_ _0711_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__a211o_1
X_2002_ _0231_ _0232_ _0233_ _1162_ _0234_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__o32a_1
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1648_ _0806_ _0938_ _0984_ _0989_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__a31o_1
X_2697_ clknet_2_1__leaf_clk _0173_ net62 VGND VGND VPWR VPWR PC.i_mem_addr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1717_ _0885_ _0896_ _0908_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__a21bo_2
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1579_ _0629_ _0918_ _0919_ _0920_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__o22a_2
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2416__16 clknet_1_1__leaf__0515_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__inv_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2620_ net74 _0096_ net59 VGND VGND VPWR VPWR ALU.flags_to_alu\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2551_ PC.i_mem_addr\[8\] _0586_ _0542_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1502_ ALU.immediate\[3\] _0674_ _0843_ _0830_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__o211a_2
X_2482_ ByteBuffer.instr\[20\] _0639_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1433_ _0764_ _0769_ _0773_ _0774_ RegFile.A\[5\] VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__o32a_2
XFILLER_0_37_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1295_ _0626_ _0635_ _0636_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__and3b_1
X_1364_ _0622_ _0701_ _0702_ _0626_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1982_ _1139_ _0909_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2534_ ALU.immediate\[6\] _0969_ _0519_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__mux2_1
X_2603_ clknet_2_0__leaf_clk _0079_ net59 VGND VGND VPWR VPWR ByteBuffer.instr\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_2396_ _0490_ ALU.immediate\[3\] _0408_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__mux2_1
X_1416_ _0619_ _0622_ ByteBuffer.instr\[21\] VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__a21bo_1
X_1347_ RegFile.H\[6\] net53 _0688_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1278_ ByteBuffer.instr\[17\] VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2250_ _0419_ _0422_ net2 VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2181_ _0345_ _0359_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1965_ _0195_ _0197_ _0198_ _0199_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__or4b_1
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2517_ _0556_ _0557_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__nor2_1
X_1896_ net49 _1123_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2379_ _0500_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold8 _0000_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1750_ _1091_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__buf_6
XFILLER_0_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1681_ _1003_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2302_ PC.i_mem_addr\[3\] _0451_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__or2_1
X_2233_ _0407_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__clkbuf_4
X_2164_ _0275_ net47 _0336_ net138 VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2095_ _0300_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__clkbuf_1
X_1879_ _1206_ _1209_ _1219_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__or3b_1
X_1948_ _0997_ _0183_ _1043_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_2437__36 clknet_1_1__leaf__0516_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__inv_2
XFILLER_0_15_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1733_ _1066_ _0959_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__nor2_1
X_1802_ _1057_ _1060_ _1062_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__o21ai_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1595_ _0935_ _0936_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__nor2_2
XFILLER_0_40_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1664_ RegFile.A\[5\] _0704_ _1005_ _0630_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__o211a_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _1149_ _1079_ _1207_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__o21ai_1
X_2147_ _0647_ _0328_ _0330_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2078_ _0291_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1380_ RegFile.H\[3\] _0707_ _0709_ RegFile.D\[3\] VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__a22o_1
X_2001_ _1059_ _1123_ _1141_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2696_ clknet_2_1__leaf_clk _0172_ net62 VGND VGND VPWR VPWR PC.i_mem_addr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1716_ _0675_ _0867_ _0869_ _0880_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1647_ _0984_ _0985_ _0988_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__a21bo_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1578_ RegFile.L\[4\] _0680_ _0685_ RegFile.C\[4\] VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__a22o_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2550_ net46 _0583_ _0584_ _0585_ ALU.immediate\[8\] VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2481_ _0678_ _0524_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__nor2_1
X_1501_ _0655_ _0838_ _0839_ _0842_ _0828_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__a311o_1
X_1432_ _0760_ _0652_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__or2_2
X_1363_ _0699_ _0703_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__nor2_8
XFILLER_0_37_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1294_ _0624_ _0622_ ByteBuffer.instr\[21\] VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2679_ net69 _0155_ net59 VGND VGND VPWR VPWR RegFile.A\[5\] sky130_fd_sc_hd__dfrtp_4
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1981_ _0883_ _1172_ _1168_ _1058_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2533_ _0571_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__clkbuf_1
X_2602_ clknet_2_0__leaf_clk _0078_ net59 VGND VGND VPWR VPWR ByteBuffer.instr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2395_ _0508_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
X_1415_ ByteBuffer.instr\[22\] _0642_ _0635_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__or3_2
X_1346_ RegFile.D\[6\] _0683_ net52 RegFile.B\[6\] _0687_ VGND VGND VPWR VPWR _0688_
+ sky130_fd_sc_hd__a221o_1
X_1277_ ByteBuffer.instr\[16\] VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2180_ _0354_ _0358_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1895_ _1151_ _1134_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1964_ _1256_ _1175_ _0816_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2516_ PC.i_mem_addr\[3\] _0551_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2447_ clknet_1_0__leaf__0514_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__buf_1
XFILLER_0_11_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1329_ _0670_ _0661_ _0639_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__or3_1
X_2378_ _0434_ _0624_ _0497_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__mux2_1
X_2458__56 clknet_1_1__leaf__0517_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__inv_2
XFILLER_0_34_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold9 ALU.flags_to_alu\[1\] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1680_ _1020_ _1021_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__nand2_2
X_2301_ _0203_ _0454_ _0458_ _0441_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__o211a_1
XFILLER_0_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2232_ ByteBuffer.counter\[1\] _0659_ ByteBuffer.counter\[0\] VGND VGND VPWR VPWR
+ _0407_ sky130_fd_sc_hd__or3b_1
XFILLER_0_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2163_ _0273_ net47 _0336_ net139 VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2094_ RegFile.E\[5\] _0273_ _0297_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__mux2_1
X_1947_ _0736_ _1082_ _0734_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__a21boi_1
X_1878_ _1100_ _1210_ _1212_ _1213_ _1218_ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__o221a_1
XFILLER_0_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1732_ _1071_ _1072_ _1073_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__a21o_1
X_1801_ _1137_ _1142_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1663_ RegFile.B\[5\] _0705_ _1004_ _0711_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__a211o_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ _0922_ _0934_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2215_ _1124_ _0391_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2146_ _0329_ _0696_ _0618_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__a21o_1
X_2077_ RegFile.D\[5\] _1247_ _0288_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2000_ _1109_ _1123_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2695_ clknet_2_2__leaf_clk _0171_ net63 VGND VGND VPWR VPWR PC.i_mem_addr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1646_ _0986_ _0970_ _0982_ _0987_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__o31a_1
X_1715_ _0816_ _0831_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__xor2_4
XFILLER_0_5_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1577_ ALU.flags_to_alu\[4\] _0687_ _0683_ RegFile.E\[4\] _0654_ VGND VGND VPWR VPWR
+ _0919_ sky130_fd_sc_hd__a221o_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2129_ _0273_ RegFile.L\[5\] _0316_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2480_ ByteBuffer.instr\[19\] _0639_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__nand2_1
X_1500_ ALU.flags_to_alu\[3\] _0704_ _0841_ _0629_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__o211a_1
X_1293_ ByteBuffer.instr\[17\] _0624_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__xor2_4
XFILLER_0_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1362_ _0699_ _0703_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__nand2_8
X_1431_ RegFile.L\[5\] _0770_ _0771_ RegFile.B\[5\] net51 VGND VGND VPWR VPWR _0773_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2421__21 clknet_1_1__leaf__0515_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__inv_2
X_1629_ RegFile.A\[6\] _0792_ _0704_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__or3_1
X_2678_ net68 _0154_ net58 VGND VGND VPWR VPWR RegFile.A\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1980_ _1139_ _0213_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2532_ PC.i_mem_addr\[5\] _0570_ _0542_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__mux2_1
X_2601_ clknet_2_1__leaf_clk _0077_ net62 VGND VGND VPWR VPWR ALU.immediate\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1414_ _0754_ _0755_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__nand2_2
XFILLER_0_48_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1276_ ByteBuffer.instr\[19\] VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__inv_2
X_2394_ _0434_ ALU.immediate\[2\] _0408_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__mux2_1
X_1345_ _0686_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire56 _0706_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1894_ _0806_ _1210_ _1229_ _1213_ _1233_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__o221a_1
X_1963_ _1210_ _1168_ _1057_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2515_ PC.i_mem_addr\[3\] _0551_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1328_ _0645_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__clkinv_4
X_2377_ _0499_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2300_ PC.i_mem_addr\[2\] _0451_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__or2_1
X_2231_ ByteBuffer.counter\[1\] ByteBuffer.next_counter\[0\] VGND VGND VPWR VPWR _0406_
+ sky130_fd_sc_hd__nand2_4
X_2162_ net142 _0336_ _0343_ _0344_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2093_ _0299_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1946_ _1273_ _0179_ _0181_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__o21a_2
X_1877_ _1070_ _1172_ _1216_ _1217_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1800_ _1139_ _1141_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1731_ _0781_ _0782_ _0802_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1662_ RegFile.H\[5\] _0707_ _0709_ RegFile.D\[5\] VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__a22o_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _1096_ _1125_ _0986_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__a21o_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1593_ _0922_ _0934_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2145_ _0619_ _0620_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__nand2_1
X_2428__27 clknet_1_0__leaf__0516_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__inv_2
X_2076_ _0290_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1929_ _1022_ _1266_ _1267_ _1092_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2442__41 clknet_1_1__leaf__0516_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__inv_2
XFILLER_0_22_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2694_ clknet_2_2__leaf_clk _0170_ net63 VGND VGND VPWR VPWR PC.i_mem_addr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1714_ _0855_ _0844_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__nor2_1
X_1645_ _0947_ _0959_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1576_ _0914_ _0916_ _0917_ _0774_ RegFile.A\[4\] VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__o32a_1
XFILLER_0_67_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2059_ _0278_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__clkbuf_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2128_ _0318_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1430_ _0638_ net57 _0650_ _0760_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__nor4_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1292_ ByteBuffer.instr\[20\] _0633_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__nand2_1
X_1361_ _0622_ _0701_ _0702_ _0626_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__o22a_4
XFILLER_0_26_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1628_ _0780_ _0969_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__nand2_4
X_1559_ net57 _0650_ _0762_ _0684_ ALU.flags_to_alu\[0\] VGND VGND VPWR VPWR _0901_
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_1_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2677_ net67 _0153_ net58 VGND VGND VPWR VPWR RegFile.A\[3\] sky130_fd_sc_hd__dfrtp_4
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2600_ clknet_2_1__leaf_clk _0076_ net62 VGND VGND VPWR VPWR ALU.immediate\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2531_ _0566_ _0569_ net46 VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__mux2_1
X_1413_ _0749_ _0753_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2393_ _0507_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1344_ _0684_ _0677_ _0679_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__and3_1
Xwire46 _0540_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_4
XFILLER_0_58_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1962_ _0855_ _1165_ _1164_ _0196_ _1166_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1893_ _1073_ _1168_ _1231_ _1232_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2514_ ALU.immediate\[3\] _0853_ _0519_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__mux2_1
X_2376_ _0435_ _0622_ _0497_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__mux2_1
X_1327_ _0667_ _0668_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2449__47 clknet_1_0__leaf__0517_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__inv_2
XFILLER_0_52_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2230_ net132 _0659_ VGND VGND VPWR VPWR ByteBuffer.next_counter\[0\] sky130_fd_sc_hd__nor2_1
X_2161_ _1201_ _0271_ _0334_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__o21a_1
X_2092_ RegFile.E\[6\] _0271_ _0297_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__mux2_1
X_1945_ _0180_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2463__61 clknet_1_0__leaf__0517_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__inv_2
X_1876_ _1175_ _1174_ _1069_ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2359_ _0434_ ALU.immediate\[10\] _0406_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1730_ _0780_ _0921_ _0929_ _0933_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__nand4_2
X_1592_ ALU.immediate\[4\] _0675_ _0929_ _0933_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1661_ RegFile.A\[5\] _0652_ _0676_ _1002_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__o211a_2
XFILLER_0_21_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ _0619_ _0668_ _0620_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__a21oi_1
X_2213_ _0281_ _0390_ _0334_ net137 VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2075_ RegFile.D\[6\] _1225_ _0288_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__mux2_1
X_1928_ _1022_ _1266_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__nand2_1
X_1859_ _1200_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1713_ _0756_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2693_ clknet_2_2__leaf_clk _0169_ net63 VGND VGND VPWR VPWR PC.i_mem_addr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1644_ _0947_ _0959_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__and2_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1575_ RegFile.L\[4\] _0770_ _0771_ RegFile.B\[4\] net51 VGND VGND VPWR VPWR _0917_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2127_ _0271_ RegFile.L\[6\] _0316_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2058_ RegFile.C\[3\] _0277_ _0269_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__mux2_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1360_ ByteBuffer.instr\[21\] _0667_ _0668_ _0696_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1291_ _0619_ _0622_ _0624_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_58_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2676_ net66 _0152_ net58 VGND VGND VPWR VPWR RegFile.A\[2\] sky130_fd_sc_hd__dfrtp_4
X_1489_ ALU.immediate\[2\] _0674_ _0829_ _0830_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__o211a_4
X_1558_ net57 _0650_ _0766_ _0684_ RegFile.D\[0\] VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__o2111a_1
X_1627_ _0654_ _0966_ _0967_ _0968_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__o2bb2a_2
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2412__12 clknet_1_1__leaf__0515_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__inv_2
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2530_ _0567_ _0568_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1412_ _0749_ _0753_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__nand2_1
X_2392_ _0435_ ALU.immediate\[1\] _0408_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__mux2_1
X_1343_ _0677_ _0679_ _0684_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_64_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2659_ net113 _0135_ net60 VGND VGND VPWR VPWR RegFile.C\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1892_ _1174_ _1175_ _0781_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1961_ _0675_ _0867_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__nor2_1
X_2513_ _0554_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1326_ ByteBuffer.instr\[20\] ByteBuffer.instr\[21\] VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__nand2b_1
X_2375_ _0498_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2160_ _1201_ _0342_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap1 _0772_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__buf_1
X_2091_ _0298_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1944_ _1093_ _1145_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__nor2_1
X_1875_ _0781_ _1214_ _1076_ _1168_ _1215_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__o221a_1
XFILLER_0_43_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2427_ clknet_1_0__leaf__0514_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__buf_1
X_2358_ _0488_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
X_2289_ ByteBuffer.instr\[19\] _0621_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__or2_2
X_1309_ _0638_ _0646_ _0650_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1591_ _0930_ _0931_ _0932_ _0693_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__o31a_1
X_1660_ RegFile.H\[5\] net53 _1001_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2143_ _0263_ _0326_ _1201_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__mux2_1
X_2212_ net47 VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2074_ _0289_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1927_ _1000_ _1085_ _1043_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1858_ _1196_ _0627_ _1199_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__or3b_1
XFILLER_0_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1789_ _0983_ _1128_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2692_ clknet_2_3__leaf_clk _0168_ net63 VGND VGND VPWR VPWR PC.i_mem_addr\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_1712_ _0746_ _1053_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__nand2_1
X_1643_ _0804_ _0935_ _0805_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_5_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2433__32 clknet_1_1__leaf__0516_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__inv_2
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1574_ ALU.flags_to_alu\[4\] _0765_ _0767_ RegFile.D\[4\] _0915_ VGND VGND VPWR VPWR
+ _0916_ sky130_fd_sc_hd__a221o_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2057_ _0182_ _0261_ _0262_ net6 VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__a22o_2
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2126_ _0317_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1290_ ByteBuffer.instr\[23\] ByteBuffer.instr\[22\] VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_37_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1626_ RegFile.L\[6\] _0680_ _0685_ RegFile.C\[6\] VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__a22o_1
X_2675_ net65 _0151_ net60 VGND VGND VPWR VPWR RegFile.A\[1\] sky130_fd_sc_hd__dfrtp_4
X_1488_ _0664_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__inv_2
X_1557_ net57 _0650_ _0762_ _0638_ RegFile.H\[0\] VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__o2111a_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2109_ _0308_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1411_ ALU.immediate\[8\] _0675_ _0693_ _0752_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__a22o_1
X_2391_ _0506_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
X_1342_ _0637_ _0634_ _0632_ _0622_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2589_ _0617_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__clkbuf_1
X_2658_ net112 _0134_ net61 VGND VGND VPWR VPWR RegFile.C\[0\] sky130_fd_sc_hd__dfrtp_1
X_1609_ RegFile.E\[7\] _0789_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1891_ _1071_ _1172_ _1214_ _0922_ _1230_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__o221a_1
X_1960_ _1062_ _1172_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2512_ PC.i_mem_addr\[2\] _0553_ _0542_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1325_ _0622_ _0624_ ByteBuffer.instr\[19\] _0619_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__or4bb_1
X_2374_ _0425_ _0619_ _0497_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2090_ RegFile.E\[7\] _0263_ _0297_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1943_ _1146_ _1274_ _0174_ _1161_ _0178_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__a221o_1
X_1874_ _1066_ _1165_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2357_ _0435_ ALU.immediate\[9\] _0406_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__mux2_1
X_2288_ _0261_ _0412_ _0441_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__a21boi_2
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1308_ _0649_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__clkbuf_4
X_2454__52 clknet_1_1__leaf__0517_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__inv_2
XFILLER_0_15_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1590_ RegFile.E\[4\] _0699_ net55 _0654_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__a31o_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2142_ _1183_ _0325_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__nand2_1
X_2211_ _0389_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
X_2073_ RegFile.D\[7\] _1184_ _0288_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1788_ _0960_ _1129_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1926_ _1227_ _1249_ _1263_ _1264_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__a211o_2
X_1857_ _0632_ _1197_ _1198_ _0663_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2419__19 clknet_1_0__leaf__0515_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__inv_2
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2691_ clknet_2_2__leaf_clk _0167_ net63 VGND VGND VPWR VPWR PC.i_mem_addr\[9\] sky130_fd_sc_hd__dfrtp_1
X_1711_ _0991_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1642_ _0960_ _0983_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ RegFile.C\[4\] _0638_ _0681_ _0760_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__and4_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2125_ _0263_ RegFile.L\[7\] _0316_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__mux2_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2056_ _0276_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__clkbuf_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1909_ _1248_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2674_ net128 _0150_ net61 VGND VGND VPWR VPWR RegFile.A\[0\] sky130_fd_sc_hd__dfrtp_2
X_1625_ ALU.flags_to_alu\[6\] _0687_ _0683_ RegFile.E\[6\] _0654_ VGND VGND VPWR VPWR
+ _0967_ sky130_fd_sc_hd__a221o_1
X_1556_ RegFile.L\[0\] _0770_ _0771_ RegFile.B\[0\] _0897_ VGND VGND VPWR VPWR _0898_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ _0654_ _0823_ _0824_ _0827_ _0828_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__a311o_1
XFILLER_0_49_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2039_ _1182_ _0261_ _0262_ net10 VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__a22o_1
X_2108_ _1184_ RegFile.H\[7\] net48 VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1410_ RegFile.A\[0\] _0704_ _0751_ _0630_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__o211a_1
X_2390_ _0425_ ALU.immediate\[0\] _0408_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1341_ _0682_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__buf_4
XFILLER_0_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2588_ PC.i_mem_addr\[15\] _0616_ _0542_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__mux2_1
X_1539_ _0869_ _0880_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__nand2_1
X_2657_ net111 _0133_ net58 VGND VGND VPWR VPWR RegFile.D\[7\] sky130_fd_sc_hd__dfrtp_2
X_1608_ RegFile.C\[7\] _0793_ _0786_ RegFile.D\[7\] VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1890_ _1069_ _1165_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2511_ _0549_ _0552_ net46 VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__mux2_1
X_2373_ _0496_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1324_ _0633_ _0665_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__or2_2
XFILLER_0_24_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1942_ _1113_ _1210_ _0177_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1873_ _1122_ _1163_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__or2_2
XFILLER_0_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2356_ _0487_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1307_ _0620_ _0647_ _0648_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2287_ _0449_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2210_ ALU.flags_to_alu\[2\] _0388_ _0334_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2141_ _0630_ _1094_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__nand2_1
X_2072_ _0286_ _0287_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__nor2_4
X_1925_ _0937_ _1114_ _1116_ _1124_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1787_ _1100_ _1128_ _1070_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__o21ai_1
X_1856_ ByteBuffer.instr\[19\] _0660_ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2339_ _0724_ _0476_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2690_ clknet_2_3__leaf_clk _0166_ net63 VGND VGND VPWR VPWR PC.i_mem_addr\[8\] sky130_fd_sc_hd__dfrtp_1
X_1710_ _0726_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__inv_2
X_1641_ _0970_ _0982_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1572_ RegFile.E\[4\] _0761_ _0763_ RegFile.H\[4\] VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__a22o_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2124_ _0267_ _0306_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__nand2_4
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2055_ RegFile.C\[4\] _0275_ _0269_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1839_ _1130_ _1166_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1908_ RegFile.A\[5\] _1247_ _1203_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput40 net40 VGND VGND VPWR VPWR gpo[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1555_ RegFile.C\[0\] _0638_ _0681_ _0760_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__and4_1
X_2673_ net127 _0149_ net60 VGND VGND VPWR VPWR RegFile.B\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1624_ _0961_ _0963_ _0964_ net50 _0965_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__a32o_1
X_1486_ _0664_ _0692_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__or2_2
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2107_ _0630_ _0264_ _0306_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2038_ ByteBuffer.instr\[19\] net1 net4 _0260_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__and4_2
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1340_ _0638_ _0681_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2656_ net110 _0132_ net59 VGND VGND VPWR VPWR RegFile.D\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2587_ ALU.immediate\[15\] _0585_ _0615_ _0540_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__a22o_1
X_1538_ _0654_ _0876_ _0879_ _0828_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__a211o_1
X_1607_ ALU.flags_to_alu\[7\] _0788_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__and2_1
X_1469_ RegFile.E\[2\] _0761_ _0771_ RegFile.B\[2\] VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2510_ _0550_ _0551_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2372_ ByteBuffer.counter\[0\] ByteBuffer.counter\[1\] _0659_ VGND VGND VPWR VPWR
+ _0496_ sky130_fd_sc_hd__or3_1
X_1323_ _0622_ _0618_ _0647_ _0619_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2639_ net93 _0115_ net58 VGND VGND VPWR VPWR RegFile.H\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1941_ _1061_ _1172_ _1256_ _1056_ _0176_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__o221a_1
X_1872_ _1092_ _1160_ _1151_ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2355_ _0425_ ALU.immediate\[8\] _0406_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__mux2_1
X_1306_ ByteBuffer.instr\[23\] ByteBuffer.instr\[22\] VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__and2_2
X_2286_ RegFile.A\[7\] net1 VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ _0324_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2071_ _0655_ _0266_ _0268_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__o21ai_4
X_1924_ _1093_ _1136_ _1213_ _1252_ _1262_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__o221ai_1
X_1855_ _0645_ _0700_ _0661_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__a21o_1
X_1786_ _0806_ _1127_ _1074_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2269_ _0410_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__inv_2
X_2407_ clknet_1_1__leaf__0514_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__buf_1
X_2338_ _0479_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2469__3 clknet_1_0__leaf__0514_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__inv_2
XFILLER_0_53_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1571_ _0855_ _0844_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__or2b_1
X_1640_ _0693_ _0978_ _0981_ _0675_ ALU.immediate\[6\] VGND VGND VPWR VPWR _0982_
+ sky130_fd_sc_hd__a32o_4
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ _0315_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2054_ _1265_ _0261_ _0262_ net7 VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__a22o_2
XFILLER_0_29_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2424__24 clknet_1_1__leaf__0515_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__inv_2
X_1838_ _1158_ _1161_ _1179_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__a21o_1
X_1907_ _0655_ _1239_ _1246_ _0631_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__a22o_2
XFILLER_0_29_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1769_ _0868_ _0881_ _1108_ _1110_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput41 net41 VGND VGND VPWR VPWR gpo[5] sky130_fd_sc_hd__clkbuf_4
Xoutput30 net30 VGND VGND VPWR VPWR gpo[26] sky130_fd_sc_hd__buf_2
XFILLER_0_50_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2672_ net126 _0148_ net59 VGND VGND VPWR VPWR RegFile.B\[6\] sky130_fd_sc_hd__dfrtp_2
X_1554_ _0629_ _0892_ _0895_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__o21ai_4
X_1623_ RegFile.A\[6\] VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__inv_2
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1485_ ALU.flags_to_alu\[2\] _0704_ _0826_ _0629_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__o211a_1
.ends

