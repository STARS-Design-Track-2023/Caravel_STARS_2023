VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO silly_synthesizer
  CLASS BLOCK ;
  FOREIGN silly_synthesizer ;
  ORIGIN 0.000 0.000 ;
  SIZE 231.685 BY 242.405 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 231.440 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 231.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 231.440 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END clk
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 227.685 221.040 231.685 221.640 ;
    END
  END cs
  PIN gpio[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 209.390 238.405 209.670 242.405 ;
    END
  END gpio[0]
  PIN gpio[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 238.405 119.510 242.405 ;
    END
  END gpio[10]
  PIN gpio[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END gpio[11]
  PIN gpio[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END gpio[12]
  PIN gpio[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 227.685 34.040 231.685 34.640 ;
    END
  END gpio[13]
  PIN gpio[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END gpio[14]
  PIN gpio[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 227.685 173.440 231.685 174.040 ;
    END
  END gpio[15]
  PIN gpio[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END gpio[16]
  PIN gpio[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END gpio[1]
  PIN gpio[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END gpio[2]
  PIN gpio[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END gpio[3]
  PIN gpio[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 238.405 74.430 242.405 ;
    END
  END gpio[4]
  PIN gpio[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 227.685 125.840 231.685 126.440 ;
    END
  END gpio[5]
  PIN gpio[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END gpio[6]
  PIN gpio[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 164.310 238.405 164.590 242.405 ;
    END
  END gpio[7]
  PIN gpio[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END gpio[8]
  PIN gpio[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END gpio[9]
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 238.405 32.570 242.405 ;
    END
  END nrst
  PIN pwm
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 227.685 81.640 231.685 82.240 ;
    END
  END pwm
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 225.860 231.285 ;
      LAYER met1 ;
        RECT 0.070 10.640 226.710 231.440 ;
      LAYER met2 ;
        RECT 0.100 238.125 32.010 239.090 ;
        RECT 32.850 238.125 73.870 239.090 ;
        RECT 74.710 238.125 118.950 239.090 ;
        RECT 119.790 238.125 164.030 239.090 ;
        RECT 164.870 238.125 209.110 239.090 ;
        RECT 209.950 238.125 226.690 239.090 ;
        RECT 0.100 4.280 226.690 238.125 ;
        RECT 0.650 4.000 41.670 4.280 ;
        RECT 42.510 4.000 86.750 4.280 ;
        RECT 87.590 4.000 131.830 4.280 ;
        RECT 132.670 4.000 173.690 4.280 ;
        RECT 174.530 4.000 218.770 4.280 ;
        RECT 219.610 4.000 226.690 4.280 ;
      LAYER met3 ;
        RECT 4.400 230.840 227.685 231.705 ;
        RECT 4.000 222.040 227.685 230.840 ;
        RECT 4.000 220.640 227.285 222.040 ;
        RECT 4.000 184.640 227.685 220.640 ;
        RECT 4.400 183.240 227.685 184.640 ;
        RECT 4.000 174.440 227.685 183.240 ;
        RECT 4.000 173.040 227.285 174.440 ;
        RECT 4.000 140.440 227.685 173.040 ;
        RECT 4.400 139.040 227.685 140.440 ;
        RECT 4.000 126.840 227.685 139.040 ;
        RECT 4.000 125.440 227.285 126.840 ;
        RECT 4.000 92.840 227.685 125.440 ;
        RECT 4.400 91.440 227.685 92.840 ;
        RECT 4.000 82.640 227.685 91.440 ;
        RECT 4.000 81.240 227.285 82.640 ;
        RECT 4.000 45.240 227.685 81.240 ;
        RECT 4.400 43.840 227.685 45.240 ;
        RECT 4.000 35.040 227.685 43.840 ;
        RECT 4.000 33.640 227.285 35.040 ;
        RECT 4.000 10.715 227.685 33.640 ;
      LAYER met4 ;
        RECT 61.935 34.175 97.440 173.225 ;
        RECT 99.840 34.175 166.225 173.225 ;
  END
END silly_synthesizer
END LIBRARY

