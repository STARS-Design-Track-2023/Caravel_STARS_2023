magic
tech sky130A
magscale 1 2
timestamp 1693969699
<< viali >>
rect 1685 27081 1719 27115
rect 3893 27081 3927 27115
rect 15761 27081 15795 27115
rect 11069 27013 11103 27047
rect 13185 27013 13219 27047
rect 1777 26945 1811 26979
rect 4169 26945 4203 26979
rect 7389 26945 7423 26979
rect 10793 26945 10827 26979
rect 10977 26945 11011 26979
rect 11161 26945 11195 26979
rect 11713 26945 11747 26979
rect 13093 26945 13127 26979
rect 15669 26945 15703 26979
rect 16773 26945 16807 26979
rect 19441 26945 19475 26979
rect 21005 26945 21039 26979
rect 23489 26945 23523 26979
rect 10609 26877 10643 26911
rect 13369 26877 13403 26911
rect 20729 26877 20763 26911
rect 7205 26741 7239 26775
rect 9965 26741 9999 26775
rect 11345 26741 11379 26775
rect 11897 26741 11931 26775
rect 12725 26741 12759 26775
rect 16957 26741 16991 26775
rect 19625 26741 19659 26775
rect 23305 26741 23339 26775
rect 10701 26537 10735 26571
rect 20808 26537 20842 26571
rect 12909 26469 12943 26503
rect 15393 26469 15427 26503
rect 15945 26469 15979 26503
rect 5917 26401 5951 26435
rect 7389 26401 7423 26435
rect 7481 26401 7515 26435
rect 13553 26401 13587 26435
rect 16497 26401 16531 26435
rect 17417 26401 17451 26435
rect 20545 26401 20579 26435
rect 22293 26401 22327 26435
rect 5641 26333 5675 26367
rect 8953 26333 8987 26367
rect 11345 26333 11379 26367
rect 12449 26333 12483 26367
rect 12817 26333 12851 26367
rect 14657 26333 14691 26367
rect 14841 26333 14875 26367
rect 15117 26333 15151 26367
rect 15209 26333 15243 26367
rect 15761 26333 15795 26367
rect 16405 26333 16439 26367
rect 17509 26333 17543 26367
rect 18797 26333 18831 26367
rect 22477 26333 22511 26367
rect 23029 26333 23063 26367
rect 9229 26265 9263 26299
rect 13369 26265 13403 26299
rect 14105 26265 14139 26299
rect 15025 26265 15059 26299
rect 16313 26265 16347 26299
rect 16773 26265 16807 26299
rect 18153 26265 18187 26299
rect 8125 26197 8159 26231
rect 10793 26197 10827 26231
rect 11897 26197 11931 26231
rect 12633 26197 12667 26231
rect 13277 26197 13311 26231
rect 15577 26197 15611 26231
rect 18245 26197 18279 26231
rect 10241 25993 10275 26027
rect 13921 25993 13955 26027
rect 14013 25993 14047 26027
rect 7941 25925 7975 25959
rect 12449 25925 12483 25959
rect 16957 25925 16991 25959
rect 18797 25925 18831 25959
rect 22201 25925 22235 25959
rect 10425 25857 10459 25891
rect 11345 25857 11379 25891
rect 11897 25857 11931 25891
rect 14749 25857 14783 25891
rect 21281 25857 21315 25891
rect 6101 25789 6135 25823
rect 6469 25789 6503 25823
rect 8217 25789 8251 25823
rect 8493 25789 8527 25823
rect 8769 25789 8803 25823
rect 10885 25789 10919 25823
rect 12173 25789 12207 25823
rect 14565 25789 14599 25823
rect 15025 25789 15059 25823
rect 16681 25789 16715 25823
rect 18429 25789 18463 25823
rect 18521 25789 18555 25823
rect 20637 25789 20671 25823
rect 21925 25789 21959 25823
rect 5549 25653 5583 25687
rect 11161 25653 11195 25687
rect 12081 25653 12115 25687
rect 16497 25653 16531 25687
rect 20269 25653 20303 25687
rect 21189 25653 21223 25687
rect 21465 25653 21499 25687
rect 23673 25653 23707 25687
rect 8953 25449 8987 25483
rect 10320 25449 10354 25483
rect 11805 25449 11839 25483
rect 12160 25449 12194 25483
rect 13645 25449 13679 25483
rect 16957 25449 16991 25483
rect 21005 25449 21039 25483
rect 25881 25449 25915 25483
rect 9229 25381 9263 25415
rect 16221 25381 16255 25415
rect 5273 25313 5307 25347
rect 7205 25313 7239 25347
rect 9781 25313 9815 25347
rect 10057 25313 10091 25347
rect 11897 25313 11931 25347
rect 14473 25313 14507 25347
rect 14749 25313 14783 25347
rect 17509 25313 17543 25347
rect 17785 25313 17819 25347
rect 19533 25313 19567 25347
rect 21097 25313 21131 25347
rect 21373 25313 21407 25347
rect 22845 25313 22879 25347
rect 23489 25313 23523 25347
rect 24961 25313 24995 25347
rect 1409 25245 1443 25279
rect 4997 25245 5031 25279
rect 6837 25245 6871 25279
rect 8585 25245 8619 25279
rect 9137 25245 9171 25279
rect 9689 25245 9723 25279
rect 17325 25245 17359 25279
rect 17417 25245 17451 25279
rect 18337 25245 18371 25279
rect 18521 25245 18555 25279
rect 18797 25245 18831 25279
rect 18889 25245 18923 25279
rect 19257 25245 19291 25279
rect 25697 25245 25731 25279
rect 18705 25177 18739 25211
rect 22937 25177 22971 25211
rect 1593 25109 1627 25143
rect 6745 25109 6779 25143
rect 8769 25109 8803 25143
rect 9597 25109 9631 25143
rect 19073 25109 19107 25143
rect 24409 25109 24443 25143
rect 8769 24905 8803 24939
rect 9137 24905 9171 24939
rect 11529 24905 11563 24939
rect 11897 24905 11931 24939
rect 7021 24837 7055 24871
rect 15945 24837 15979 24871
rect 23857 24837 23891 24871
rect 6469 24769 6503 24803
rect 7205 24769 7239 24803
rect 9229 24769 9263 24803
rect 9597 24769 9631 24803
rect 13001 24769 13035 24803
rect 15577 24769 15611 24803
rect 15670 24769 15704 24803
rect 15853 24769 15887 24803
rect 16083 24769 16117 24803
rect 16865 24769 16899 24803
rect 21557 24769 21591 24803
rect 21925 24769 21959 24803
rect 4445 24701 4479 24735
rect 4721 24701 4755 24735
rect 7297 24701 7331 24735
rect 9413 24701 9447 24735
rect 9873 24701 9907 24735
rect 11989 24701 12023 24735
rect 12173 24701 12207 24735
rect 13277 24701 13311 24735
rect 14841 24701 14875 24735
rect 15393 24701 15427 24735
rect 16957 24701 16991 24735
rect 17233 24701 17267 24735
rect 19717 24701 19751 24735
rect 21281 24701 21315 24735
rect 24133 24701 24167 24735
rect 7573 24633 7607 24667
rect 14749 24633 14783 24667
rect 18705 24633 18739 24667
rect 6193 24565 6227 24599
rect 7205 24565 7239 24599
rect 11345 24565 11379 24599
rect 16221 24565 16255 24599
rect 16681 24565 16715 24599
rect 19073 24565 19107 24599
rect 19809 24565 19843 24599
rect 22017 24565 22051 24599
rect 22385 24565 22419 24599
rect 5825 24361 5859 24395
rect 10149 24361 10183 24395
rect 12081 24361 12115 24395
rect 13093 24361 13127 24395
rect 16392 24361 16426 24395
rect 17969 24361 18003 24395
rect 20821 24361 20855 24395
rect 23489 24361 23523 24395
rect 15209 24293 15243 24327
rect 18797 24293 18831 24327
rect 21649 24293 21683 24327
rect 8217 24225 8251 24259
rect 11069 24225 11103 24259
rect 11253 24225 11287 24259
rect 12173 24225 12207 24259
rect 12725 24225 12759 24259
rect 13277 24225 13311 24259
rect 15025 24225 15059 24259
rect 15853 24225 15887 24259
rect 16129 24225 16163 24259
rect 18429 24225 18463 24259
rect 18613 24225 18647 24259
rect 20269 24225 20303 24259
rect 21097 24225 21131 24259
rect 21189 24225 21223 24259
rect 22477 24225 22511 24259
rect 23121 24225 23155 24259
rect 5641 24157 5675 24191
rect 5825 24157 5859 24191
rect 10333 24157 10367 24191
rect 10977 24157 11011 24191
rect 11437 24157 11471 24191
rect 11530 24157 11564 24191
rect 11805 24157 11839 24191
rect 11943 24157 11977 24191
rect 12909 24157 12943 24191
rect 13553 24157 13587 24191
rect 14289 24157 14323 24191
rect 14473 24157 14507 24191
rect 15669 24157 15703 24191
rect 18981 24157 19015 24191
rect 19809 24157 19843 24191
rect 22293 24157 22327 24191
rect 23213 24157 23247 24191
rect 23673 24157 23707 24191
rect 11713 24089 11747 24123
rect 18337 24089 18371 24123
rect 19257 24089 19291 24123
rect 21281 24089 21315 24123
rect 7573 24021 7607 24055
rect 10609 24021 10643 24055
rect 13461 24021 13495 24055
rect 13921 24021 13955 24055
rect 14105 24021 14139 24055
rect 15577 24021 15611 24055
rect 17877 24021 17911 24055
rect 20361 24021 20395 24055
rect 20453 24021 20487 24055
rect 21741 24021 21775 24055
rect 23397 24021 23431 24055
rect 5273 23817 5307 23851
rect 8309 23817 8343 23851
rect 14933 23817 14967 23851
rect 15853 23817 15887 23851
rect 19993 23817 20027 23851
rect 20361 23817 20395 23851
rect 21281 23817 21315 23851
rect 5181 23749 5215 23783
rect 6101 23749 6135 23783
rect 13461 23749 13495 23783
rect 19625 23749 19659 23783
rect 21189 23749 21223 23783
rect 23949 23749 23983 23783
rect 4813 23681 4847 23715
rect 6009 23681 6043 23715
rect 9045 23681 9079 23715
rect 9321 23681 9355 23715
rect 10793 23681 10827 23715
rect 12909 23681 12943 23715
rect 13185 23681 13219 23715
rect 15209 23681 15243 23715
rect 16681 23681 16715 23715
rect 19073 23681 19107 23715
rect 19257 23681 19291 23715
rect 19350 23681 19384 23715
rect 19533 23681 19567 23715
rect 19722 23681 19756 23715
rect 20453 23681 20487 23715
rect 22109 23681 22143 23715
rect 22385 23681 22419 23715
rect 4721 23613 4755 23647
rect 5089 23613 5123 23647
rect 5825 23613 5859 23647
rect 6561 23613 6595 23647
rect 6837 23613 6871 23647
rect 12633 23613 12667 23647
rect 16957 23613 16991 23647
rect 18429 23613 18463 23647
rect 20637 23613 20671 23647
rect 21465 23613 21499 23647
rect 22201 23613 22235 23647
rect 22477 23613 22511 23647
rect 24225 23613 24259 23647
rect 4537 23477 4571 23511
rect 8401 23477 8435 23511
rect 9137 23477 9171 23511
rect 10609 23477 10643 23511
rect 11989 23477 12023 23511
rect 13001 23477 13035 23511
rect 18521 23477 18555 23511
rect 19901 23477 19935 23511
rect 20821 23477 20855 23511
rect 21925 23477 21959 23511
rect 22109 23477 22143 23511
rect 8769 23273 8803 23307
rect 16589 23273 16623 23307
rect 18061 23273 18095 23307
rect 22109 23273 22143 23307
rect 22293 23273 22327 23307
rect 23305 23273 23339 23307
rect 6929 23205 6963 23239
rect 4077 23137 4111 23171
rect 7021 23137 7055 23171
rect 9045 23137 9079 23171
rect 10517 23137 10551 23171
rect 11989 23137 12023 23171
rect 17417 23137 17451 23171
rect 21005 23137 21039 23171
rect 21925 23137 21959 23171
rect 22661 23137 22695 23171
rect 22845 23137 22879 23171
rect 24133 23137 24167 23171
rect 6377 23069 6411 23103
rect 6745 23069 6779 23103
rect 10241 23069 10275 23103
rect 12541 23069 12575 23103
rect 12817 23069 12851 23103
rect 12909 23069 12943 23103
rect 13093 23069 13127 23103
rect 16037 23069 16071 23103
rect 16405 23069 16439 23103
rect 17601 23069 17635 23103
rect 17693 23069 17727 23103
rect 18613 23069 18647 23103
rect 18889 23069 18923 23103
rect 19257 23069 19291 23103
rect 21649 23069 21683 23103
rect 22109 23069 22143 23103
rect 4353 23001 4387 23035
rect 6101 23001 6135 23035
rect 6561 23001 6595 23035
rect 6653 23001 6687 23035
rect 7297 23001 7331 23035
rect 9873 23001 9907 23035
rect 16221 23001 16255 23035
rect 16313 23001 16347 23035
rect 19533 23001 19567 23035
rect 21833 23001 21867 23035
rect 18797 22933 18831 22967
rect 19073 22933 19107 22967
rect 21097 22933 21131 22967
rect 22937 22933 22971 22967
rect 23581 22933 23615 22967
rect 4905 22729 4939 22763
rect 7297 22729 7331 22763
rect 11529 22729 11563 22763
rect 11897 22729 11931 22763
rect 20821 22729 20855 22763
rect 6929 22661 6963 22695
rect 8493 22661 8527 22695
rect 19349 22661 19383 22695
rect 4997 22593 5031 22627
rect 5365 22593 5399 22627
rect 5825 22593 5859 22627
rect 6745 22593 6779 22627
rect 7021 22593 7055 22627
rect 7113 22593 7147 22627
rect 8217 22593 8251 22627
rect 11161 22593 11195 22627
rect 14657 22593 14691 22627
rect 19073 22593 19107 22627
rect 21465 22593 21499 22627
rect 22017 22593 22051 22627
rect 22293 22593 22327 22627
rect 2697 22525 2731 22559
rect 2973 22525 3007 22559
rect 4445 22525 4479 22559
rect 10057 22525 10091 22559
rect 10609 22525 10643 22559
rect 11989 22525 12023 22559
rect 12173 22525 12207 22559
rect 12909 22525 12943 22559
rect 14749 22525 14783 22559
rect 14933 22525 14967 22559
rect 16037 22525 16071 22559
rect 22569 22525 22603 22559
rect 22201 22457 22235 22491
rect 9965 22389 9999 22423
rect 10977 22389 11011 22423
rect 12357 22389 12391 22423
rect 14289 22389 14323 22423
rect 15485 22389 15519 22423
rect 20913 22389 20947 22423
rect 24041 22389 24075 22423
rect 22477 22185 22511 22219
rect 14749 22117 14783 22151
rect 22385 22117 22419 22151
rect 9781 22049 9815 22083
rect 10701 22049 10735 22083
rect 13277 22049 13311 22083
rect 15209 22049 15243 22083
rect 15393 22049 15427 22083
rect 15577 22049 15611 22083
rect 17233 22049 17267 22083
rect 19349 22049 19383 22083
rect 22937 22049 22971 22083
rect 23029 22049 23063 22083
rect 5549 21981 5583 22015
rect 9137 21981 9171 22015
rect 10057 21981 10091 22015
rect 10425 21981 10459 22015
rect 13737 21981 13771 22015
rect 14289 21981 14323 22015
rect 14657 21981 14691 22015
rect 15117 21981 15151 22015
rect 16129 21981 16163 22015
rect 16313 21981 16347 22015
rect 17601 21981 17635 22015
rect 18429 21981 18463 22015
rect 20269 21981 20303 22015
rect 20453 21981 20487 22015
rect 20637 21981 20671 22015
rect 20729 21981 20763 22015
rect 21097 21981 21131 22015
rect 21925 21981 21959 22015
rect 5825 21913 5859 21947
rect 9689 21913 9723 21947
rect 10241 21913 10275 21947
rect 10333 21913 10367 21947
rect 10977 21913 11011 21947
rect 12541 21913 12575 21947
rect 14381 21913 14415 21947
rect 14473 21913 14507 21947
rect 16957 21913 16991 21947
rect 17785 21913 17819 21947
rect 20177 21913 20211 21947
rect 21557 21913 21591 21947
rect 7297 21845 7331 21879
rect 8953 21845 8987 21879
rect 9229 21845 9263 21879
rect 9597 21845 9631 21879
rect 10609 21845 10643 21879
rect 12449 21845 12483 21879
rect 13921 21845 13955 21879
rect 14105 21845 14139 21879
rect 16497 21845 16531 21879
rect 16589 21845 16623 21879
rect 17049 21845 17083 21879
rect 17417 21845 17451 21879
rect 20361 21845 20395 21879
rect 22845 21845 22879 21879
rect 11529 21641 11563 21675
rect 11897 21641 11931 21675
rect 15853 21641 15887 21675
rect 23213 21641 23247 21675
rect 6377 21573 6411 21607
rect 8585 21573 8619 21607
rect 13553 21573 13587 21607
rect 13645 21573 13679 21607
rect 14289 21573 14323 21607
rect 16957 21573 16991 21607
rect 19717 21573 19751 21607
rect 22293 21573 22327 21607
rect 1777 21505 1811 21539
rect 2789 21505 2823 21539
rect 7113 21505 7147 21539
rect 8309 21505 8343 21539
rect 10701 21505 10735 21539
rect 11989 21505 12023 21539
rect 13277 21505 13311 21539
rect 13370 21505 13404 21539
rect 13742 21505 13776 21539
rect 16405 21505 16439 21539
rect 16681 21505 16715 21539
rect 19441 21505 19475 21539
rect 21925 21505 21959 21539
rect 23765 21505 23799 21539
rect 25697 21505 25731 21539
rect 3065 21437 3099 21471
rect 4813 21437 4847 21471
rect 8033 21437 8067 21471
rect 10057 21437 10091 21471
rect 12173 21437 12207 21471
rect 13093 21437 13127 21471
rect 14013 21437 14047 21471
rect 15761 21437 15795 21471
rect 21189 21437 21223 21471
rect 1501 21301 1535 21335
rect 7389 21301 7423 21335
rect 10149 21301 10183 21335
rect 12541 21301 12575 21335
rect 13921 21301 13955 21335
rect 18429 21301 18463 21335
rect 25881 21301 25915 21335
rect 3157 21097 3191 21131
rect 6193 21097 6227 21131
rect 9137 21097 9171 21131
rect 15853 21097 15887 21131
rect 21649 21097 21683 21131
rect 21998 21097 22032 21131
rect 23489 21097 23523 21131
rect 6377 21029 6411 21063
rect 7113 21029 7147 21063
rect 7665 21029 7699 21063
rect 4445 20961 4479 20995
rect 7849 20961 7883 20995
rect 9689 20961 9723 20995
rect 16497 20961 16531 20995
rect 16773 20961 16807 20995
rect 18245 20961 18279 20995
rect 18889 20961 18923 20995
rect 19533 20961 19567 20995
rect 21741 20961 21775 20995
rect 3341 20893 3375 20927
rect 5549 20893 5583 20927
rect 5825 20893 5859 20927
rect 6009 20893 6043 20927
rect 6561 20893 6595 20927
rect 6745 20893 6779 20927
rect 6883 20893 6917 20927
rect 7021 20893 7055 20927
rect 7573 20893 7607 20927
rect 9505 20893 9539 20927
rect 12541 20893 12575 20927
rect 13737 20893 13771 20927
rect 14105 20893 14139 20927
rect 19257 20893 19291 20927
rect 21465 20893 21499 20927
rect 4169 20825 4203 20859
rect 5687 20825 5721 20859
rect 5917 20825 5951 20859
rect 6653 20825 6687 20859
rect 7297 20825 7331 20859
rect 7481 20825 7515 20859
rect 13277 20825 13311 20859
rect 14381 20825 14415 20859
rect 18337 20825 18371 20859
rect 3801 20757 3835 20791
rect 4261 20757 4295 20791
rect 7849 20757 7883 20791
rect 9597 20757 9631 20791
rect 13921 20757 13955 20791
rect 21005 20757 21039 20791
rect 6745 20553 6779 20587
rect 6929 20553 6963 20587
rect 9413 20553 9447 20587
rect 11989 20553 12023 20587
rect 14841 20553 14875 20587
rect 17049 20553 17083 20587
rect 17509 20553 17543 20587
rect 23305 20553 23339 20587
rect 25237 20553 25271 20587
rect 6377 20485 6411 20519
rect 9781 20485 9815 20519
rect 16037 20485 16071 20519
rect 18337 20485 18371 20519
rect 22017 20485 22051 20519
rect 22753 20485 22787 20519
rect 23213 20485 23247 20519
rect 2329 20417 2363 20451
rect 2605 20417 2639 20451
rect 3249 20417 3283 20451
rect 5089 20417 5123 20451
rect 5917 20417 5951 20451
rect 6101 20417 6135 20451
rect 6193 20417 6227 20451
rect 6561 20417 6595 20451
rect 6837 20417 6871 20451
rect 7021 20417 7055 20451
rect 9321 20417 9355 20451
rect 9873 20417 9907 20451
rect 10333 20417 10367 20451
rect 12081 20417 12115 20451
rect 15853 20417 15887 20451
rect 16129 20417 16163 20451
rect 16221 20417 16255 20451
rect 17141 20417 17175 20451
rect 17601 20417 17635 20451
rect 18613 20417 18647 20451
rect 18706 20417 18740 20451
rect 18889 20417 18923 20451
rect 18981 20417 19015 20451
rect 19097 20417 19131 20451
rect 20637 20417 20671 20451
rect 23857 20417 23891 20451
rect 23949 20417 23983 20451
rect 24041 20417 24075 20451
rect 24225 20417 24259 20451
rect 25053 20417 25087 20451
rect 3341 20349 3375 20383
rect 3525 20349 3559 20383
rect 5181 20349 5215 20383
rect 9965 20349 9999 20383
rect 10885 20349 10919 20383
rect 12265 20349 12299 20383
rect 13093 20349 13127 20383
rect 13369 20349 13403 20383
rect 16957 20349 16991 20383
rect 23397 20349 23431 20383
rect 2881 20281 2915 20315
rect 5457 20281 5491 20315
rect 5733 20281 5767 20315
rect 16405 20281 16439 20315
rect 2145 20213 2179 20247
rect 2421 20213 2455 20247
rect 9137 20213 9171 20247
rect 11621 20213 11655 20247
rect 19257 20213 19291 20247
rect 20913 20213 20947 20247
rect 21097 20213 21131 20247
rect 22845 20213 22879 20247
rect 23673 20213 23707 20247
rect 4445 20009 4479 20043
rect 4905 20009 4939 20043
rect 4997 20009 5031 20043
rect 8033 20009 8067 20043
rect 10701 20009 10735 20043
rect 23305 20009 23339 20043
rect 24961 20009 24995 20043
rect 21833 19941 21867 19975
rect 1869 19873 1903 19907
rect 4537 19873 4571 19907
rect 6193 19873 6227 19907
rect 6285 19873 6319 19907
rect 8953 19873 8987 19907
rect 9229 19873 9263 19907
rect 11161 19873 11195 19907
rect 13461 19873 13495 19907
rect 13553 19873 13587 19907
rect 17877 19873 17911 19907
rect 22477 19873 22511 19907
rect 22753 19873 22787 19907
rect 25053 19873 25087 19907
rect 1593 19805 1627 19839
rect 4261 19805 4295 19839
rect 4445 19805 4479 19839
rect 4721 19805 4755 19839
rect 5181 19805 5215 19839
rect 5365 19805 5399 19839
rect 5457 19805 5491 19839
rect 5733 19805 5767 19839
rect 5917 19805 5951 19839
rect 8769 19805 8803 19839
rect 10885 19805 10919 19839
rect 14657 19805 14691 19839
rect 16865 19805 16899 19839
rect 18889 19805 18923 19839
rect 20913 19805 20947 19839
rect 22293 19805 22327 19839
rect 23397 19805 23431 19839
rect 24409 19805 24443 19839
rect 24685 19805 24719 19839
rect 24961 19805 24995 19839
rect 25237 19805 25271 19839
rect 3617 19737 3651 19771
rect 5825 19737 5859 19771
rect 6055 19737 6089 19771
rect 6561 19737 6595 19771
rect 11437 19737 11471 19771
rect 13369 19737 13403 19771
rect 14105 19737 14139 19771
rect 22201 19737 22235 19771
rect 24869 19737 24903 19771
rect 5549 19669 5583 19703
rect 8585 19669 8619 19703
rect 11069 19669 11103 19703
rect 12909 19669 12943 19703
rect 13001 19669 13035 19703
rect 16313 19669 16347 19703
rect 17325 19669 17359 19703
rect 17693 19669 17727 19703
rect 17785 19669 17819 19703
rect 18337 19669 18371 19703
rect 20729 19669 20763 19703
rect 24041 19669 24075 19703
rect 24501 19669 24535 19703
rect 25421 19669 25455 19703
rect 3709 19465 3743 19499
rect 4077 19465 4111 19499
rect 5273 19465 5307 19499
rect 5733 19465 5767 19499
rect 7113 19465 7147 19499
rect 16497 19465 16531 19499
rect 21649 19465 21683 19499
rect 24409 19465 24443 19499
rect 1869 19397 1903 19431
rect 3617 19397 3651 19431
rect 8677 19397 8711 19431
rect 22845 19397 22879 19431
rect 1593 19329 1627 19363
rect 5457 19329 5491 19363
rect 5641 19329 5675 19363
rect 5917 19329 5951 19363
rect 6101 19329 6135 19363
rect 6193 19329 6227 19363
rect 6377 19329 6411 19363
rect 6469 19329 6503 19363
rect 7757 19329 7791 19363
rect 8401 19329 8435 19363
rect 11161 19329 11195 19363
rect 11529 19329 11563 19363
rect 14749 19329 14783 19363
rect 16865 19329 16899 19363
rect 24225 19329 24259 19363
rect 25053 19329 25087 19363
rect 4169 19261 4203 19295
rect 4261 19261 4295 19295
rect 10149 19261 10183 19295
rect 10793 19261 10827 19295
rect 11805 19261 11839 19295
rect 15025 19261 15059 19295
rect 17141 19261 17175 19295
rect 17417 19261 17451 19295
rect 19165 19261 19199 19295
rect 19901 19261 19935 19295
rect 20177 19261 20211 19295
rect 22109 19261 22143 19295
rect 23489 19261 23523 19295
rect 11345 19193 11379 19227
rect 13277 19193 13311 19227
rect 17049 19193 17083 19227
rect 10241 19125 10275 19159
rect 18889 19125 18923 19159
rect 19809 19125 19843 19159
rect 22937 19125 22971 19159
rect 23673 19125 23707 19159
rect 5181 18921 5215 18955
rect 5733 18921 5767 18955
rect 9321 18921 9355 18955
rect 14933 18921 14967 18955
rect 22201 18921 22235 18955
rect 10977 18853 11011 18887
rect 12541 18853 12575 18887
rect 15577 18853 15611 18887
rect 15669 18853 15703 18887
rect 1593 18785 1627 18819
rect 6009 18785 6043 18819
rect 9873 18785 9907 18819
rect 16221 18785 16255 18819
rect 17141 18785 17175 18819
rect 19717 18785 19751 18819
rect 19809 18785 19843 18819
rect 20453 18785 20487 18819
rect 22385 18785 22419 18819
rect 22753 18785 22787 18819
rect 3617 18717 3651 18751
rect 5365 18717 5399 18751
rect 5549 18717 5583 18751
rect 5641 18717 5675 18751
rect 5733 18717 5767 18751
rect 5825 18717 5859 18751
rect 9689 18717 9723 18751
rect 10425 18717 10459 18751
rect 10609 18717 10643 18751
rect 10793 18717 10827 18751
rect 11897 18717 11931 18751
rect 12045 18717 12079 18751
rect 12403 18717 12437 18751
rect 14749 18717 14783 18751
rect 15025 18717 15059 18751
rect 15393 18717 15427 18751
rect 16037 18717 16071 18751
rect 16497 18717 16531 18751
rect 16865 18717 16899 18751
rect 19625 18717 19659 18751
rect 24179 18717 24213 18751
rect 24593 18717 24627 18751
rect 1869 18649 1903 18683
rect 9781 18649 9815 18683
rect 10701 18649 10735 18683
rect 12173 18649 12207 18683
rect 12265 18649 12299 18683
rect 15209 18649 15243 18683
rect 15301 18649 15335 18683
rect 16681 18649 16715 18683
rect 16773 18649 16807 18683
rect 17417 18649 17451 18683
rect 20729 18649 20763 18683
rect 16129 18581 16163 18615
rect 17049 18581 17083 18615
rect 18889 18581 18923 18615
rect 19257 18581 19291 18615
rect 24501 18581 24535 18615
rect 2237 18377 2271 18411
rect 2697 18377 2731 18411
rect 3525 18377 3559 18411
rect 6929 18377 6963 18411
rect 9505 18377 9539 18411
rect 17417 18377 17451 18411
rect 21005 18377 21039 18411
rect 3065 18309 3099 18343
rect 10609 18309 10643 18343
rect 10701 18309 10735 18343
rect 21557 18309 21591 18343
rect 23397 18309 23431 18343
rect 2421 18241 2455 18275
rect 3157 18241 3191 18275
rect 5365 18241 5399 18275
rect 5549 18241 5583 18275
rect 6561 18241 6595 18275
rect 6653 18241 6687 18275
rect 7757 18241 7791 18275
rect 10241 18241 10275 18275
rect 10425 18241 10459 18275
rect 10793 18241 10827 18275
rect 12265 18241 12299 18275
rect 12403 18241 12437 18275
rect 12541 18241 12575 18275
rect 12633 18241 12667 18275
rect 12730 18241 12764 18275
rect 15853 18241 15887 18275
rect 17601 18241 17635 18275
rect 19809 18241 19843 18275
rect 21189 18241 21223 18275
rect 21281 18241 21315 18275
rect 3341 18173 3375 18207
rect 4169 18173 4203 18207
rect 6469 18173 6503 18207
rect 6745 18173 6779 18207
rect 8033 18173 8067 18207
rect 13369 18173 13403 18207
rect 13645 18173 13679 18207
rect 15117 18173 15151 18207
rect 17233 18173 17267 18207
rect 19533 18173 19567 18207
rect 20453 18173 20487 18207
rect 21649 18173 21683 18207
rect 23673 18173 23707 18207
rect 10977 18105 11011 18139
rect 5549 18037 5583 18071
rect 9689 18037 9723 18071
rect 12909 18037 12943 18071
rect 15301 18037 15335 18071
rect 16681 18037 16715 18071
rect 18061 18037 18095 18071
rect 19901 18037 19935 18071
rect 21925 18037 21959 18071
rect 5733 17833 5767 17867
rect 6193 17833 6227 17867
rect 7665 17833 7699 17867
rect 13645 17833 13679 17867
rect 15853 17833 15887 17867
rect 18797 17833 18831 17867
rect 22109 17833 22143 17867
rect 23765 17833 23799 17867
rect 23949 17833 23983 17867
rect 11345 17765 11379 17799
rect 15945 17765 15979 17799
rect 23029 17765 23063 17799
rect 5181 17697 5215 17731
rect 6837 17697 6871 17731
rect 8309 17697 8343 17731
rect 12081 17697 12115 17731
rect 13185 17697 13219 17731
rect 14105 17697 14139 17731
rect 16497 17697 16531 17731
rect 17877 17697 17911 17731
rect 23121 17697 23155 17731
rect 4997 17629 5031 17663
rect 5273 17629 5307 17663
rect 5365 17629 5399 17663
rect 5457 17629 5491 17663
rect 5825 17629 5859 17663
rect 6009 17629 6043 17663
rect 6377 17629 6411 17663
rect 6469 17629 6503 17663
rect 6561 17629 6595 17663
rect 6653 17629 6687 17663
rect 7205 17629 7239 17663
rect 7573 17629 7607 17663
rect 7849 17629 7883 17663
rect 7941 17629 7975 17663
rect 10885 17629 10919 17663
rect 11161 17629 11195 17663
rect 13461 17629 13495 17663
rect 13737 17629 13771 17663
rect 16313 17629 16347 17663
rect 17049 17629 17083 17663
rect 17197 17629 17231 17663
rect 17514 17629 17548 17663
rect 18153 17629 18187 17663
rect 18613 17629 18647 17663
rect 21649 17629 21683 17663
rect 22017 17629 22051 17663
rect 22293 17629 22327 17663
rect 22385 17629 22419 17663
rect 22477 17629 22511 17663
rect 22661 17629 22695 17663
rect 22845 17629 22879 17663
rect 23857 17629 23891 17663
rect 7389 17561 7423 17595
rect 8033 17561 8067 17595
rect 8171 17561 8205 17595
rect 11805 17561 11839 17595
rect 12633 17561 12667 17595
rect 14381 17561 14415 17595
rect 17325 17561 17359 17595
rect 17417 17561 17451 17595
rect 22753 17561 22787 17595
rect 10241 17493 10275 17527
rect 11437 17493 11471 17527
rect 11897 17493 11931 17527
rect 13921 17493 13955 17527
rect 16405 17493 16439 17527
rect 17693 17493 17727 17527
rect 18061 17493 18095 17527
rect 18521 17493 18555 17527
rect 21833 17493 21867 17527
rect 4629 17289 4663 17323
rect 7113 17289 7147 17323
rect 9781 17289 9815 17323
rect 11069 17289 11103 17323
rect 13277 17289 13311 17323
rect 14289 17289 14323 17323
rect 14749 17289 14783 17323
rect 18429 17289 18463 17323
rect 23305 17289 23339 17323
rect 3617 17221 3651 17255
rect 6561 17221 6595 17255
rect 9689 17221 9723 17255
rect 14657 17221 14691 17255
rect 15669 17221 15703 17255
rect 19961 17221 19995 17255
rect 20177 17221 20211 17255
rect 4169 17153 4203 17187
rect 4461 17153 4495 17187
rect 4997 17153 5031 17187
rect 5365 17153 5399 17187
rect 5549 17153 5583 17187
rect 6193 17153 6227 17187
rect 6377 17153 6411 17187
rect 6837 17153 6871 17187
rect 9045 17153 9079 17187
rect 10333 17153 10367 17187
rect 10977 17153 11011 17187
rect 15577 17153 15611 17187
rect 16681 17153 16715 17187
rect 18521 17153 18555 17187
rect 19073 17153 19107 17187
rect 21373 17153 21407 17187
rect 21557 17153 21591 17187
rect 23949 17153 23983 17187
rect 25973 17153 26007 17187
rect 1593 17085 1627 17119
rect 1869 17085 1903 17119
rect 4261 17085 4295 17119
rect 7113 17077 7147 17111
rect 9873 17085 9907 17119
rect 11253 17085 11287 17119
rect 11529 17085 11563 17119
rect 11805 17085 11839 17119
rect 14933 17085 14967 17119
rect 15853 17085 15887 17119
rect 17233 17085 17267 17119
rect 6929 17017 6963 17051
rect 9321 17017 9355 17051
rect 10609 17017 10643 17051
rect 18797 17017 18831 17051
rect 4445 16949 4479 16983
rect 6193 16949 6227 16983
rect 6745 16949 6779 16983
rect 8861 16949 8895 16983
rect 10517 16949 10551 16983
rect 15209 16949 15243 16983
rect 19809 16949 19843 16983
rect 19993 16949 20027 16983
rect 21557 16949 21591 16983
rect 25789 16949 25823 16983
rect 2145 16745 2179 16779
rect 4813 16745 4847 16779
rect 6101 16745 6135 16779
rect 10701 16745 10735 16779
rect 12541 16745 12575 16779
rect 14657 16745 14691 16779
rect 15282 16745 15316 16779
rect 18429 16745 18463 16779
rect 18613 16745 18647 16779
rect 19349 16745 19383 16779
rect 23581 16745 23615 16779
rect 1501 16609 1535 16643
rect 3341 16609 3375 16643
rect 3985 16609 4019 16643
rect 4353 16609 4387 16643
rect 5457 16609 5491 16643
rect 7021 16609 7055 16643
rect 10793 16609 10827 16643
rect 11069 16609 11103 16643
rect 13185 16609 13219 16643
rect 15025 16609 15059 16643
rect 16773 16609 16807 16643
rect 17325 16609 17359 16643
rect 17417 16609 17451 16643
rect 19993 16609 20027 16643
rect 21189 16609 21223 16643
rect 22109 16609 22143 16643
rect 2329 16541 2363 16575
rect 4169 16541 4203 16575
rect 5181 16541 5215 16575
rect 6101 16541 6135 16575
rect 6285 16541 6319 16575
rect 6561 16541 6595 16575
rect 6745 16541 6779 16575
rect 8585 16541 8619 16575
rect 8953 16541 8987 16575
rect 12633 16541 12667 16575
rect 14473 16541 14507 16575
rect 14933 16541 14967 16575
rect 18245 16541 18279 16575
rect 18981 16541 19015 16575
rect 19809 16541 19843 16575
rect 20729 16541 20763 16575
rect 21097 16541 21131 16575
rect 21833 16541 21867 16575
rect 1777 16473 1811 16507
rect 4445 16473 4479 16507
rect 4629 16473 4663 16507
rect 6653 16473 6687 16507
rect 6883 16473 6917 16507
rect 9229 16473 9263 16507
rect 17233 16473 17267 16507
rect 17693 16473 17727 16507
rect 18613 16473 18647 16507
rect 19625 16473 19659 16507
rect 2697 16405 2731 16439
rect 3065 16405 3099 16439
rect 3157 16405 3191 16439
rect 6009 16405 6043 16439
rect 6377 16405 6411 16439
rect 8769 16405 8803 16439
rect 14749 16405 14783 16439
rect 16865 16405 16899 16439
rect 5641 16201 5675 16235
rect 6929 16201 6963 16235
rect 7665 16201 7699 16235
rect 10149 16201 10183 16235
rect 16313 16201 16347 16235
rect 20821 16201 20855 16235
rect 2973 16133 3007 16167
rect 14841 16133 14875 16167
rect 17877 16133 17911 16167
rect 19625 16133 19659 16167
rect 22109 16133 22143 16167
rect 23857 16133 23891 16167
rect 25513 16133 25547 16167
rect 2237 16065 2271 16099
rect 2513 16065 2547 16099
rect 3065 16065 3099 16099
rect 5365 16065 5399 16099
rect 5549 16065 5583 16099
rect 7573 16065 7607 16099
rect 8401 16065 8435 16099
rect 10793 16065 10827 16099
rect 16681 16065 16715 16099
rect 16829 16065 16863 16099
rect 16957 16065 16991 16099
rect 17049 16065 17083 16099
rect 17187 16065 17221 16099
rect 18245 16065 18279 16099
rect 18429 16065 18463 16099
rect 18889 16065 18923 16099
rect 19165 16097 19199 16131
rect 19717 16065 19751 16099
rect 19901 16065 19935 16099
rect 19993 16065 20027 16099
rect 20913 16065 20947 16099
rect 21833 16065 21867 16099
rect 3249 15997 3283 16031
rect 5089 15997 5123 16031
rect 5457 15997 5491 16031
rect 7849 15997 7883 16031
rect 7941 15997 7975 16031
rect 8033 15997 8067 16031
rect 8125 15997 8159 16031
rect 14565 15997 14599 16031
rect 20177 15997 20211 16031
rect 21649 15997 21683 16031
rect 25789 15997 25823 16031
rect 2605 15929 2639 15963
rect 5181 15929 5215 15963
rect 19165 15929 19199 15963
rect 2053 15861 2087 15895
rect 2329 15861 2363 15895
rect 8664 15861 8698 15895
rect 10241 15861 10275 15895
rect 17325 15861 17359 15895
rect 21005 15861 21039 15895
rect 24041 15861 24075 15895
rect 1856 15657 1890 15691
rect 3801 15657 3835 15691
rect 6929 15657 6963 15691
rect 9229 15657 9263 15691
rect 17049 15657 17083 15691
rect 19257 15657 19291 15691
rect 23213 15657 23247 15691
rect 23489 15657 23523 15691
rect 17233 15589 17267 15623
rect 19993 15589 20027 15623
rect 1593 15521 1627 15555
rect 4353 15521 4387 15555
rect 5181 15521 5215 15555
rect 9781 15521 9815 15555
rect 12541 15521 12575 15555
rect 19533 15521 19567 15555
rect 22293 15521 22327 15555
rect 24409 15521 24443 15555
rect 7021 15453 7055 15487
rect 9597 15453 9631 15487
rect 11529 15453 11563 15487
rect 11897 15453 11931 15487
rect 14105 15453 14139 15487
rect 17325 15453 17359 15487
rect 18521 15453 18555 15487
rect 18613 15453 18647 15487
rect 18890 15453 18924 15487
rect 19073 15453 19107 15487
rect 20177 15453 20211 15487
rect 20361 15453 20395 15487
rect 20453 15453 20487 15487
rect 23673 15453 23707 15487
rect 3617 15385 3651 15419
rect 5457 15385 5491 15419
rect 7297 15385 7331 15419
rect 12449 15385 12483 15419
rect 16865 15385 16899 15419
rect 17693 15385 17727 15419
rect 17877 15385 17911 15419
rect 19993 15385 20027 15419
rect 20729 15385 20763 15419
rect 23029 15385 23063 15419
rect 4169 15317 4203 15351
rect 4261 15317 4295 15351
rect 8769 15317 8803 15351
rect 9689 15317 9723 15351
rect 11345 15317 11379 15351
rect 11713 15317 11747 15351
rect 11989 15317 12023 15351
rect 12357 15317 12391 15351
rect 14289 15317 14323 15351
rect 17075 15317 17109 15351
rect 19441 15317 19475 15351
rect 20269 15317 20303 15351
rect 22201 15317 22235 15351
rect 22937 15317 22971 15351
rect 23229 15317 23263 15351
rect 23397 15317 23431 15351
rect 25053 15317 25087 15351
rect 4169 15113 4203 15147
rect 6469 15113 6503 15147
rect 6929 15113 6963 15147
rect 10977 15113 11011 15147
rect 11345 15113 11379 15147
rect 1869 15045 1903 15079
rect 7481 15045 7515 15079
rect 11805 15045 11839 15079
rect 15301 15045 15335 15079
rect 17937 15045 17971 15079
rect 18153 15045 18187 15079
rect 25513 15045 25547 15079
rect 1593 14977 1627 15011
rect 3617 14977 3651 15011
rect 4077 14977 4111 15011
rect 6377 14977 6411 15011
rect 6653 14977 6687 15011
rect 7205 14977 7239 15011
rect 8861 14977 8895 15011
rect 11529 14977 11563 15011
rect 19993 14977 20027 15011
rect 21189 14977 21223 15011
rect 21373 14977 21407 15011
rect 25789 14977 25823 15011
rect 4261 14909 4295 14943
rect 7113 14909 7147 14943
rect 7573 14909 7607 14943
rect 8217 14909 8251 14943
rect 10793 14909 10827 14943
rect 10885 14909 10919 14943
rect 18245 14909 18279 14943
rect 19717 14909 19751 14943
rect 21281 14909 21315 14943
rect 21465 14909 21499 14943
rect 6653 14841 6687 14875
rect 21005 14841 21039 14875
rect 3709 14773 3743 14807
rect 13277 14773 13311 14807
rect 14013 14773 14047 14807
rect 17785 14773 17819 14807
rect 17969 14773 18003 14807
rect 24041 14773 24075 14807
rect 6929 14569 6963 14603
rect 19809 14569 19843 14603
rect 22753 14569 22787 14603
rect 23397 14569 23431 14603
rect 24593 14569 24627 14603
rect 18705 14501 18739 14535
rect 18797 14501 18831 14535
rect 19349 14501 19383 14535
rect 22937 14501 22971 14535
rect 6561 14433 6595 14467
rect 6653 14433 6687 14467
rect 6745 14433 6779 14467
rect 10793 14433 10827 14467
rect 11253 14433 11287 14467
rect 12725 14433 12759 14467
rect 14381 14433 14415 14467
rect 18337 14433 18371 14467
rect 19901 14433 19935 14467
rect 20361 14433 20395 14467
rect 22109 14433 22143 14467
rect 3157 14365 3191 14399
rect 3525 14365 3559 14399
rect 6469 14365 6503 14399
rect 7941 14365 7975 14399
rect 8125 14365 8159 14399
rect 9689 14365 9723 14399
rect 10057 14365 10091 14399
rect 10977 14365 11011 14399
rect 14105 14365 14139 14399
rect 19717 14365 19751 14399
rect 19809 14365 19843 14399
rect 22385 14365 22419 14399
rect 22477 14365 22511 14399
rect 23121 14365 23155 14399
rect 23213 14365 23247 14399
rect 24593 14365 24627 14399
rect 24685 14365 24719 14399
rect 25053 14365 25087 14399
rect 2789 14297 2823 14331
rect 10609 14297 10643 14331
rect 21833 14297 21867 14331
rect 22845 14297 22879 14331
rect 23581 14297 23615 14331
rect 3341 14229 3375 14263
rect 8309 14229 8343 14263
rect 9505 14229 9539 14263
rect 9873 14229 9907 14263
rect 10149 14229 10183 14263
rect 10517 14229 10551 14263
rect 15853 14229 15887 14263
rect 19257 14229 19291 14263
rect 20177 14229 20211 14263
rect 22201 14229 22235 14263
rect 24961 14229 24995 14263
rect 25697 14229 25731 14263
rect 11529 14025 11563 14059
rect 14105 14025 14139 14059
rect 14473 14025 14507 14059
rect 14565 14025 14599 14059
rect 16681 14025 16715 14059
rect 17141 14025 17175 14059
rect 21189 14025 21223 14059
rect 21931 14025 21965 14059
rect 22201 14025 22235 14059
rect 23949 14025 23983 14059
rect 3065 13957 3099 13991
rect 5549 13957 5583 13991
rect 5917 13957 5951 13991
rect 6009 13957 6043 13991
rect 6469 13957 6503 13991
rect 9229 13957 9263 13991
rect 9873 13957 9907 13991
rect 11897 13957 11931 13991
rect 11989 13957 12023 13991
rect 18061 13957 18095 13991
rect 21557 13957 21591 13991
rect 22017 13957 22051 13991
rect 23581 13957 23615 13991
rect 25421 13957 25455 13991
rect 2789 13889 2823 13923
rect 4997 13889 5031 13923
rect 5825 13889 5859 13923
rect 6193 13889 6227 13923
rect 6377 13889 6411 13923
rect 6555 13889 6589 13923
rect 7205 13889 7239 13923
rect 14933 13889 14967 13923
rect 16405 13889 16439 13923
rect 17049 13889 17083 13923
rect 21097 13889 21131 13923
rect 21281 13889 21315 13923
rect 21373 13889 21407 13923
rect 21649 13889 21683 13923
rect 21833 13889 21867 13923
rect 22109 13889 22143 13923
rect 22385 13889 22419 13923
rect 22845 13889 22879 13923
rect 23765 13889 23799 13923
rect 4813 13821 4847 13855
rect 6929 13821 6963 13855
rect 7021 13821 7055 13855
rect 7389 13821 7423 13855
rect 7757 13821 7791 13855
rect 9505 13821 9539 13855
rect 9597 13821 9631 13855
rect 11345 13821 11379 13855
rect 12173 13821 12207 13855
rect 14657 13821 14691 13855
rect 17325 13821 17359 13855
rect 19809 13821 19843 13855
rect 20085 13821 20119 13855
rect 22477 13821 22511 13855
rect 25697 13821 25731 13855
rect 21373 13753 21407 13787
rect 5641 13685 5675 13719
rect 15025 13685 15059 13719
rect 16221 13685 16255 13719
rect 22753 13685 22787 13719
rect 3893 13481 3927 13515
rect 5917 13481 5951 13515
rect 6837 13481 6871 13515
rect 13921 13481 13955 13515
rect 17785 13481 17819 13515
rect 21741 13481 21775 13515
rect 22293 13481 22327 13515
rect 24225 13481 24259 13515
rect 24409 13481 24443 13515
rect 24869 13481 24903 13515
rect 25053 13481 25087 13515
rect 3157 13413 3191 13447
rect 7205 13413 7239 13447
rect 7389 13413 7423 13447
rect 13185 13413 13219 13447
rect 14933 13413 14967 13447
rect 25881 13413 25915 13447
rect 5365 13345 5399 13379
rect 6561 13345 6595 13379
rect 6745 13345 6779 13379
rect 7573 13345 7607 13379
rect 11989 13345 12023 13379
rect 14657 13345 14691 13379
rect 16313 13345 16347 13379
rect 18521 13345 18555 13379
rect 22477 13345 22511 13379
rect 25145 13345 25179 13379
rect 1409 13277 1443 13311
rect 5641 13277 5675 13311
rect 5825 13277 5859 13311
rect 6101 13277 6135 13311
rect 6469 13277 6503 13311
rect 7021 13277 7055 13311
rect 7297 13277 7331 13311
rect 7849 13277 7883 13311
rect 8217 13277 8251 13311
rect 8769 13277 8803 13311
rect 13185 13277 13219 13311
rect 13369 13277 13403 13311
rect 13737 13277 13771 13311
rect 13921 13277 13955 13311
rect 14381 13277 14415 13311
rect 15393 13277 15427 13311
rect 16037 13277 16071 13311
rect 17969 13277 18003 13311
rect 21925 13277 21959 13311
rect 22109 13277 22143 13311
rect 24685 13277 24719 13311
rect 24961 13277 24995 13311
rect 25329 13277 25363 13311
rect 25697 13277 25731 13311
rect 1685 13209 1719 13243
rect 7665 13209 7699 13243
rect 9045 13209 9079 13243
rect 9413 13209 9447 13243
rect 14197 13209 14231 13243
rect 15209 13209 15243 13243
rect 22385 13209 22419 13243
rect 22753 13209 22787 13243
rect 25053 13209 25087 13243
rect 6285 13141 6319 13175
rect 7573 13141 7607 13175
rect 12633 13141 12667 13175
rect 14565 13141 14599 13175
rect 15117 13141 15151 13175
rect 15577 13141 15611 13175
rect 25513 13141 25547 13175
rect 3157 12937 3191 12971
rect 7573 12937 7607 12971
rect 12173 12937 12207 12971
rect 12541 12937 12575 12971
rect 13185 12937 13219 12971
rect 14565 12937 14599 12971
rect 22477 12937 22511 12971
rect 25237 12937 25271 12971
rect 15393 12869 15427 12903
rect 23765 12869 23799 12903
rect 1409 12801 1443 12835
rect 4261 12801 4295 12835
rect 4353 12801 4387 12835
rect 4537 12801 4571 12835
rect 4813 12801 4847 12835
rect 6561 12801 6595 12835
rect 6837 12801 6871 12835
rect 6929 12801 6963 12835
rect 7113 12801 7147 12835
rect 7941 12801 7975 12835
rect 8033 12801 8067 12835
rect 10885 12801 10919 12835
rect 10977 12801 11011 12835
rect 11253 12801 11287 12835
rect 12081 12801 12115 12835
rect 13369 12801 13403 12835
rect 13645 12801 13679 12835
rect 13829 12801 13863 12835
rect 14004 12801 14038 12835
rect 14105 12801 14139 12835
rect 14381 12801 14415 12835
rect 14657 12801 14691 12835
rect 14933 12801 14967 12835
rect 15117 12801 15151 12835
rect 15485 12801 15519 12835
rect 15577 12801 15611 12835
rect 15945 12801 15979 12835
rect 16221 12801 16255 12835
rect 16405 12801 16439 12835
rect 19901 12801 19935 12835
rect 19993 12801 20027 12835
rect 23489 12801 23523 12835
rect 1685 12733 1719 12767
rect 5549 12733 5583 12767
rect 7849 12733 7883 12767
rect 8309 12733 8343 12767
rect 11161 12733 11195 12767
rect 12633 12733 12667 12767
rect 12725 12733 12759 12767
rect 15761 12733 15795 12767
rect 16313 12733 16347 12767
rect 16957 12733 16991 12767
rect 17233 12733 17267 12767
rect 18705 12733 18739 12767
rect 19349 12733 19383 12767
rect 23029 12733 23063 12767
rect 6745 12665 6779 12699
rect 9781 12665 9815 12699
rect 15945 12665 15979 12699
rect 4721 12597 4755 12631
rect 6377 12597 6411 12631
rect 7021 12597 7055 12631
rect 7757 12597 7791 12631
rect 10701 12597 10735 12631
rect 11897 12597 11931 12631
rect 18797 12597 18831 12631
rect 20177 12597 20211 12631
rect 1593 12393 1627 12427
rect 8953 12393 8987 12427
rect 12633 12393 12667 12427
rect 13369 12393 13403 12427
rect 15577 12393 15611 12427
rect 17325 12393 17359 12427
rect 22201 12393 22235 12427
rect 6653 12325 6687 12359
rect 4353 12257 4387 12291
rect 4721 12257 4755 12291
rect 9597 12257 9631 12291
rect 10517 12257 10551 12291
rect 12541 12257 12575 12291
rect 13185 12257 13219 12291
rect 15117 12257 15151 12291
rect 18061 12257 18095 12291
rect 18153 12257 18187 12291
rect 1409 12189 1443 12223
rect 1777 12189 1811 12223
rect 5549 12189 5583 12223
rect 6193 12189 6227 12223
rect 6285 12189 6319 12223
rect 6561 12189 6595 12223
rect 6837 12189 6871 12223
rect 6929 12189 6963 12223
rect 7021 12189 7055 12223
rect 7205 12189 7239 12223
rect 9078 12189 9112 12223
rect 9505 12189 9539 12223
rect 13553 12189 13587 12223
rect 13645 12189 13679 12223
rect 13921 12189 13955 12223
rect 14105 12189 14139 12223
rect 14289 12189 14323 12223
rect 14555 12167 14589 12201
rect 14657 12189 14691 12223
rect 14841 12189 14875 12223
rect 14933 12189 14967 12223
rect 15209 12189 15243 12223
rect 17509 12189 17543 12223
rect 17969 12189 18003 12223
rect 20177 12189 20211 12223
rect 20453 12189 20487 12223
rect 2053 12121 2087 12155
rect 4169 12121 4203 12155
rect 6377 12121 6411 12155
rect 10793 12121 10827 12155
rect 13737 12121 13771 12155
rect 20729 12121 20763 12155
rect 3525 12053 3559 12087
rect 3801 12053 3835 12087
rect 4261 12053 4295 12087
rect 6009 12053 6043 12087
rect 9137 12053 9171 12087
rect 14473 12053 14507 12087
rect 15577 12053 15611 12087
rect 15761 12053 15795 12087
rect 17601 12053 17635 12087
rect 19625 12053 19659 12087
rect 2697 11849 2731 11883
rect 5641 11849 5675 11883
rect 14381 11849 14415 11883
rect 15669 11849 15703 11883
rect 24961 11849 24995 11883
rect 25237 11849 25271 11883
rect 4537 11781 4571 11815
rect 10425 11781 10459 11815
rect 11161 11781 11195 11815
rect 11897 11781 11931 11815
rect 13737 11781 13771 11815
rect 13921 11781 13955 11815
rect 14565 11781 14599 11815
rect 2881 11713 2915 11747
rect 4813 11713 4847 11747
rect 5825 11713 5859 11747
rect 5917 11713 5951 11747
rect 6193 11713 6227 11747
rect 6469 11713 6503 11747
rect 6561 11713 6595 11747
rect 6745 11713 6779 11747
rect 9873 11713 9907 11747
rect 10057 11713 10091 11747
rect 10333 11711 10367 11745
rect 11621 11713 11655 11747
rect 13645 11713 13679 11747
rect 14289 11713 14323 11747
rect 14933 11713 14967 11747
rect 15025 11713 15059 11747
rect 15301 11713 15335 11747
rect 15393 11713 15427 11747
rect 15761 11713 15795 11747
rect 15945 11713 15979 11747
rect 18429 11713 18463 11747
rect 20361 11713 20395 11747
rect 21281 11713 21315 11747
rect 21465 11713 21499 11747
rect 21833 11713 21867 11747
rect 22109 11713 22143 11747
rect 23213 11713 23247 11747
rect 25053 11713 25087 11747
rect 4905 11645 4939 11679
rect 5549 11645 5583 11679
rect 13369 11645 13403 11679
rect 15669 11645 15703 11679
rect 18705 11645 18739 11679
rect 20821 11645 20855 11679
rect 21097 11645 21131 11679
rect 23489 11645 23523 11679
rect 9873 11577 9907 11611
rect 13921 11577 13955 11611
rect 15485 11577 15519 11611
rect 3065 11509 3099 11543
rect 6101 11509 6135 11543
rect 6745 11509 6779 11543
rect 10241 11509 10275 11543
rect 14565 11509 14599 11543
rect 15853 11509 15887 11543
rect 20177 11509 20211 11543
rect 22017 11509 22051 11543
rect 22293 11509 22327 11543
rect 6285 11305 6319 11339
rect 7941 11305 7975 11339
rect 8953 11305 8987 11339
rect 10885 11305 10919 11339
rect 18613 11305 18647 11339
rect 24409 11305 24443 11339
rect 25329 11305 25363 11339
rect 6653 11237 6687 11271
rect 7205 11237 7239 11271
rect 25145 11237 25179 11271
rect 5641 11169 5675 11203
rect 6101 11169 6135 11203
rect 6561 11169 6595 11203
rect 8125 11169 8159 11203
rect 11345 11169 11379 11203
rect 11621 11169 11655 11203
rect 11897 11169 11931 11203
rect 14749 11169 14783 11203
rect 17969 11169 18003 11203
rect 19257 11169 19291 11203
rect 21097 11169 21131 11203
rect 22845 11169 22879 11203
rect 23673 11169 23707 11203
rect 3065 11101 3099 11135
rect 5825 11101 5859 11135
rect 5917 11101 5951 11135
rect 6009 11101 6043 11135
rect 6469 11101 6503 11135
rect 6745 11101 6779 11135
rect 7573 11101 7607 11135
rect 8217 11101 8251 11135
rect 9137 11101 9171 11135
rect 9229 11101 9263 11135
rect 9505 11101 9539 11135
rect 9597 11101 9631 11135
rect 10793 11101 10827 11135
rect 11069 11101 11103 11135
rect 11161 11101 11195 11135
rect 11437 11101 11471 11135
rect 14473 11101 14507 11135
rect 14565 11101 14599 11135
rect 17233 11101 17267 11135
rect 18797 11101 18831 11135
rect 18981 11101 19015 11135
rect 19073 11101 19107 11135
rect 24961 11101 24995 11135
rect 25697 11101 25731 11135
rect 9321 11033 9355 11067
rect 10057 11033 10091 11067
rect 13645 11033 13679 11067
rect 14749 11033 14783 11067
rect 19533 11033 19567 11067
rect 22569 11033 22603 11067
rect 22937 11033 22971 11067
rect 3617 10965 3651 10999
rect 7113 10965 7147 10999
rect 17049 10965 17083 10999
rect 17325 10965 17359 10999
rect 21005 10965 21039 10999
rect 25329 10965 25363 10999
rect 6377 10761 6411 10795
rect 6745 10761 6779 10795
rect 7097 10761 7131 10795
rect 8953 10761 8987 10795
rect 9597 10761 9631 10795
rect 11069 10761 11103 10795
rect 16681 10761 16715 10795
rect 17049 10761 17083 10795
rect 17509 10761 17543 10795
rect 19349 10761 19383 10795
rect 20177 10761 20211 10795
rect 1501 10693 1535 10727
rect 3249 10693 3283 10727
rect 4077 10693 4111 10727
rect 7297 10693 7331 10727
rect 8769 10693 8803 10727
rect 17141 10693 17175 10727
rect 17969 10693 18003 10727
rect 19717 10693 19751 10727
rect 20821 10693 20855 10727
rect 3525 10625 3559 10659
rect 3893 10625 3927 10659
rect 5825 10625 5859 10659
rect 5917 10625 5951 10659
rect 6561 10625 6595 10659
rect 6837 10625 6871 10659
rect 7389 10625 7423 10659
rect 7573 10625 7607 10659
rect 8585 10625 8619 10659
rect 8861 10625 8895 10659
rect 9137 10625 9171 10659
rect 9965 10625 9999 10659
rect 10057 10625 10091 10659
rect 10425 10625 10459 10659
rect 10609 10625 10643 10659
rect 10701 10625 10735 10659
rect 10793 10625 10827 10659
rect 16313 10625 16347 10659
rect 17877 10625 17911 10659
rect 19073 10625 19107 10659
rect 19257 10625 19291 10659
rect 19533 10625 19567 10659
rect 19809 10625 19843 10659
rect 20361 10625 20395 10659
rect 20729 10625 20763 10659
rect 22017 10625 22051 10659
rect 22201 10625 22235 10659
rect 3617 10557 3651 10591
rect 5641 10557 5675 10591
rect 5733 10557 5767 10591
rect 10149 10557 10183 10591
rect 17325 10557 17359 10591
rect 18061 10557 18095 10591
rect 19165 10557 19199 10591
rect 19901 10557 19935 10591
rect 20085 10557 20119 10591
rect 21373 10557 21407 10591
rect 22477 10557 22511 10591
rect 24225 10557 24259 10591
rect 24501 10557 24535 10591
rect 25237 10557 25271 10591
rect 25789 10557 25823 10591
rect 9137 10489 9171 10523
rect 3709 10421 3743 10455
rect 5457 10421 5491 10455
rect 6929 10421 6963 10455
rect 7113 10421 7147 10455
rect 7573 10421 7607 10455
rect 8401 10421 8435 10455
rect 16129 10421 16163 10455
rect 21833 10421 21867 10455
rect 25145 10421 25179 10455
rect 5917 10217 5951 10251
rect 6101 10217 6135 10251
rect 6653 10217 6687 10251
rect 7941 10217 7975 10251
rect 8401 10217 8435 10251
rect 9045 10217 9079 10251
rect 9873 10217 9907 10251
rect 10609 10217 10643 10251
rect 15932 10217 15966 10251
rect 20164 10217 20198 10251
rect 22201 10217 22235 10251
rect 22477 10217 22511 10251
rect 25421 10217 25455 10251
rect 2881 10081 2915 10115
rect 4905 10081 4939 10115
rect 5549 10081 5583 10115
rect 5733 10081 5767 10115
rect 6745 10081 6779 10115
rect 9689 10081 9723 10115
rect 14565 10081 14599 10115
rect 14749 10081 14783 10115
rect 15669 10081 15703 10115
rect 19901 10081 19935 10115
rect 2605 10013 2639 10047
rect 2789 10013 2823 10047
rect 3801 10013 3835 10047
rect 3985 10013 4019 10047
rect 4261 10013 4295 10047
rect 5457 10013 5491 10047
rect 5641 10013 5675 10047
rect 6377 10013 6411 10047
rect 6469 10013 6503 10047
rect 7941 10013 7975 10047
rect 8125 10013 8159 10047
rect 8401 10013 8435 10047
rect 8769 10013 8803 10047
rect 8953 10013 8987 10047
rect 9137 10013 9171 10047
rect 9413 10013 9447 10047
rect 9505 10013 9539 10047
rect 9781 10013 9815 10047
rect 10057 10013 10091 10047
rect 10149 10013 10183 10047
rect 10333 10013 10367 10047
rect 10425 10013 10459 10047
rect 10517 10013 10551 10047
rect 10701 10013 10735 10047
rect 10793 10013 10827 10047
rect 14933 10013 14967 10047
rect 21833 10013 21867 10047
rect 22017 10013 22051 10047
rect 24225 10013 24259 10047
rect 25145 10013 25179 10047
rect 25605 10013 25639 10047
rect 25881 10013 25915 10047
rect 4445 9945 4479 9979
rect 4537 9945 4571 9979
rect 4721 9945 4755 9979
rect 6009 9945 6043 9979
rect 6929 9945 6963 9979
rect 7113 9945 7147 9979
rect 23949 9945 23983 9979
rect 24409 9945 24443 9979
rect 25789 9945 25823 9979
rect 2421 9877 2455 9911
rect 8585 9877 8619 9911
rect 9229 9877 9263 9911
rect 14105 9877 14139 9911
rect 14473 9877 14507 9911
rect 15117 9877 15151 9911
rect 17417 9877 17451 9911
rect 21649 9877 21683 9911
rect 8677 9673 8711 9707
rect 9137 9673 9171 9707
rect 10149 9673 10183 9707
rect 10701 9673 10735 9707
rect 10885 9673 10919 9707
rect 14841 9673 14875 9707
rect 23443 9673 23477 9707
rect 25881 9673 25915 9707
rect 2329 9605 2363 9639
rect 3249 9605 3283 9639
rect 3893 9605 3927 9639
rect 4353 9605 4387 9639
rect 9965 9605 9999 9639
rect 15301 9605 15335 9639
rect 16957 9605 16991 9639
rect 20821 9605 20855 9639
rect 2053 9537 2087 9571
rect 2973 9537 3007 9571
rect 4077 9537 4111 9571
rect 4169 9537 4203 9571
rect 4445 9537 4479 9571
rect 4537 9537 4571 9571
rect 4721 9537 4755 9571
rect 6745 9537 6779 9571
rect 8493 9537 8527 9571
rect 8677 9537 8711 9571
rect 8861 9537 8895 9571
rect 9689 9537 9723 9571
rect 9781 9537 9815 9571
rect 10333 9537 10367 9571
rect 10793 9537 10827 9571
rect 10885 9537 10919 9571
rect 11062 9537 11096 9571
rect 11149 9537 11183 9571
rect 11345 9537 11379 9571
rect 12725 9537 12759 9571
rect 15209 9537 15243 9571
rect 16681 9537 16715 9571
rect 24869 9537 24903 9571
rect 25237 9537 25271 9571
rect 25421 9537 25455 9571
rect 2329 9469 2363 9503
rect 2697 9469 2731 9503
rect 6653 9469 6687 9503
rect 8953 9469 8987 9503
rect 9137 9469 9171 9503
rect 9965 9469 9999 9503
rect 10517 9469 10551 9503
rect 13001 9469 13035 9503
rect 14749 9469 14783 9503
rect 15485 9469 15519 9503
rect 18613 9469 18647 9503
rect 19901 9469 19935 9503
rect 20637 9469 20671 9503
rect 21373 9469 21407 9503
rect 22385 9469 22419 9503
rect 2789 9401 2823 9435
rect 3617 9401 3651 9435
rect 4169 9401 4203 9435
rect 6377 9401 6411 9435
rect 11161 9401 11195 9435
rect 19349 9401 19383 9435
rect 2145 9333 2179 9367
rect 2881 9333 2915 9367
rect 3065 9333 3099 9367
rect 3249 9333 3283 9367
rect 3709 9333 3743 9367
rect 4721 9333 4755 9367
rect 6561 9333 6595 9367
rect 18429 9333 18463 9367
rect 19257 9333 19291 9367
rect 20085 9333 20119 9367
rect 21833 9333 21867 9367
rect 25697 9333 25731 9367
rect 5641 9129 5675 9163
rect 6745 9129 6779 9163
rect 10149 9129 10183 9163
rect 13277 9129 13311 9163
rect 7481 9061 7515 9095
rect 8217 9061 8251 9095
rect 1685 8993 1719 9027
rect 3433 8993 3467 9027
rect 4445 8993 4479 9027
rect 7665 8993 7699 9027
rect 11897 8993 11931 9027
rect 14197 8993 14231 9027
rect 15669 8993 15703 9027
rect 15945 8993 15979 9027
rect 16681 8993 16715 9027
rect 16773 8993 16807 9027
rect 18429 8993 18463 9027
rect 18613 8993 18647 9027
rect 20177 8993 20211 9027
rect 22293 8993 22327 9027
rect 1409 8925 1443 8959
rect 3801 8925 3835 8959
rect 3985 8925 4019 8959
rect 4261 8925 4295 8959
rect 4721 8925 4755 8959
rect 4813 8925 4847 8959
rect 5089 8925 5123 8959
rect 5273 8925 5307 8959
rect 5549 8925 5583 8959
rect 6653 8925 6687 8959
rect 6837 8925 6871 8959
rect 7481 8925 7515 8959
rect 7757 8925 7791 8959
rect 7941 8925 7975 8959
rect 8309 8925 8343 8959
rect 10057 8925 10091 8959
rect 10241 8925 10275 8959
rect 13461 8925 13495 8959
rect 18061 8925 18095 8959
rect 4537 8857 4571 8891
rect 5457 8857 5491 8891
rect 7113 8857 7147 8891
rect 17325 8857 17359 8891
rect 20453 8857 20487 8891
rect 22569 8857 22603 8891
rect 11253 8789 11287 8823
rect 11621 8789 11655 8823
rect 11713 8789 11747 8823
rect 16865 8789 16899 8823
rect 17233 8789 17267 8823
rect 18705 8789 18739 8823
rect 19073 8789 19107 8823
rect 21925 8789 21959 8823
rect 24041 8789 24075 8823
rect 1593 8585 1627 8619
rect 2605 8585 2639 8619
rect 7573 8585 7607 8619
rect 8217 8585 8251 8619
rect 10885 8585 10919 8619
rect 11621 8585 11655 8619
rect 20729 8585 20763 8619
rect 21833 8585 21867 8619
rect 23765 8585 23799 8619
rect 25605 8585 25639 8619
rect 5917 8517 5951 8551
rect 6009 8517 6043 8551
rect 7849 8517 7883 8551
rect 13093 8517 13127 8551
rect 16313 8517 16347 8551
rect 18153 8517 18187 8551
rect 19993 8517 20027 8551
rect 21189 8517 21223 8551
rect 1409 8449 1443 8483
rect 2053 8449 2087 8483
rect 2145 8449 2179 8483
rect 2421 8449 2455 8483
rect 2693 8449 2727 8483
rect 2881 8449 2915 8483
rect 3157 8449 3191 8483
rect 3341 8449 3375 8483
rect 3617 8449 3651 8483
rect 3893 8449 3927 8483
rect 3985 8449 4019 8483
rect 4169 8449 4203 8483
rect 4261 8449 4295 8483
rect 4905 8449 4939 8483
rect 5089 8449 5123 8483
rect 5820 8449 5854 8483
rect 6193 8449 6227 8483
rect 7757 8449 7791 8483
rect 7941 8449 7975 8483
rect 8125 8449 8159 8483
rect 8585 8449 8619 8483
rect 10517 8449 10551 8483
rect 11069 8449 11103 8483
rect 11713 8449 11747 8483
rect 12081 8449 12115 8483
rect 12357 8449 12391 8483
rect 12725 8449 12759 8483
rect 12909 8449 12943 8483
rect 13185 8449 13219 8483
rect 14197 8449 14231 8483
rect 14933 8449 14967 8483
rect 15853 8449 15887 8483
rect 16129 8449 16163 8483
rect 16497 8449 16531 8483
rect 16957 8449 16991 8483
rect 17417 8449 17451 8483
rect 20913 8449 20947 8483
rect 23857 8449 23891 8483
rect 2329 8381 2363 8415
rect 3525 8381 3559 8415
rect 4813 8381 4847 8415
rect 5917 8381 5951 8415
rect 6653 8381 6687 8415
rect 7389 8381 7423 8415
rect 8493 8381 8527 8415
rect 10425 8381 10459 8415
rect 11345 8381 11379 8415
rect 16037 8381 16071 8415
rect 18245 8381 18279 8415
rect 20269 8381 20303 8415
rect 21097 8381 21131 8415
rect 22385 8381 22419 8415
rect 23213 8381 23247 8415
rect 24133 8381 24167 8415
rect 2237 8313 2271 8347
rect 4353 8313 4387 8347
rect 4445 8313 4479 8347
rect 4905 8313 4939 8347
rect 15669 8313 15703 8347
rect 2421 8245 2455 8279
rect 3709 8245 3743 8279
rect 8401 8245 8435 8279
rect 11161 8245 11195 8279
rect 11253 8245 11287 8279
rect 13277 8245 13311 8279
rect 17141 8245 17175 8279
rect 21189 8245 21223 8279
rect 2881 8041 2915 8075
rect 5549 8041 5583 8075
rect 7481 8041 7515 8075
rect 10885 8041 10919 8075
rect 22477 8041 22511 8075
rect 7665 7973 7699 8007
rect 7941 7973 7975 8007
rect 14105 7973 14139 8007
rect 4997 7905 5031 7939
rect 11345 7905 11379 7939
rect 12633 7905 12667 7939
rect 12909 7905 12943 7939
rect 14381 7905 14415 7939
rect 15301 7905 15335 7939
rect 16589 7905 16623 7939
rect 17049 7905 17083 7939
rect 19901 7905 19935 7939
rect 21649 7905 21683 7939
rect 21925 7905 21959 7939
rect 24961 7905 24995 7939
rect 25697 7905 25731 7939
rect 25973 7905 26007 7939
rect 2881 7837 2915 7871
rect 3065 7837 3099 7871
rect 3801 7837 3835 7871
rect 3985 7837 4019 7871
rect 5181 7837 5215 7871
rect 5825 7837 5859 7871
rect 6101 7837 6135 7871
rect 6469 7837 6503 7871
rect 6837 7837 6871 7871
rect 7389 7837 7423 7871
rect 7573 7837 7607 7871
rect 7941 7837 7975 7871
rect 8125 7837 8159 7871
rect 11069 7837 11103 7871
rect 11253 7837 11287 7871
rect 11437 7837 11471 7871
rect 12265 7837 12299 7871
rect 12449 7837 12483 7871
rect 13001 7837 13035 7871
rect 14473 7837 14507 7871
rect 15669 7837 15703 7871
rect 16037 7837 16071 7871
rect 16497 7837 16531 7871
rect 16681 7837 16715 7871
rect 19441 7837 19475 7871
rect 22293 7837 22327 7871
rect 22385 7837 22419 7871
rect 5089 7769 5123 7803
rect 17325 7769 17359 7803
rect 19073 7769 19107 7803
rect 22017 7769 22051 7803
rect 3985 7701 4019 7735
rect 19257 7701 19291 7735
rect 22109 7701 22143 7735
rect 24409 7701 24443 7735
rect 7021 7497 7055 7531
rect 8769 7497 8803 7531
rect 11713 7497 11747 7531
rect 15485 7497 15519 7531
rect 17509 7497 17543 7531
rect 20729 7497 20763 7531
rect 21097 7497 21131 7531
rect 25421 7497 25455 7531
rect 7205 7429 7239 7463
rect 9413 7429 9447 7463
rect 13093 7429 13127 7463
rect 18981 7429 19015 7463
rect 23305 7429 23339 7463
rect 23949 7429 23983 7463
rect 6377 7361 6411 7395
rect 6837 7361 6871 7395
rect 7389 7361 7423 7395
rect 8677 7361 8711 7395
rect 8861 7361 8895 7395
rect 9321 7361 9355 7395
rect 9505 7361 9539 7395
rect 11713 7361 11747 7395
rect 11897 7361 11931 7395
rect 12173 7361 12207 7395
rect 12633 7361 12667 7395
rect 13461 7361 13495 7395
rect 14749 7361 14783 7395
rect 15117 7361 15151 7395
rect 15669 7361 15703 7395
rect 15853 7361 15887 7395
rect 17325 7361 17359 7395
rect 20913 7361 20947 7395
rect 21189 7361 21223 7395
rect 6469 7293 6503 7327
rect 6653 7293 6687 7327
rect 14657 7293 14691 7327
rect 15761 7293 15795 7327
rect 15945 7293 15979 7327
rect 19257 7293 19291 7327
rect 23581 7293 23615 7327
rect 23673 7293 23707 7327
rect 11989 7157 12023 7191
rect 13921 7157 13955 7191
rect 15025 7157 15059 7191
rect 15301 7157 15335 7191
rect 16681 7157 16715 7191
rect 21833 7157 21867 7191
rect 5917 6953 5951 6987
rect 7021 6953 7055 6987
rect 11148 6953 11182 6987
rect 13093 6953 13127 6987
rect 13829 6953 13863 6987
rect 21557 6953 21591 6987
rect 21741 6953 21775 6987
rect 24133 6953 24167 6987
rect 24409 6953 24443 6987
rect 25145 6953 25179 6987
rect 12633 6885 12667 6919
rect 14381 6885 14415 6919
rect 22385 6885 22419 6919
rect 2605 6817 2639 6851
rect 6377 6817 6411 6851
rect 10885 6817 10919 6851
rect 15117 6817 15151 6851
rect 15577 6817 15611 6851
rect 16313 6817 16347 6851
rect 16681 6817 16715 6851
rect 17049 6817 17083 6851
rect 23029 6817 23063 6851
rect 24501 6817 24535 6851
rect 25697 6817 25731 6851
rect 2421 6749 2455 6783
rect 2697 6749 2731 6783
rect 2973 6749 3007 6783
rect 3525 6749 3559 6783
rect 6101 6749 6135 6783
rect 6285 6749 6319 6783
rect 8309 6749 8343 6783
rect 8493 6749 8527 6783
rect 9413 6749 9447 6783
rect 9597 6749 9631 6783
rect 9873 6749 9907 6783
rect 12909 6749 12943 6783
rect 13093 6749 13127 6783
rect 13737 6749 13771 6783
rect 13921 6749 13955 6783
rect 14105 6749 14139 6783
rect 14841 6749 14875 6783
rect 16865 6749 16899 6783
rect 17417 6749 17451 6783
rect 17601 6749 17635 6783
rect 18797 6749 18831 6783
rect 21649 6749 21683 6783
rect 21925 6749 21959 6783
rect 22090 6749 22124 6783
rect 22201 6749 22235 6783
rect 22293 6749 22327 6783
rect 23489 6749 23523 6783
rect 24409 6749 24443 6783
rect 9229 6681 9263 6715
rect 2237 6613 2271 6647
rect 9689 6613 9723 6647
rect 17417 6613 17451 6647
rect 18613 6613 18647 6647
rect 21189 6613 21223 6647
rect 24777 6613 24811 6647
rect 6193 6409 6227 6443
rect 6561 6409 6595 6443
rect 7941 6409 7975 6443
rect 8585 6409 8619 6443
rect 11989 6409 12023 6443
rect 12449 6409 12483 6443
rect 13185 6409 13219 6443
rect 13737 6409 13771 6443
rect 16957 6409 16991 6443
rect 20085 6409 20119 6443
rect 1685 6341 1719 6375
rect 9321 6341 9355 6375
rect 12081 6341 12115 6375
rect 18061 6341 18095 6375
rect 1409 6273 1443 6307
rect 5549 6273 5583 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 7757 6273 7791 6307
rect 8033 6273 8067 6307
rect 8125 6273 8159 6307
rect 9045 6273 9079 6307
rect 13369 6273 13403 6307
rect 13553 6273 13587 6307
rect 13645 6273 13679 6307
rect 13829 6273 13863 6307
rect 14197 6273 14231 6307
rect 14657 6273 14691 6307
rect 14933 6273 14967 6307
rect 15301 6273 15335 6307
rect 15393 6273 15427 6307
rect 17141 6273 17175 6307
rect 17233 6273 17267 6307
rect 17509 6273 17543 6307
rect 18337 6273 18371 6307
rect 21649 6273 21683 6307
rect 23581 6273 23615 6307
rect 25421 6273 25455 6307
rect 5273 6205 5307 6239
rect 6929 6205 6963 6239
rect 11897 6205 11931 6239
rect 14473 6205 14507 6239
rect 17417 6205 17451 6239
rect 18613 6205 18647 6239
rect 23305 6205 23339 6239
rect 25145 6205 25179 6239
rect 17601 6137 17635 6171
rect 17693 6137 17727 6171
rect 23673 6137 23707 6171
rect 3157 6069 3191 6103
rect 7573 6069 7607 6103
rect 8401 6069 8435 6103
rect 10793 6069 10827 6103
rect 14289 6069 14323 6103
rect 14841 6069 14875 6103
rect 15025 6069 15059 6103
rect 15577 6069 15611 6103
rect 21557 6069 21591 6103
rect 21833 6069 21867 6103
rect 5273 5865 5307 5899
rect 6745 5865 6779 5899
rect 8217 5865 8251 5899
rect 8953 5865 8987 5899
rect 9137 5865 9171 5899
rect 10149 5865 10183 5899
rect 11621 5865 11655 5899
rect 13277 5865 13311 5899
rect 15945 5865 15979 5899
rect 19257 5865 19291 5899
rect 22753 5865 22787 5899
rect 11437 5797 11471 5831
rect 15393 5797 15427 5831
rect 4997 5729 5031 5763
rect 5549 5729 5583 5763
rect 6469 5729 6503 5763
rect 7573 5729 7607 5763
rect 9965 5729 9999 5763
rect 10609 5729 10643 5763
rect 10701 5729 10735 5763
rect 11713 5729 11747 5763
rect 13093 5729 13127 5763
rect 18086 5729 18120 5763
rect 18521 5729 18555 5763
rect 18613 5729 18647 5763
rect 19717 5729 19751 5763
rect 19809 5729 19843 5763
rect 22201 5729 22235 5763
rect 22477 5729 22511 5763
rect 4905 5661 4939 5695
rect 5825 5661 5859 5695
rect 6561 5661 6595 5695
rect 6745 5661 6779 5695
rect 7088 5661 7122 5695
rect 8401 5661 8435 5695
rect 8677 5661 8711 5695
rect 9873 5661 9907 5695
rect 11805 5661 11839 5695
rect 13369 5661 13403 5695
rect 15577 5661 15611 5695
rect 15853 5661 15887 5695
rect 16037 5661 16071 5695
rect 17601 5661 17635 5695
rect 17969 5661 18003 5695
rect 23029 5661 23063 5695
rect 7205 5593 7239 5627
rect 9321 5593 9355 5627
rect 15761 5593 15795 5627
rect 19625 5593 19659 5627
rect 20453 5593 20487 5627
rect 6929 5525 6963 5559
rect 7297 5525 7331 5559
rect 8585 5525 8619 5559
rect 9121 5525 9155 5559
rect 9505 5525 9539 5559
rect 10517 5525 10551 5559
rect 12817 5525 12851 5559
rect 17877 5525 17911 5559
rect 18245 5525 18279 5559
rect 18705 5525 18739 5559
rect 19073 5525 19107 5559
rect 22569 5525 22603 5559
rect 4813 5321 4847 5355
rect 5549 5321 5583 5355
rect 5641 5321 5675 5355
rect 6009 5321 6043 5355
rect 8125 5321 8159 5355
rect 9045 5321 9079 5355
rect 17601 5321 17635 5355
rect 18153 5321 18187 5355
rect 20361 5321 20395 5355
rect 23489 5321 23523 5355
rect 6745 5253 6779 5287
rect 18245 5253 18279 5287
rect 18429 5253 18463 5287
rect 4721 5185 4755 5219
rect 4899 5185 4933 5219
rect 5181 5185 5215 5219
rect 5825 5185 5859 5219
rect 6101 5185 6135 5219
rect 7481 5185 7515 5219
rect 8125 5185 8159 5219
rect 8309 5185 8343 5219
rect 9137 5185 9171 5219
rect 9321 5185 9355 5219
rect 9597 5185 9631 5219
rect 9689 5183 9723 5217
rect 13185 5185 13219 5219
rect 13277 5185 13311 5219
rect 13461 5185 13495 5219
rect 16129 5185 16163 5219
rect 17049 5185 17083 5219
rect 17141 5185 17175 5219
rect 17325 5185 17359 5219
rect 17417 5185 17451 5219
rect 17785 5185 17819 5219
rect 17969 5185 18003 5219
rect 18061 5185 18095 5219
rect 18153 5185 18187 5219
rect 5273 5117 5307 5151
rect 13093 5117 13127 5151
rect 16037 5117 16071 5151
rect 18613 5117 18647 5151
rect 18889 5117 18923 5151
rect 22845 5117 22879 5151
rect 8861 4981 8895 5015
rect 12817 4981 12851 5015
rect 13001 4981 13035 5015
rect 13369 4981 13403 5015
rect 16865 4981 16899 5015
rect 5825 4777 5859 4811
rect 6101 4777 6135 4811
rect 7021 4777 7055 4811
rect 9045 4777 9079 4811
rect 9505 4777 9539 4811
rect 16589 4777 16623 4811
rect 18889 4777 18923 4811
rect 9321 4641 9355 4675
rect 9781 4641 9815 4675
rect 9965 4641 9999 4675
rect 10609 4641 10643 4675
rect 12909 4641 12943 4675
rect 13645 4641 13679 4675
rect 16129 4641 16163 4675
rect 16957 4641 16991 4675
rect 1777 4573 1811 4607
rect 5733 4573 5767 4607
rect 5917 4573 5951 4607
rect 6009 4583 6043 4617
rect 6193 4573 6227 4607
rect 6929 4573 6963 4607
rect 7113 4573 7147 4607
rect 9597 4573 9631 4607
rect 16865 4573 16899 4607
rect 19073 4573 19107 4607
rect 1409 4505 1443 4539
rect 10885 4505 10919 4539
rect 16037 4505 16071 4539
rect 25605 4505 25639 4539
rect 10057 4437 10091 4471
rect 10425 4437 10459 4471
rect 12357 4437 12391 4471
rect 15577 4437 15611 4471
rect 15945 4437 15979 4471
rect 25881 4437 25915 4471
rect 6469 4233 6503 4267
rect 9505 4233 9539 4267
rect 10885 4233 10919 4267
rect 11529 4233 11563 4267
rect 13645 4233 13679 4267
rect 9689 4165 9723 4199
rect 10977 4165 11011 4199
rect 13185 4165 13219 4199
rect 15761 4165 15795 4199
rect 17049 4165 17083 4199
rect 7113 4097 7147 4131
rect 7481 4097 7515 4131
rect 10057 4097 10091 4131
rect 10333 4097 10367 4131
rect 11713 4097 11747 4131
rect 11989 4097 12023 4131
rect 13737 4097 13771 4131
rect 15209 4097 15243 4131
rect 15853 4097 15887 4131
rect 17141 4097 17175 4131
rect 17785 4097 17819 4131
rect 17877 4097 17911 4131
rect 23581 4097 23615 4131
rect 7665 4029 7699 4063
rect 7941 4029 7975 4063
rect 10701 4029 10735 4063
rect 12357 4029 12391 4063
rect 13829 4029 13863 4063
rect 16037 4029 16071 4063
rect 17233 4029 17267 4063
rect 17601 4029 17635 4063
rect 21833 4029 21867 4063
rect 23305 4029 23339 4063
rect 9413 3961 9447 3995
rect 11345 3961 11379 3995
rect 15393 3961 15427 3995
rect 9689 3893 9723 3927
rect 10149 3893 10183 3927
rect 11805 3893 11839 3927
rect 13277 3893 13311 3927
rect 15025 3893 15059 3927
rect 16681 3893 16715 3927
rect 18245 3893 18279 3927
rect 7389 3689 7423 3723
rect 8309 3689 8343 3723
rect 10504 3689 10538 3723
rect 11989 3689 12023 3723
rect 13829 3689 13863 3723
rect 16221 3689 16255 3723
rect 18061 3689 18095 3723
rect 22477 3689 22511 3723
rect 5641 3553 5675 3587
rect 7941 3553 7975 3587
rect 8125 3553 8159 3587
rect 9505 3553 9539 3587
rect 10241 3553 10275 3587
rect 12081 3553 12115 3587
rect 16313 3553 16347 3587
rect 19717 3553 19751 3587
rect 21465 3553 21499 3587
rect 21833 3553 21867 3587
rect 7849 3485 7883 3519
rect 8493 3485 8527 3519
rect 9321 3485 9355 3519
rect 14197 3485 14231 3519
rect 14473 3485 14507 3519
rect 18153 3485 18187 3519
rect 5917 3417 5951 3451
rect 12357 3417 12391 3451
rect 14749 3417 14783 3451
rect 16589 3417 16623 3451
rect 19993 3417 20027 3451
rect 7481 3349 7515 3383
rect 8953 3349 8987 3383
rect 9413 3349 9447 3383
rect 14381 3349 14415 3383
rect 18337 3349 18371 3383
rect 6561 3145 6595 3179
rect 8401 3145 8435 3179
rect 12265 3145 12299 3179
rect 12541 3145 12575 3179
rect 16129 3145 16163 3179
rect 16497 3145 16531 3179
rect 17141 3145 17175 3179
rect 9873 3077 9907 3111
rect 11805 3077 11839 3111
rect 11897 3077 11931 3111
rect 14657 3077 14691 3111
rect 18613 3077 18647 3111
rect 6745 3009 6779 3043
rect 10149 3009 10183 3043
rect 12725 3009 12759 3043
rect 14381 3009 14415 3043
rect 16313 3009 16347 3043
rect 11713 2941 11747 2975
rect 18889 2941 18923 2975
rect 20085 2601 20119 2635
rect 25789 2601 25823 2635
rect 1777 2397 1811 2431
rect 4353 2397 4387 2431
rect 7941 2397 7975 2431
rect 12081 2397 12115 2431
rect 15945 2397 15979 2431
rect 20269 2397 20303 2431
rect 25973 2397 26007 2431
rect 1409 2329 1443 2363
rect 3985 2329 4019 2363
rect 11713 2329 11747 2363
rect 15577 2329 15611 2363
rect 24501 2329 24535 2363
rect 8033 2261 8067 2295
rect 24593 2261 24627 2295
<< metal1 >>
rect 1104 27226 26472 27248
rect 1104 27174 7252 27226
rect 7304 27174 7316 27226
rect 7368 27174 7380 27226
rect 7432 27174 7444 27226
rect 7496 27174 7508 27226
rect 7560 27174 13554 27226
rect 13606 27174 13618 27226
rect 13670 27174 13682 27226
rect 13734 27174 13746 27226
rect 13798 27174 13810 27226
rect 13862 27174 19856 27226
rect 19908 27174 19920 27226
rect 19972 27174 19984 27226
rect 20036 27174 20048 27226
rect 20100 27174 20112 27226
rect 20164 27174 26158 27226
rect 26210 27174 26222 27226
rect 26274 27174 26286 27226
rect 26338 27174 26350 27226
rect 26402 27174 26414 27226
rect 26466 27174 26472 27226
rect 1104 27152 26472 27174
rect 1673 27115 1731 27121
rect 1673 27081 1685 27115
rect 1719 27112 1731 27115
rect 2774 27112 2780 27124
rect 1719 27084 2780 27112
rect 1719 27081 1731 27084
rect 1673 27075 1731 27081
rect 2774 27072 2780 27084
rect 2832 27072 2838 27124
rect 3234 27072 3240 27124
rect 3292 27112 3298 27124
rect 3881 27115 3939 27121
rect 3881 27112 3893 27115
rect 3292 27084 3893 27112
rect 3292 27072 3298 27084
rect 3881 27081 3893 27084
rect 3927 27081 3939 27115
rect 3881 27075 3939 27081
rect 7098 27072 7104 27124
rect 7156 27072 7162 27124
rect 11606 27072 11612 27124
rect 11664 27072 11670 27124
rect 15194 27112 15200 27124
rect 12406 27084 15200 27112
rect 1762 26936 1768 26988
rect 1820 26936 1826 26988
rect 4157 26979 4215 26985
rect 4157 26945 4169 26979
rect 4203 26976 4215 26979
rect 5074 26976 5080 26988
rect 4203 26948 5080 26976
rect 4203 26945 4215 26948
rect 4157 26939 4215 26945
rect 5074 26936 5080 26948
rect 5132 26936 5138 26988
rect 7116 26976 7144 27072
rect 11057 27047 11115 27053
rect 11057 27013 11069 27047
rect 11103 27044 11115 27047
rect 11103 27016 11376 27044
rect 11103 27013 11115 27016
rect 11057 27007 11115 27013
rect 11348 26988 11376 27016
rect 7377 26979 7435 26985
rect 7377 26976 7389 26979
rect 7116 26948 7389 26976
rect 7377 26945 7389 26948
rect 7423 26945 7435 26979
rect 7377 26939 7435 26945
rect 10781 26979 10839 26985
rect 10781 26945 10793 26979
rect 10827 26976 10839 26979
rect 10827 26948 10861 26976
rect 10827 26945 10839 26948
rect 10781 26939 10839 26945
rect 10597 26911 10655 26917
rect 10597 26877 10609 26911
rect 10643 26908 10655 26911
rect 10796 26908 10824 26939
rect 10962 26936 10968 26988
rect 11020 26936 11026 26988
rect 11149 26979 11207 26985
rect 11149 26945 11161 26979
rect 11195 26945 11207 26979
rect 11149 26939 11207 26945
rect 10643 26880 10824 26908
rect 11164 26908 11192 26939
rect 11330 26936 11336 26988
rect 11388 26936 11394 26988
rect 11624 26976 11652 27072
rect 11701 26979 11759 26985
rect 11701 26976 11713 26979
rect 11624 26948 11713 26976
rect 11701 26945 11713 26948
rect 11747 26945 11759 26979
rect 12406 26976 12434 27084
rect 15194 27072 15200 27084
rect 15252 27072 15258 27124
rect 15746 27072 15752 27124
rect 15804 27072 15810 27124
rect 19334 27072 19340 27124
rect 19392 27072 19398 27124
rect 23474 27072 23480 27124
rect 23532 27072 23538 27124
rect 13173 27047 13231 27053
rect 13173 27013 13185 27047
rect 13219 27044 13231 27047
rect 13446 27044 13452 27056
rect 13219 27016 13452 27044
rect 13219 27013 13231 27016
rect 13173 27007 13231 27013
rect 13446 27004 13452 27016
rect 13504 27004 13510 27056
rect 11701 26939 11759 26945
rect 11808 26948 12434 26976
rect 13081 26979 13139 26985
rect 11808 26908 11836 26948
rect 13081 26945 13093 26979
rect 13127 26976 13139 26979
rect 13998 26976 14004 26988
rect 13127 26948 14004 26976
rect 13127 26945 13139 26948
rect 13081 26939 13139 26945
rect 13998 26936 14004 26948
rect 14056 26936 14062 26988
rect 15654 26936 15660 26988
rect 15712 26936 15718 26988
rect 16761 26979 16819 26985
rect 16761 26945 16773 26979
rect 16807 26976 16819 26979
rect 17126 26976 17132 26988
rect 16807 26948 17132 26976
rect 16807 26945 16819 26948
rect 16761 26939 16819 26945
rect 17126 26936 17132 26948
rect 17184 26936 17190 26988
rect 19352 26976 19380 27072
rect 19429 26979 19487 26985
rect 19429 26976 19441 26979
rect 19352 26948 19441 26976
rect 19429 26945 19441 26948
rect 19475 26945 19487 26979
rect 20990 26976 20996 26988
rect 19429 26939 19487 26945
rect 19536 26948 20996 26976
rect 11164 26880 11836 26908
rect 13357 26911 13415 26917
rect 10643 26877 10655 26880
rect 10597 26871 10655 26877
rect 10796 26784 10824 26880
rect 13357 26877 13369 26911
rect 13403 26908 13415 26911
rect 14918 26908 14924 26920
rect 13403 26880 14924 26908
rect 13403 26877 13415 26880
rect 13357 26871 13415 26877
rect 14918 26868 14924 26880
rect 14976 26868 14982 26920
rect 15378 26868 15384 26920
rect 15436 26908 15442 26920
rect 19536 26908 19564 26948
rect 20990 26936 20996 26948
rect 21048 26936 21054 26988
rect 23492 26985 23520 27072
rect 23477 26979 23535 26985
rect 23477 26945 23489 26979
rect 23523 26945 23535 26979
rect 23477 26939 23535 26945
rect 15436 26880 19564 26908
rect 15436 26868 15442 26880
rect 20714 26868 20720 26920
rect 20772 26868 20778 26920
rect 7190 26732 7196 26784
rect 7248 26732 7254 26784
rect 9766 26732 9772 26784
rect 9824 26772 9830 26784
rect 9953 26775 10011 26781
rect 9953 26772 9965 26775
rect 9824 26744 9965 26772
rect 9824 26732 9830 26744
rect 9953 26741 9965 26744
rect 9999 26741 10011 26775
rect 9953 26735 10011 26741
rect 10778 26732 10784 26784
rect 10836 26732 10842 26784
rect 11333 26775 11391 26781
rect 11333 26741 11345 26775
rect 11379 26772 11391 26775
rect 11422 26772 11428 26784
rect 11379 26744 11428 26772
rect 11379 26741 11391 26744
rect 11333 26735 11391 26741
rect 11422 26732 11428 26744
rect 11480 26732 11486 26784
rect 11885 26775 11943 26781
rect 11885 26741 11897 26775
rect 11931 26772 11943 26775
rect 12250 26772 12256 26784
rect 11931 26744 12256 26772
rect 11931 26741 11943 26744
rect 11885 26735 11943 26741
rect 12250 26732 12256 26744
rect 12308 26732 12314 26784
rect 12434 26732 12440 26784
rect 12492 26772 12498 26784
rect 12713 26775 12771 26781
rect 12713 26772 12725 26775
rect 12492 26744 12725 26772
rect 12492 26732 12498 26744
rect 12713 26741 12725 26744
rect 12759 26741 12771 26775
rect 12713 26735 12771 26741
rect 16945 26775 17003 26781
rect 16945 26741 16957 26775
rect 16991 26772 17003 26775
rect 17034 26772 17040 26784
rect 16991 26744 17040 26772
rect 16991 26741 17003 26744
rect 16945 26735 17003 26741
rect 17034 26732 17040 26744
rect 17092 26732 17098 26784
rect 19610 26732 19616 26784
rect 19668 26732 19674 26784
rect 22462 26732 22468 26784
rect 22520 26772 22526 26784
rect 23293 26775 23351 26781
rect 23293 26772 23305 26775
rect 22520 26744 23305 26772
rect 22520 26732 22526 26744
rect 23293 26741 23305 26744
rect 23339 26741 23351 26775
rect 23293 26735 23351 26741
rect 1104 26682 26312 26704
rect 1104 26630 4101 26682
rect 4153 26630 4165 26682
rect 4217 26630 4229 26682
rect 4281 26630 4293 26682
rect 4345 26630 4357 26682
rect 4409 26630 10403 26682
rect 10455 26630 10467 26682
rect 10519 26630 10531 26682
rect 10583 26630 10595 26682
rect 10647 26630 10659 26682
rect 10711 26630 16705 26682
rect 16757 26630 16769 26682
rect 16821 26630 16833 26682
rect 16885 26630 16897 26682
rect 16949 26630 16961 26682
rect 17013 26630 23007 26682
rect 23059 26630 23071 26682
rect 23123 26630 23135 26682
rect 23187 26630 23199 26682
rect 23251 26630 23263 26682
rect 23315 26630 26312 26682
rect 1104 26608 26312 26630
rect 7190 26528 7196 26580
rect 7248 26528 7254 26580
rect 10689 26571 10747 26577
rect 10689 26537 10701 26571
rect 10735 26568 10747 26571
rect 10778 26568 10784 26580
rect 10735 26540 10784 26568
rect 10735 26537 10747 26540
rect 10689 26531 10747 26537
rect 10778 26528 10784 26540
rect 10836 26528 10842 26580
rect 14918 26528 14924 26580
rect 14976 26568 14982 26580
rect 20796 26571 20854 26577
rect 14976 26540 16068 26568
rect 14976 26528 14982 26540
rect 5905 26435 5963 26441
rect 5905 26401 5917 26435
rect 5951 26432 5963 26435
rect 7208 26432 7236 26528
rect 12897 26503 12955 26509
rect 12897 26469 12909 26503
rect 12943 26469 12955 26503
rect 15286 26500 15292 26512
rect 12897 26463 12955 26469
rect 13556 26472 15292 26500
rect 5951 26404 7236 26432
rect 7377 26435 7435 26441
rect 5951 26401 5963 26404
rect 5905 26395 5963 26401
rect 7377 26401 7389 26435
rect 7423 26432 7435 26435
rect 7469 26435 7527 26441
rect 7469 26432 7481 26435
rect 7423 26404 7481 26432
rect 7423 26401 7435 26404
rect 7377 26395 7435 26401
rect 7469 26401 7481 26404
rect 7515 26401 7527 26435
rect 7469 26395 7527 26401
rect 5629 26367 5687 26373
rect 5629 26333 5641 26367
rect 5675 26333 5687 26367
rect 5629 26327 5687 26333
rect 5644 26296 5672 26327
rect 8478 26324 8484 26376
rect 8536 26364 8542 26376
rect 8941 26367 8999 26373
rect 8941 26364 8953 26367
rect 8536 26336 8953 26364
rect 8536 26324 8542 26336
rect 8941 26333 8953 26336
rect 8987 26333 8999 26367
rect 8941 26327 8999 26333
rect 11330 26324 11336 26376
rect 11388 26324 11394 26376
rect 11790 26324 11796 26376
rect 11848 26364 11854 26376
rect 12437 26367 12495 26373
rect 12437 26364 12449 26367
rect 11848 26336 12449 26364
rect 11848 26324 11854 26336
rect 12437 26333 12449 26336
rect 12483 26333 12495 26367
rect 12437 26327 12495 26333
rect 12805 26367 12863 26373
rect 12805 26333 12817 26367
rect 12851 26364 12863 26367
rect 12912 26364 12940 26463
rect 13556 26441 13584 26472
rect 15286 26460 15292 26472
rect 15344 26460 15350 26512
rect 15381 26503 15439 26509
rect 15381 26469 15393 26503
rect 15427 26500 15439 26503
rect 15470 26500 15476 26512
rect 15427 26472 15476 26500
rect 15427 26469 15439 26472
rect 15381 26463 15439 26469
rect 15470 26460 15476 26472
rect 15528 26460 15534 26512
rect 15933 26503 15991 26509
rect 15933 26469 15945 26503
rect 15979 26469 15991 26503
rect 15933 26463 15991 26469
rect 13541 26435 13599 26441
rect 13541 26401 13553 26435
rect 13587 26401 13599 26435
rect 14550 26432 14556 26444
rect 13541 26395 13599 26401
rect 13832 26404 14556 26432
rect 13832 26364 13860 26404
rect 14550 26392 14556 26404
rect 14608 26392 14614 26444
rect 14660 26404 15148 26432
rect 12851 26336 12940 26364
rect 13280 26336 13860 26364
rect 12851 26333 12863 26336
rect 12805 26327 12863 26333
rect 7650 26296 7656 26308
rect 5460 26268 5672 26296
rect 7130 26268 7656 26296
rect 4982 26188 4988 26240
rect 5040 26228 5046 26240
rect 5460 26228 5488 26268
rect 7650 26256 7656 26268
rect 7708 26256 7714 26308
rect 8846 26256 8852 26308
rect 8904 26296 8910 26308
rect 9217 26299 9275 26305
rect 9217 26296 9229 26299
rect 8904 26268 9229 26296
rect 8904 26256 8910 26268
rect 9217 26265 9229 26268
rect 9263 26265 9275 26299
rect 13280 26296 13308 26336
rect 13906 26324 13912 26376
rect 13964 26364 13970 26376
rect 14660 26373 14688 26404
rect 15120 26373 15148 26404
rect 14645 26367 14703 26373
rect 14645 26364 14657 26367
rect 13964 26336 14657 26364
rect 13964 26324 13970 26336
rect 14645 26333 14657 26336
rect 14691 26333 14703 26367
rect 14645 26327 14703 26333
rect 14829 26367 14887 26373
rect 14829 26333 14841 26367
rect 14875 26333 14887 26367
rect 14829 26327 14887 26333
rect 15105 26367 15163 26373
rect 15105 26333 15117 26367
rect 15151 26333 15163 26367
rect 15105 26327 15163 26333
rect 9217 26259 9275 26265
rect 9600 26268 9706 26296
rect 10442 26268 13308 26296
rect 13357 26299 13415 26305
rect 5040 26200 5488 26228
rect 5040 26188 5046 26200
rect 8018 26188 8024 26240
rect 8076 26228 8082 26240
rect 8113 26231 8171 26237
rect 8113 26228 8125 26231
rect 8076 26200 8125 26228
rect 8076 26188 8082 26200
rect 8113 26197 8125 26200
rect 8159 26197 8171 26231
rect 8113 26191 8171 26197
rect 8202 26188 8208 26240
rect 8260 26228 8266 26240
rect 9600 26228 9628 26268
rect 13357 26265 13369 26299
rect 13403 26296 13415 26299
rect 14093 26299 14151 26305
rect 14093 26296 14105 26299
rect 13403 26268 14105 26296
rect 13403 26265 13415 26268
rect 13357 26259 13415 26265
rect 14093 26265 14105 26268
rect 14139 26265 14151 26299
rect 14844 26296 14872 26327
rect 15194 26324 15200 26376
rect 15252 26324 15258 26376
rect 15749 26367 15807 26373
rect 15749 26333 15761 26367
rect 15795 26364 15807 26367
rect 15948 26364 15976 26463
rect 16040 26432 16068 26540
rect 20796 26537 20808 26571
rect 20842 26568 20854 26571
rect 20842 26540 22094 26568
rect 20842 26537 20854 26540
rect 20796 26531 20854 26537
rect 16485 26435 16543 26441
rect 16485 26432 16497 26435
rect 16040 26404 16497 26432
rect 16485 26401 16497 26404
rect 16531 26401 16543 26435
rect 16485 26395 16543 26401
rect 17405 26435 17463 26441
rect 17405 26401 17417 26435
rect 17451 26432 17463 26435
rect 20533 26435 20591 26441
rect 17451 26404 17724 26432
rect 17451 26401 17463 26404
rect 17405 26395 17463 26401
rect 17696 26376 17724 26404
rect 20533 26401 20545 26435
rect 20579 26432 20591 26435
rect 20898 26432 20904 26444
rect 20579 26404 20904 26432
rect 20579 26401 20591 26404
rect 20533 26395 20591 26401
rect 20898 26392 20904 26404
rect 20956 26392 20962 26444
rect 15795 26336 15976 26364
rect 16393 26367 16451 26373
rect 15795 26333 15807 26336
rect 15749 26327 15807 26333
rect 16393 26333 16405 26367
rect 16439 26364 16451 26367
rect 17310 26364 17316 26376
rect 16439 26336 17316 26364
rect 16439 26333 16451 26336
rect 16393 26327 16451 26333
rect 17310 26324 17316 26336
rect 17368 26324 17374 26376
rect 17494 26324 17500 26376
rect 17552 26324 17558 26376
rect 17678 26324 17684 26376
rect 17736 26324 17742 26376
rect 18414 26324 18420 26376
rect 18472 26364 18478 26376
rect 18785 26367 18843 26373
rect 18785 26364 18797 26367
rect 18472 26336 18797 26364
rect 18472 26324 18478 26336
rect 18785 26333 18797 26336
rect 18831 26333 18843 26367
rect 22066 26364 22094 26540
rect 22281 26435 22339 26441
rect 22281 26401 22293 26435
rect 22327 26432 22339 26435
rect 22830 26432 22836 26444
rect 22327 26404 22836 26432
rect 22327 26401 22339 26404
rect 22281 26395 22339 26401
rect 22830 26392 22836 26404
rect 22888 26392 22894 26444
rect 22465 26367 22523 26373
rect 22465 26364 22477 26367
rect 18785 26327 18843 26333
rect 14093 26259 14151 26265
rect 14568 26268 14872 26296
rect 15013 26299 15071 26305
rect 14568 26240 14596 26268
rect 15013 26265 15025 26299
rect 15059 26265 15071 26299
rect 15013 26259 15071 26265
rect 16301 26299 16359 26305
rect 16301 26265 16313 26299
rect 16347 26296 16359 26299
rect 16761 26299 16819 26305
rect 16761 26296 16773 26299
rect 16347 26268 16773 26296
rect 16347 26265 16359 26268
rect 16301 26259 16359 26265
rect 16761 26265 16773 26268
rect 16807 26265 16819 26299
rect 16761 26259 16819 26265
rect 18141 26299 18199 26305
rect 18141 26265 18153 26299
rect 18187 26296 18199 26299
rect 18506 26296 18512 26308
rect 18187 26268 18512 26296
rect 18187 26265 18199 26268
rect 18141 26259 18199 26265
rect 8260 26200 9628 26228
rect 8260 26188 8266 26200
rect 9950 26188 9956 26240
rect 10008 26228 10014 26240
rect 10781 26231 10839 26237
rect 10781 26228 10793 26231
rect 10008 26200 10793 26228
rect 10008 26188 10014 26200
rect 10781 26197 10793 26200
rect 10827 26197 10839 26231
rect 10781 26191 10839 26197
rect 11882 26188 11888 26240
rect 11940 26188 11946 26240
rect 12526 26188 12532 26240
rect 12584 26228 12590 26240
rect 12621 26231 12679 26237
rect 12621 26228 12633 26231
rect 12584 26200 12633 26228
rect 12584 26188 12590 26200
rect 12621 26197 12633 26200
rect 12667 26197 12679 26231
rect 12621 26191 12679 26197
rect 13265 26231 13323 26237
rect 13265 26197 13277 26231
rect 13311 26228 13323 26231
rect 13446 26228 13452 26240
rect 13311 26200 13452 26228
rect 13311 26197 13323 26200
rect 13265 26191 13323 26197
rect 13446 26188 13452 26200
rect 13504 26188 13510 26240
rect 14550 26188 14556 26240
rect 14608 26188 14614 26240
rect 14826 26188 14832 26240
rect 14884 26228 14890 26240
rect 15028 26228 15056 26259
rect 18506 26256 18512 26268
rect 18564 26256 18570 26308
rect 14884 26200 15056 26228
rect 14884 26188 14890 26200
rect 15562 26188 15568 26240
rect 15620 26188 15626 26240
rect 17402 26188 17408 26240
rect 17460 26228 17466 26240
rect 18233 26231 18291 26237
rect 18233 26228 18245 26231
rect 17460 26200 18245 26228
rect 17460 26188 17466 26200
rect 18233 26197 18245 26200
rect 18279 26197 18291 26231
rect 21928 26228 21956 26350
rect 22066 26336 22477 26364
rect 22465 26333 22477 26336
rect 22511 26333 22523 26367
rect 22465 26327 22523 26333
rect 23017 26367 23075 26373
rect 23017 26333 23029 26367
rect 23063 26333 23075 26367
rect 23017 26327 23075 26333
rect 22094 26256 22100 26308
rect 22152 26296 22158 26308
rect 23032 26296 23060 26327
rect 22152 26268 23060 26296
rect 22152 26256 22158 26268
rect 22738 26228 22744 26240
rect 21928 26200 22744 26228
rect 18233 26191 18291 26197
rect 22738 26188 22744 26200
rect 22796 26188 22802 26240
rect 1104 26138 26472 26160
rect 1104 26086 7252 26138
rect 7304 26086 7316 26138
rect 7368 26086 7380 26138
rect 7432 26086 7444 26138
rect 7496 26086 7508 26138
rect 7560 26086 13554 26138
rect 13606 26086 13618 26138
rect 13670 26086 13682 26138
rect 13734 26086 13746 26138
rect 13798 26086 13810 26138
rect 13862 26086 19856 26138
rect 19908 26086 19920 26138
rect 19972 26086 19984 26138
rect 20036 26086 20048 26138
rect 20100 26086 20112 26138
rect 20164 26086 26158 26138
rect 26210 26086 26222 26138
rect 26274 26086 26286 26138
rect 26338 26086 26350 26138
rect 26402 26086 26414 26138
rect 26466 26086 26472 26138
rect 1104 26064 26472 26086
rect 10229 26027 10287 26033
rect 10229 25993 10241 26027
rect 10275 26024 10287 26027
rect 11330 26024 11336 26036
rect 10275 25996 11336 26024
rect 10275 25993 10287 25996
rect 10229 25987 10287 25993
rect 11330 25984 11336 25996
rect 11388 25984 11394 26036
rect 11440 25996 12756 26024
rect 7466 25916 7472 25968
rect 7524 25916 7530 25968
rect 7929 25959 7987 25965
rect 7929 25925 7941 25959
rect 7975 25956 7987 25959
rect 8018 25956 8024 25968
rect 7975 25928 8024 25956
rect 7975 25925 7987 25928
rect 7929 25919 7987 25925
rect 8018 25916 8024 25928
rect 8076 25916 8082 25968
rect 11440 25956 11468 25996
rect 12342 25956 12348 25968
rect 10336 25928 11468 25956
rect 11900 25928 12348 25956
rect 10336 25888 10364 25928
rect 9890 25860 10364 25888
rect 10413 25891 10471 25897
rect 10413 25857 10425 25891
rect 10459 25857 10471 25891
rect 10413 25851 10471 25857
rect 5902 25780 5908 25832
rect 5960 25820 5966 25832
rect 6089 25823 6147 25829
rect 6089 25820 6101 25823
rect 5960 25792 6101 25820
rect 5960 25780 5966 25792
rect 6089 25789 6101 25792
rect 6135 25820 6147 25823
rect 6457 25823 6515 25829
rect 6457 25820 6469 25823
rect 6135 25792 6469 25820
rect 6135 25789 6147 25792
rect 6089 25783 6147 25789
rect 6457 25789 6469 25792
rect 6503 25789 6515 25823
rect 6457 25783 6515 25789
rect 6914 25780 6920 25832
rect 6972 25820 6978 25832
rect 8205 25823 8263 25829
rect 8205 25820 8217 25823
rect 6972 25792 8217 25820
rect 6972 25780 6978 25792
rect 8205 25789 8217 25792
rect 8251 25820 8263 25823
rect 8478 25820 8484 25832
rect 8251 25792 8484 25820
rect 8251 25789 8263 25792
rect 8205 25783 8263 25789
rect 8478 25780 8484 25792
rect 8536 25780 8542 25832
rect 8754 25780 8760 25832
rect 8812 25780 8818 25832
rect 10428 25752 10456 25851
rect 10888 25832 10916 25928
rect 11330 25848 11336 25900
rect 11388 25848 11394 25900
rect 11900 25897 11928 25928
rect 12342 25916 12348 25928
rect 12400 25916 12406 25968
rect 12437 25959 12495 25965
rect 12437 25925 12449 25959
rect 12483 25956 12495 25959
rect 12526 25956 12532 25968
rect 12483 25928 12532 25956
rect 12483 25925 12495 25928
rect 12437 25919 12495 25925
rect 12526 25916 12532 25928
rect 12584 25916 12590 25968
rect 12728 25956 12756 25996
rect 13906 25984 13912 26036
rect 13964 25984 13970 26036
rect 13998 25984 14004 26036
rect 14056 25984 14062 26036
rect 15378 25984 15384 26036
rect 15436 25984 15442 26036
rect 18248 25996 18920 26024
rect 12728 25928 12926 25956
rect 14642 25916 14648 25968
rect 14700 25956 14706 25968
rect 15396 25956 15424 25984
rect 18248 25968 18276 25996
rect 16945 25959 17003 25965
rect 14700 25928 15502 25956
rect 14700 25916 14706 25928
rect 16945 25925 16957 25959
rect 16991 25956 17003 25959
rect 17034 25956 17040 25968
rect 16991 25928 17040 25956
rect 16991 25925 17003 25928
rect 16945 25919 17003 25925
rect 17034 25916 17040 25928
rect 17092 25916 17098 25968
rect 18230 25956 18236 25968
rect 18170 25928 18236 25956
rect 18230 25916 18236 25928
rect 18288 25916 18294 25968
rect 18506 25916 18512 25968
rect 18564 25956 18570 25968
rect 18785 25959 18843 25965
rect 18785 25956 18797 25959
rect 18564 25928 18797 25956
rect 18564 25916 18570 25928
rect 18785 25925 18797 25928
rect 18831 25925 18843 25959
rect 18892 25956 18920 25996
rect 22189 25959 22247 25965
rect 18892 25928 19274 25956
rect 18785 25919 18843 25925
rect 22189 25925 22201 25959
rect 22235 25956 22247 25959
rect 22462 25956 22468 25968
rect 22235 25928 22468 25956
rect 22235 25925 22247 25928
rect 22189 25919 22247 25925
rect 22462 25916 22468 25928
rect 22520 25916 22526 25968
rect 22738 25916 22744 25968
rect 22796 25916 22802 25968
rect 11885 25891 11943 25897
rect 11885 25857 11897 25891
rect 11931 25857 11943 25891
rect 11885 25851 11943 25857
rect 14458 25848 14464 25900
rect 14516 25888 14522 25900
rect 14737 25891 14795 25897
rect 14737 25888 14749 25891
rect 14516 25860 14749 25888
rect 14516 25848 14522 25860
rect 14737 25857 14749 25860
rect 14783 25857 14795 25891
rect 14737 25851 14795 25857
rect 20806 25848 20812 25900
rect 20864 25888 20870 25900
rect 21269 25891 21327 25897
rect 21269 25888 21281 25891
rect 20864 25860 21281 25888
rect 20864 25848 20870 25860
rect 21269 25857 21281 25860
rect 21315 25857 21327 25891
rect 21269 25851 21327 25857
rect 10870 25780 10876 25832
rect 10928 25780 10934 25832
rect 11974 25780 11980 25832
rect 12032 25820 12038 25832
rect 12161 25823 12219 25829
rect 12161 25820 12173 25823
rect 12032 25792 12173 25820
rect 12032 25780 12038 25792
rect 12161 25789 12173 25792
rect 12207 25820 12219 25823
rect 14476 25820 14504 25848
rect 12207 25792 14504 25820
rect 12207 25789 12219 25792
rect 12161 25783 12219 25789
rect 14550 25780 14556 25832
rect 14608 25780 14614 25832
rect 15013 25823 15071 25829
rect 15013 25789 15025 25823
rect 15059 25820 15071 25823
rect 15562 25820 15568 25832
rect 15059 25792 15568 25820
rect 15059 25789 15071 25792
rect 15013 25783 15071 25789
rect 15562 25780 15568 25792
rect 15620 25780 15626 25832
rect 16574 25780 16580 25832
rect 16632 25820 16638 25832
rect 16669 25823 16727 25829
rect 16669 25820 16681 25823
rect 16632 25792 16681 25820
rect 16632 25780 16638 25792
rect 16669 25789 16681 25792
rect 16715 25789 16727 25823
rect 16669 25783 16727 25789
rect 18414 25780 18420 25832
rect 18472 25780 18478 25832
rect 18509 25823 18567 25829
rect 18509 25789 18521 25823
rect 18555 25789 18567 25823
rect 18509 25783 18567 25789
rect 10428 25724 12296 25752
rect 5350 25644 5356 25696
rect 5408 25684 5414 25696
rect 5537 25687 5595 25693
rect 5537 25684 5549 25687
rect 5408 25656 5549 25684
rect 5408 25644 5414 25656
rect 5537 25653 5549 25656
rect 5583 25653 5595 25687
rect 5537 25647 5595 25653
rect 7466 25644 7472 25696
rect 7524 25684 7530 25696
rect 10428 25684 10456 25724
rect 7524 25656 10456 25684
rect 7524 25644 7530 25656
rect 10778 25644 10784 25696
rect 10836 25684 10842 25696
rect 11149 25687 11207 25693
rect 11149 25684 11161 25687
rect 10836 25656 11161 25684
rect 10836 25644 10842 25656
rect 11149 25653 11161 25656
rect 11195 25653 11207 25687
rect 11149 25647 11207 25653
rect 12069 25687 12127 25693
rect 12069 25653 12081 25687
rect 12115 25684 12127 25687
rect 12158 25684 12164 25696
rect 12115 25656 12164 25684
rect 12115 25653 12127 25656
rect 12069 25647 12127 25653
rect 12158 25644 12164 25656
rect 12216 25644 12222 25696
rect 12268 25684 12296 25724
rect 12618 25684 12624 25696
rect 12268 25656 12624 25684
rect 12618 25644 12624 25656
rect 12676 25644 12682 25696
rect 16485 25687 16543 25693
rect 16485 25653 16497 25687
rect 16531 25684 16543 25687
rect 17678 25684 17684 25696
rect 16531 25656 17684 25684
rect 16531 25653 16543 25656
rect 16485 25647 16543 25653
rect 17678 25644 17684 25656
rect 17736 25644 17742 25696
rect 18524 25684 18552 25783
rect 20622 25780 20628 25832
rect 20680 25780 20686 25832
rect 20898 25780 20904 25832
rect 20956 25820 20962 25832
rect 21913 25823 21971 25829
rect 21913 25820 21925 25823
rect 20956 25792 21925 25820
rect 20956 25780 20962 25792
rect 21913 25789 21925 25792
rect 21959 25789 21971 25823
rect 21913 25783 21971 25789
rect 19242 25684 19248 25696
rect 18524 25656 19248 25684
rect 19242 25644 19248 25656
rect 19300 25644 19306 25696
rect 20254 25644 20260 25696
rect 20312 25644 20318 25696
rect 21174 25644 21180 25696
rect 21232 25644 21238 25696
rect 21450 25644 21456 25696
rect 21508 25644 21514 25696
rect 23658 25644 23664 25696
rect 23716 25644 23722 25696
rect 1104 25594 26312 25616
rect 1104 25542 4101 25594
rect 4153 25542 4165 25594
rect 4217 25542 4229 25594
rect 4281 25542 4293 25594
rect 4345 25542 4357 25594
rect 4409 25542 10403 25594
rect 10455 25542 10467 25594
rect 10519 25542 10531 25594
rect 10583 25542 10595 25594
rect 10647 25542 10659 25594
rect 10711 25542 16705 25594
rect 16757 25542 16769 25594
rect 16821 25542 16833 25594
rect 16885 25542 16897 25594
rect 16949 25542 16961 25594
rect 17013 25542 23007 25594
rect 23059 25542 23071 25594
rect 23123 25542 23135 25594
rect 23187 25542 23199 25594
rect 23251 25542 23263 25594
rect 23315 25542 26312 25594
rect 1104 25520 26312 25542
rect 8754 25440 8760 25492
rect 8812 25480 8818 25492
rect 8941 25483 8999 25489
rect 8941 25480 8953 25483
rect 8812 25452 8953 25480
rect 8812 25440 8818 25452
rect 8941 25449 8953 25452
rect 8987 25449 8999 25483
rect 8941 25443 8999 25449
rect 10308 25483 10366 25489
rect 10308 25449 10320 25483
rect 10354 25480 10366 25483
rect 10778 25480 10784 25492
rect 10354 25452 10784 25480
rect 10354 25449 10366 25452
rect 10308 25443 10366 25449
rect 10778 25440 10784 25452
rect 10836 25440 10842 25492
rect 11790 25440 11796 25492
rect 11848 25440 11854 25492
rect 11974 25440 11980 25492
rect 12032 25440 12038 25492
rect 12158 25489 12164 25492
rect 12148 25483 12164 25489
rect 12148 25449 12160 25483
rect 12148 25443 12164 25449
rect 12158 25440 12164 25443
rect 12216 25440 12222 25492
rect 12250 25440 12256 25492
rect 12308 25480 12314 25492
rect 13633 25483 13691 25489
rect 12308 25452 13400 25480
rect 12308 25440 12314 25452
rect 9217 25415 9275 25421
rect 9217 25381 9229 25415
rect 9263 25381 9275 25415
rect 9217 25375 9275 25381
rect 5261 25347 5319 25353
rect 5261 25313 5273 25347
rect 5307 25344 5319 25347
rect 5350 25344 5356 25356
rect 5307 25316 5356 25344
rect 5307 25313 5319 25316
rect 5261 25307 5319 25313
rect 5350 25304 5356 25316
rect 5408 25304 5414 25356
rect 7193 25347 7251 25353
rect 7193 25344 7205 25347
rect 6932 25316 7205 25344
rect 934 25236 940 25288
rect 992 25276 998 25288
rect 1397 25279 1455 25285
rect 1397 25276 1409 25279
rect 992 25248 1409 25276
rect 992 25236 998 25248
rect 1397 25245 1409 25248
rect 1443 25245 1455 25279
rect 1397 25239 1455 25245
rect 4430 25236 4436 25288
rect 4488 25276 4494 25288
rect 4982 25276 4988 25288
rect 4488 25248 4988 25276
rect 4488 25236 4494 25248
rect 4982 25236 4988 25248
rect 5040 25236 5046 25288
rect 6825 25279 6883 25285
rect 6825 25245 6837 25279
rect 6871 25245 6883 25279
rect 6825 25239 6883 25245
rect 6270 25168 6276 25220
rect 6328 25168 6334 25220
rect 6840 25208 6868 25239
rect 6932 25220 6960 25316
rect 7193 25313 7205 25316
rect 7239 25344 7251 25347
rect 8202 25344 8208 25356
rect 7239 25316 8208 25344
rect 7239 25313 7251 25316
rect 7193 25307 7251 25313
rect 8202 25304 8208 25316
rect 8260 25304 8266 25356
rect 8570 25236 8576 25288
rect 8628 25236 8634 25288
rect 8846 25236 8852 25288
rect 8904 25236 8910 25288
rect 9125 25279 9183 25285
rect 9125 25245 9137 25279
rect 9171 25276 9183 25279
rect 9232 25276 9260 25375
rect 9582 25304 9588 25356
rect 9640 25344 9646 25356
rect 9769 25347 9827 25353
rect 9769 25344 9781 25347
rect 9640 25316 9781 25344
rect 9640 25304 9646 25316
rect 9769 25313 9781 25316
rect 9815 25313 9827 25347
rect 9769 25307 9827 25313
rect 9950 25304 9956 25356
rect 10008 25304 10014 25356
rect 10045 25347 10103 25353
rect 10045 25313 10057 25347
rect 10091 25344 10103 25347
rect 11885 25347 11943 25353
rect 11885 25344 11897 25347
rect 10091 25316 11897 25344
rect 10091 25313 10103 25316
rect 10045 25307 10103 25313
rect 11885 25313 11897 25316
rect 11931 25344 11943 25347
rect 11992 25344 12020 25440
rect 13372 25412 13400 25452
rect 13633 25449 13645 25483
rect 13679 25480 13691 25483
rect 14550 25480 14556 25492
rect 13679 25452 14556 25480
rect 13679 25449 13691 25452
rect 13633 25443 13691 25449
rect 14550 25440 14556 25452
rect 14608 25440 14614 25492
rect 15286 25440 15292 25492
rect 15344 25480 15350 25492
rect 16945 25483 17003 25489
rect 15344 25452 16160 25480
rect 15344 25440 15350 25452
rect 13372 25384 14596 25412
rect 11931 25316 12020 25344
rect 11931 25313 11943 25316
rect 11885 25307 11943 25313
rect 14458 25304 14464 25356
rect 14516 25304 14522 25356
rect 14568 25344 14596 25384
rect 14737 25347 14795 25353
rect 14737 25344 14749 25347
rect 14568 25316 14749 25344
rect 14737 25313 14749 25316
rect 14783 25313 14795 25347
rect 14737 25307 14795 25313
rect 15194 25304 15200 25356
rect 15252 25344 15258 25356
rect 16132 25344 16160 25452
rect 16945 25449 16957 25483
rect 16991 25480 17003 25483
rect 17126 25480 17132 25492
rect 16991 25452 17132 25480
rect 16991 25449 17003 25452
rect 16945 25443 17003 25449
rect 17126 25440 17132 25452
rect 17184 25440 17190 25492
rect 17494 25440 17500 25492
rect 17552 25440 17558 25492
rect 20993 25483 21051 25489
rect 20993 25449 21005 25483
rect 21039 25480 21051 25483
rect 22094 25480 22100 25492
rect 21039 25452 22100 25480
rect 21039 25449 21051 25452
rect 20993 25443 21051 25449
rect 22094 25440 22100 25452
rect 22152 25440 22158 25492
rect 23658 25440 23664 25492
rect 23716 25440 23722 25492
rect 25869 25483 25927 25489
rect 25869 25449 25881 25483
rect 25915 25480 25927 25483
rect 25915 25452 26372 25480
rect 25915 25449 25927 25452
rect 25869 25443 25927 25449
rect 16209 25415 16267 25421
rect 16209 25381 16221 25415
rect 16255 25412 16267 25415
rect 17512 25412 17540 25440
rect 16255 25384 17540 25412
rect 17604 25384 18920 25412
rect 16255 25381 16267 25384
rect 16209 25375 16267 25381
rect 16298 25344 16304 25356
rect 15252 25316 15976 25344
rect 16132 25316 16304 25344
rect 15252 25304 15258 25316
rect 9171 25248 9260 25276
rect 9677 25279 9735 25285
rect 9171 25245 9183 25248
rect 9125 25239 9183 25245
rect 9677 25245 9689 25279
rect 9723 25276 9735 25279
rect 9968 25276 9996 25304
rect 9723 25248 9996 25276
rect 15948 25276 15976 25316
rect 16298 25304 16304 25316
rect 16356 25344 16362 25356
rect 17497 25347 17555 25353
rect 17497 25344 17509 25347
rect 16356 25316 17509 25344
rect 16356 25304 16362 25316
rect 17497 25313 17509 25316
rect 17543 25313 17555 25347
rect 17497 25307 17555 25313
rect 15948 25248 17264 25276
rect 9723 25245 9735 25248
rect 9677 25239 9735 25245
rect 6564 25180 6868 25208
rect 1581 25143 1639 25149
rect 1581 25109 1593 25143
rect 1627 25140 1639 25143
rect 6564 25140 6592 25180
rect 6914 25168 6920 25220
rect 6972 25168 6978 25220
rect 1627 25112 6592 25140
rect 6733 25143 6791 25149
rect 1627 25109 1639 25112
rect 1581 25103 1639 25109
rect 6733 25109 6745 25143
rect 6779 25140 6791 25143
rect 7098 25140 7104 25152
rect 6779 25112 7104 25140
rect 6779 25109 6791 25112
rect 6733 25103 6791 25109
rect 7098 25100 7104 25112
rect 7156 25100 7162 25152
rect 8757 25143 8815 25149
rect 8757 25109 8769 25143
rect 8803 25140 8815 25143
rect 8864 25140 8892 25236
rect 10870 25168 10876 25220
rect 10928 25168 10934 25220
rect 12618 25168 12624 25220
rect 12676 25168 12682 25220
rect 17236 25208 17264 25248
rect 17310 25236 17316 25288
rect 17368 25236 17374 25288
rect 17402 25236 17408 25288
rect 17460 25236 17466 25288
rect 17604 25208 17632 25384
rect 17770 25304 17776 25356
rect 17828 25304 17834 25356
rect 18432 25316 18828 25344
rect 18432 25288 18460 25316
rect 18322 25236 18328 25288
rect 18380 25236 18386 25288
rect 18414 25236 18420 25288
rect 18472 25236 18478 25288
rect 18800 25285 18828 25316
rect 18892 25285 18920 25384
rect 19521 25347 19579 25353
rect 19521 25313 19533 25347
rect 19567 25344 19579 25347
rect 19610 25344 19616 25356
rect 19567 25316 19616 25344
rect 19567 25313 19579 25316
rect 19521 25307 19579 25313
rect 19610 25304 19616 25316
rect 19668 25304 19674 25356
rect 20714 25304 20720 25356
rect 20772 25304 20778 25356
rect 20898 25304 20904 25356
rect 20956 25344 20962 25356
rect 21085 25347 21143 25353
rect 21085 25344 21097 25347
rect 20956 25316 21097 25344
rect 20956 25304 20962 25316
rect 21085 25313 21097 25316
rect 21131 25313 21143 25347
rect 21085 25307 21143 25313
rect 21361 25347 21419 25353
rect 21361 25313 21373 25347
rect 21407 25344 21419 25347
rect 21450 25344 21456 25356
rect 21407 25316 21456 25344
rect 21407 25313 21419 25316
rect 21361 25307 21419 25313
rect 21450 25304 21456 25316
rect 21508 25304 21514 25356
rect 22554 25304 22560 25356
rect 22612 25344 22618 25356
rect 22833 25347 22891 25353
rect 22833 25344 22845 25347
rect 22612 25316 22845 25344
rect 22612 25304 22618 25316
rect 22833 25313 22845 25316
rect 22879 25344 22891 25347
rect 23477 25347 23535 25353
rect 23477 25344 23489 25347
rect 22879 25316 23489 25344
rect 22879 25313 22891 25316
rect 22833 25307 22891 25313
rect 23477 25313 23489 25316
rect 23523 25313 23535 25347
rect 23676 25344 23704 25440
rect 26344 25424 26372 25452
rect 26326 25372 26332 25424
rect 26384 25372 26390 25424
rect 24949 25347 25007 25353
rect 24949 25344 24961 25347
rect 23676 25316 24961 25344
rect 23477 25307 23535 25313
rect 24949 25313 24961 25316
rect 24995 25313 25007 25347
rect 24949 25307 25007 25313
rect 18509 25279 18567 25285
rect 18509 25245 18521 25279
rect 18555 25245 18567 25279
rect 18509 25239 18567 25245
rect 18785 25279 18843 25285
rect 18785 25245 18797 25279
rect 18831 25245 18843 25279
rect 18785 25239 18843 25245
rect 18877 25279 18935 25285
rect 18877 25245 18889 25279
rect 18923 25245 18935 25279
rect 18877 25239 18935 25245
rect 15962 25180 16896 25208
rect 17236 25180 17632 25208
rect 8803 25112 8892 25140
rect 8803 25109 8815 25112
rect 8757 25103 8815 25109
rect 9490 25100 9496 25152
rect 9548 25140 9554 25152
rect 9585 25143 9643 25149
rect 9585 25140 9597 25143
rect 9548 25112 9597 25140
rect 9548 25100 9554 25112
rect 9585 25109 9597 25112
rect 9631 25109 9643 25143
rect 9585 25103 9643 25109
rect 15102 25100 15108 25152
rect 15160 25140 15166 25152
rect 16040 25140 16068 25180
rect 15160 25112 16068 25140
rect 16868 25140 16896 25180
rect 17678 25168 17684 25220
rect 17736 25208 17742 25220
rect 18524 25208 18552 25239
rect 19242 25236 19248 25288
rect 19300 25236 19306 25288
rect 17736 25180 18552 25208
rect 18693 25211 18751 25217
rect 17736 25168 17742 25180
rect 18693 25177 18705 25211
rect 18739 25177 18751 25211
rect 20732 25208 20760 25304
rect 25682 25236 25688 25288
rect 25740 25236 25746 25288
rect 20732 25194 21850 25208
rect 20746 25180 21850 25194
rect 18693 25171 18751 25177
rect 18046 25140 18052 25152
rect 16868 25112 18052 25140
rect 15160 25100 15166 25112
rect 18046 25100 18052 25112
rect 18104 25100 18110 25152
rect 18138 25100 18144 25152
rect 18196 25140 18202 25152
rect 18708 25140 18736 25171
rect 21376 25152 21404 25180
rect 22646 25168 22652 25220
rect 22704 25208 22710 25220
rect 22925 25211 22983 25217
rect 22925 25208 22937 25211
rect 22704 25180 22937 25208
rect 22704 25168 22710 25180
rect 22925 25177 22937 25180
rect 22971 25177 22983 25211
rect 22925 25171 22983 25177
rect 18196 25112 18736 25140
rect 18196 25100 18202 25112
rect 18966 25100 18972 25152
rect 19024 25140 19030 25152
rect 19061 25143 19119 25149
rect 19061 25140 19073 25143
rect 19024 25112 19073 25140
rect 19024 25100 19030 25112
rect 19061 25109 19073 25112
rect 19107 25109 19119 25143
rect 19061 25103 19119 25109
rect 21358 25100 21364 25152
rect 21416 25100 21422 25152
rect 24394 25100 24400 25152
rect 24452 25100 24458 25152
rect 1104 25050 26472 25072
rect 1104 24998 7252 25050
rect 7304 24998 7316 25050
rect 7368 24998 7380 25050
rect 7432 24998 7444 25050
rect 7496 24998 7508 25050
rect 7560 24998 13554 25050
rect 13606 24998 13618 25050
rect 13670 24998 13682 25050
rect 13734 24998 13746 25050
rect 13798 24998 13810 25050
rect 13862 24998 19856 25050
rect 19908 24998 19920 25050
rect 19972 24998 19984 25050
rect 20036 24998 20048 25050
rect 20100 24998 20112 25050
rect 20164 24998 26158 25050
rect 26210 24998 26222 25050
rect 26274 24998 26286 25050
rect 26338 24998 26350 25050
rect 26402 24998 26414 25050
rect 26466 24998 26472 25050
rect 1104 24976 26472 24998
rect 8570 24896 8576 24948
rect 8628 24936 8634 24948
rect 8757 24939 8815 24945
rect 8757 24936 8769 24939
rect 8628 24908 8769 24936
rect 8628 24896 8634 24908
rect 8757 24905 8769 24908
rect 8803 24905 8815 24939
rect 8757 24899 8815 24905
rect 9125 24939 9183 24945
rect 9125 24905 9137 24939
rect 9171 24936 9183 24939
rect 9766 24936 9772 24948
rect 9171 24908 9772 24936
rect 9171 24905 9183 24908
rect 9125 24899 9183 24905
rect 9766 24896 9772 24908
rect 9824 24896 9830 24948
rect 11330 24896 11336 24948
rect 11388 24936 11394 24948
rect 11517 24939 11575 24945
rect 11517 24936 11529 24939
rect 11388 24908 11529 24936
rect 11388 24896 11394 24908
rect 11517 24905 11529 24908
rect 11563 24905 11575 24939
rect 11517 24899 11575 24905
rect 11882 24896 11888 24948
rect 11940 24896 11946 24948
rect 13170 24936 13176 24948
rect 13004 24908 13176 24936
rect 5994 24868 6000 24880
rect 5934 24840 6000 24868
rect 5994 24828 6000 24840
rect 6052 24868 6058 24880
rect 6270 24868 6276 24880
rect 6052 24840 6276 24868
rect 6052 24828 6058 24840
rect 6270 24828 6276 24840
rect 6328 24868 6334 24880
rect 7009 24871 7067 24877
rect 7009 24868 7021 24871
rect 6328 24840 7021 24868
rect 6328 24828 6334 24840
rect 7009 24837 7021 24840
rect 7055 24868 7067 24871
rect 7650 24868 7656 24880
rect 7055 24840 7656 24868
rect 7055 24837 7067 24840
rect 7009 24831 7067 24837
rect 7650 24828 7656 24840
rect 7708 24828 7714 24880
rect 8496 24840 9628 24868
rect 8496 24812 8524 24840
rect 6454 24760 6460 24812
rect 6512 24800 6518 24812
rect 6914 24800 6920 24812
rect 6512 24772 6920 24800
rect 6512 24760 6518 24772
rect 6914 24760 6920 24772
rect 6972 24760 6978 24812
rect 7098 24760 7104 24812
rect 7156 24760 7162 24812
rect 7190 24760 7196 24812
rect 7248 24760 7254 24812
rect 8478 24760 8484 24812
rect 8536 24760 8542 24812
rect 9600 24809 9628 24840
rect 9217 24803 9275 24809
rect 9217 24769 9229 24803
rect 9263 24800 9275 24803
rect 9585 24803 9643 24809
rect 9263 24772 9536 24800
rect 9263 24769 9275 24772
rect 9217 24763 9275 24769
rect 4430 24692 4436 24744
rect 4488 24692 4494 24744
rect 4706 24692 4712 24744
rect 4764 24692 4770 24744
rect 7116 24732 7144 24760
rect 9508 24744 9536 24772
rect 9585 24769 9597 24803
rect 9631 24769 9643 24803
rect 9585 24763 9643 24769
rect 10870 24760 10876 24812
rect 10928 24800 10934 24812
rect 13004 24809 13032 24908
rect 13170 24896 13176 24908
rect 13228 24936 13234 24948
rect 14274 24936 14280 24948
rect 13228 24908 14280 24936
rect 13228 24896 13234 24908
rect 14274 24896 14280 24908
rect 14332 24896 14338 24948
rect 16776 24908 18552 24936
rect 15933 24871 15991 24877
rect 15933 24868 15945 24871
rect 15396 24840 15945 24868
rect 12989 24803 13047 24809
rect 10928 24772 10994 24800
rect 10928 24760 10934 24772
rect 12989 24769 13001 24803
rect 13035 24769 13047 24803
rect 14550 24800 14556 24812
rect 14398 24772 14556 24800
rect 12989 24763 13047 24769
rect 14550 24760 14556 24772
rect 14608 24760 14614 24812
rect 7285 24735 7343 24741
rect 7285 24732 7297 24735
rect 7116 24704 7297 24732
rect 7285 24701 7297 24704
rect 7331 24701 7343 24735
rect 7285 24695 7343 24701
rect 9398 24692 9404 24744
rect 9456 24692 9462 24744
rect 9490 24692 9496 24744
rect 9548 24692 9554 24744
rect 9858 24692 9864 24744
rect 9916 24692 9922 24744
rect 11054 24692 11060 24744
rect 11112 24732 11118 24744
rect 11977 24735 12035 24741
rect 11977 24732 11989 24735
rect 11112 24704 11989 24732
rect 11112 24692 11118 24704
rect 11977 24701 11989 24704
rect 12023 24701 12035 24735
rect 11977 24695 12035 24701
rect 12161 24735 12219 24741
rect 12161 24701 12173 24735
rect 12207 24732 12219 24735
rect 12342 24732 12348 24744
rect 12207 24704 12348 24732
rect 12207 24701 12219 24704
rect 12161 24695 12219 24701
rect 12342 24692 12348 24704
rect 12400 24692 12406 24744
rect 13262 24692 13268 24744
rect 13320 24692 13326 24744
rect 13814 24692 13820 24744
rect 13872 24732 13878 24744
rect 14829 24735 14887 24741
rect 14829 24732 14841 24735
rect 13872 24704 14841 24732
rect 13872 24692 13878 24704
rect 14829 24701 14841 24704
rect 14875 24701 14887 24735
rect 14829 24695 14887 24701
rect 14918 24692 14924 24744
rect 14976 24732 14982 24744
rect 15396 24741 15424 24840
rect 15933 24837 15945 24840
rect 15979 24837 15991 24871
rect 15933 24831 15991 24837
rect 15470 24760 15476 24812
rect 15528 24800 15534 24812
rect 15565 24803 15623 24809
rect 15565 24800 15577 24803
rect 15528 24772 15577 24800
rect 15528 24760 15534 24772
rect 15565 24769 15577 24772
rect 15611 24769 15623 24803
rect 15565 24763 15623 24769
rect 15658 24803 15716 24809
rect 15658 24769 15670 24803
rect 15704 24769 15716 24803
rect 15658 24763 15716 24769
rect 15841 24803 15899 24809
rect 15841 24769 15853 24803
rect 15887 24769 15899 24803
rect 15841 24763 15899 24769
rect 15381 24735 15439 24741
rect 15381 24732 15393 24735
rect 14976 24704 15393 24732
rect 14976 24692 14982 24704
rect 15381 24701 15393 24704
rect 15427 24701 15439 24735
rect 15672 24732 15700 24763
rect 15381 24695 15439 24701
rect 15580 24704 15700 24732
rect 15856 24732 15884 24763
rect 16022 24760 16028 24812
rect 16080 24809 16086 24812
rect 16080 24803 16129 24809
rect 16080 24769 16083 24803
rect 16117 24769 16129 24803
rect 16080 24763 16129 24769
rect 16080 24760 16086 24763
rect 16776 24732 16804 24908
rect 17494 24868 17500 24880
rect 16868 24840 17500 24868
rect 16868 24809 16896 24840
rect 17494 24828 17500 24840
rect 17552 24828 17558 24880
rect 18230 24828 18236 24880
rect 18288 24828 18294 24880
rect 16853 24803 16911 24809
rect 16853 24769 16865 24803
rect 16899 24769 16911 24803
rect 18524 24800 18552 24908
rect 20898 24896 20904 24948
rect 20956 24896 20962 24948
rect 20714 24828 20720 24880
rect 20772 24828 20778 24880
rect 20916 24868 20944 24896
rect 23845 24871 23903 24877
rect 20916 24840 21588 24868
rect 18874 24800 18880 24812
rect 18524 24772 18880 24800
rect 16853 24763 16911 24769
rect 18874 24760 18880 24772
rect 18932 24760 18938 24812
rect 21560 24809 21588 24840
rect 23845 24837 23857 24871
rect 23891 24868 23903 24871
rect 24394 24868 24400 24880
rect 23891 24840 24400 24868
rect 23891 24837 23903 24840
rect 23845 24831 23903 24837
rect 24394 24828 24400 24840
rect 24452 24828 24458 24880
rect 21545 24803 21603 24809
rect 21545 24769 21557 24803
rect 21591 24769 21603 24803
rect 21545 24763 21603 24769
rect 15856 24704 16804 24732
rect 16945 24735 17003 24741
rect 7558 24624 7564 24676
rect 7616 24624 7622 24676
rect 14737 24667 14795 24673
rect 14737 24633 14749 24667
rect 14783 24664 14795 24667
rect 15194 24664 15200 24676
rect 14783 24636 15200 24664
rect 14783 24633 14795 24636
rect 14737 24627 14795 24633
rect 15194 24624 15200 24636
rect 15252 24664 15258 24676
rect 15580 24664 15608 24704
rect 15856 24664 15884 24704
rect 16945 24701 16957 24735
rect 16991 24732 17003 24735
rect 17221 24735 17279 24741
rect 16991 24704 17080 24732
rect 16991 24701 17003 24704
rect 16945 24695 17003 24701
rect 15252 24636 15608 24664
rect 15672 24636 15884 24664
rect 15252 24624 15258 24636
rect 6181 24599 6239 24605
rect 6181 24565 6193 24599
rect 6227 24596 6239 24599
rect 7193 24599 7251 24605
rect 7193 24596 7205 24599
rect 6227 24568 7205 24596
rect 6227 24565 6239 24568
rect 6181 24559 6239 24565
rect 7193 24565 7205 24568
rect 7239 24565 7251 24599
rect 7193 24559 7251 24565
rect 11333 24599 11391 24605
rect 11333 24565 11345 24599
rect 11379 24596 11391 24599
rect 11514 24596 11520 24608
rect 11379 24568 11520 24596
rect 11379 24565 11391 24568
rect 11333 24559 11391 24565
rect 11514 24556 11520 24568
rect 11572 24556 11578 24608
rect 13078 24556 13084 24608
rect 13136 24596 13142 24608
rect 15672 24596 15700 24636
rect 13136 24568 15700 24596
rect 13136 24556 13142 24568
rect 15746 24556 15752 24608
rect 15804 24596 15810 24608
rect 16209 24599 16267 24605
rect 16209 24596 16221 24599
rect 15804 24568 16221 24596
rect 15804 24556 15810 24568
rect 16209 24565 16221 24568
rect 16255 24565 16267 24599
rect 16209 24559 16267 24565
rect 16482 24556 16488 24608
rect 16540 24596 16546 24608
rect 16669 24599 16727 24605
rect 16669 24596 16681 24599
rect 16540 24568 16681 24596
rect 16540 24556 16546 24568
rect 16669 24565 16681 24568
rect 16715 24565 16727 24599
rect 17052 24596 17080 24704
rect 17221 24701 17233 24735
rect 17267 24732 17279 24735
rect 17862 24732 17868 24744
rect 17267 24704 17868 24732
rect 17267 24701 17279 24704
rect 17221 24695 17279 24701
rect 17862 24692 17868 24704
rect 17920 24692 17926 24744
rect 19242 24732 19248 24744
rect 18248 24704 19248 24732
rect 17954 24596 17960 24608
rect 17052 24568 17960 24596
rect 16669 24559 16727 24565
rect 17954 24556 17960 24568
rect 18012 24596 18018 24608
rect 18248 24596 18276 24704
rect 19242 24692 19248 24704
rect 19300 24692 19306 24744
rect 19702 24692 19708 24744
rect 19760 24692 19766 24744
rect 21266 24692 21272 24744
rect 21324 24692 21330 24744
rect 18414 24624 18420 24676
rect 18472 24664 18478 24676
rect 18693 24667 18751 24673
rect 18693 24664 18705 24667
rect 18472 24636 18705 24664
rect 18472 24624 18478 24636
rect 18693 24633 18705 24636
rect 18739 24664 18751 24667
rect 21560 24664 21588 24763
rect 21910 24760 21916 24812
rect 21968 24760 21974 24812
rect 22738 24760 22744 24812
rect 22796 24760 22802 24812
rect 24121 24735 24179 24741
rect 24121 24701 24133 24735
rect 24167 24701 24179 24735
rect 24121 24695 24179 24701
rect 18739 24636 19196 24664
rect 21560 24636 22876 24664
rect 18739 24633 18751 24636
rect 18693 24627 18751 24633
rect 19168 24608 19196 24636
rect 18012 24568 18276 24596
rect 18012 24556 18018 24568
rect 18782 24556 18788 24608
rect 18840 24596 18846 24608
rect 19061 24599 19119 24605
rect 19061 24596 19073 24599
rect 18840 24568 19073 24596
rect 18840 24556 18846 24568
rect 19061 24565 19073 24568
rect 19107 24565 19119 24599
rect 19061 24559 19119 24565
rect 19150 24556 19156 24608
rect 19208 24556 19214 24608
rect 19797 24599 19855 24605
rect 19797 24565 19809 24599
rect 19843 24596 19855 24599
rect 20622 24596 20628 24608
rect 19843 24568 20628 24596
rect 19843 24565 19855 24568
rect 19797 24559 19855 24565
rect 20622 24556 20628 24568
rect 20680 24556 20686 24608
rect 22005 24599 22063 24605
rect 22005 24565 22017 24599
rect 22051 24596 22063 24599
rect 22094 24596 22100 24608
rect 22051 24568 22100 24596
rect 22051 24565 22063 24568
rect 22005 24559 22063 24565
rect 22094 24556 22100 24568
rect 22152 24556 22158 24608
rect 22370 24556 22376 24608
rect 22428 24556 22434 24608
rect 22848 24596 22876 24636
rect 23382 24596 23388 24608
rect 22848 24568 23388 24596
rect 23382 24556 23388 24568
rect 23440 24596 23446 24608
rect 24136 24596 24164 24695
rect 23440 24568 24164 24596
rect 23440 24556 23446 24568
rect 1104 24506 26312 24528
rect 1104 24454 4101 24506
rect 4153 24454 4165 24506
rect 4217 24454 4229 24506
rect 4281 24454 4293 24506
rect 4345 24454 4357 24506
rect 4409 24454 10403 24506
rect 10455 24454 10467 24506
rect 10519 24454 10531 24506
rect 10583 24454 10595 24506
rect 10647 24454 10659 24506
rect 10711 24454 16705 24506
rect 16757 24454 16769 24506
rect 16821 24454 16833 24506
rect 16885 24454 16897 24506
rect 16949 24454 16961 24506
rect 17013 24454 23007 24506
rect 23059 24454 23071 24506
rect 23123 24454 23135 24506
rect 23187 24454 23199 24506
rect 23251 24454 23263 24506
rect 23315 24454 26312 24506
rect 1104 24432 26312 24454
rect 5813 24395 5871 24401
rect 5813 24361 5825 24395
rect 5859 24392 5871 24395
rect 7190 24392 7196 24404
rect 5859 24364 7196 24392
rect 5859 24361 5871 24364
rect 5813 24355 5871 24361
rect 7190 24352 7196 24364
rect 7248 24352 7254 24404
rect 9858 24352 9864 24404
rect 9916 24392 9922 24404
rect 10137 24395 10195 24401
rect 10137 24392 10149 24395
rect 9916 24364 10149 24392
rect 9916 24352 9922 24364
rect 10137 24361 10149 24364
rect 10183 24361 10195 24395
rect 10137 24355 10195 24361
rect 11054 24352 11060 24404
rect 11112 24352 11118 24404
rect 11698 24352 11704 24404
rect 11756 24392 11762 24404
rect 12069 24395 12127 24401
rect 12069 24392 12081 24395
rect 11756 24364 12081 24392
rect 11756 24352 11762 24364
rect 12069 24361 12081 24364
rect 12115 24361 12127 24395
rect 12069 24355 12127 24361
rect 13081 24395 13139 24401
rect 13081 24361 13093 24395
rect 13127 24392 13139 24395
rect 13262 24392 13268 24404
rect 13127 24364 13268 24392
rect 13127 24361 13139 24364
rect 13081 24355 13139 24361
rect 13262 24352 13268 24364
rect 13320 24352 13326 24404
rect 16380 24395 16438 24401
rect 16380 24361 16392 24395
rect 16426 24392 16438 24395
rect 16482 24392 16488 24404
rect 16426 24364 16488 24392
rect 16426 24361 16438 24364
rect 16380 24355 16438 24361
rect 16482 24352 16488 24364
rect 16540 24352 16546 24404
rect 17494 24352 17500 24404
rect 17552 24392 17558 24404
rect 17957 24395 18015 24401
rect 17957 24392 17969 24395
rect 17552 24364 17969 24392
rect 17552 24352 17558 24364
rect 17957 24361 17969 24364
rect 18003 24361 18015 24395
rect 17957 24355 18015 24361
rect 20806 24352 20812 24404
rect 20864 24352 20870 24404
rect 21266 24352 21272 24404
rect 21324 24392 21330 24404
rect 23477 24395 23535 24401
rect 23477 24392 23489 24395
rect 21324 24364 23489 24392
rect 21324 24352 21330 24364
rect 23477 24361 23489 24364
rect 23523 24361 23535 24395
rect 23477 24355 23535 24361
rect 9490 24284 9496 24336
rect 9548 24324 9554 24336
rect 11072 24324 11100 24352
rect 9548 24296 11100 24324
rect 9548 24284 9554 24296
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 8294 24256 8300 24268
rect 8251 24228 8300 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 8294 24216 8300 24228
rect 8352 24256 8358 24268
rect 9508 24256 9536 24284
rect 11072 24265 11100 24296
rect 11514 24284 11520 24336
rect 11572 24324 11578 24336
rect 15197 24327 15255 24333
rect 15197 24324 15209 24327
rect 11572 24296 12434 24324
rect 11572 24284 11578 24296
rect 8352 24228 9536 24256
rect 11057 24259 11115 24265
rect 8352 24216 8358 24228
rect 11057 24225 11069 24259
rect 11103 24225 11115 24259
rect 11057 24219 11115 24225
rect 11238 24216 11244 24268
rect 11296 24216 11302 24268
rect 12161 24259 12219 24265
rect 12161 24256 12173 24259
rect 11348 24228 12173 24256
rect 5442 24148 5448 24200
rect 5500 24188 5506 24200
rect 5629 24191 5687 24197
rect 5629 24188 5641 24191
rect 5500 24160 5641 24188
rect 5500 24148 5506 24160
rect 5629 24157 5641 24160
rect 5675 24157 5687 24191
rect 5629 24151 5687 24157
rect 5810 24148 5816 24200
rect 5868 24148 5874 24200
rect 10321 24191 10379 24197
rect 10321 24157 10333 24191
rect 10367 24188 10379 24191
rect 10965 24191 11023 24197
rect 10367 24160 10640 24188
rect 10367 24157 10379 24160
rect 10321 24151 10379 24157
rect 4430 24012 4436 24064
rect 4488 24052 4494 24064
rect 6454 24052 6460 24064
rect 4488 24024 6460 24052
rect 4488 24012 4494 24024
rect 6454 24012 6460 24024
rect 6512 24052 6518 24064
rect 6822 24052 6828 24064
rect 6512 24024 6828 24052
rect 6512 24012 6518 24024
rect 6822 24012 6828 24024
rect 6880 24012 6886 24064
rect 7098 24012 7104 24064
rect 7156 24052 7162 24064
rect 10612 24061 10640 24160
rect 10965 24157 10977 24191
rect 11011 24188 11023 24191
rect 11348 24188 11376 24228
rect 12161 24225 12173 24228
rect 12207 24225 12219 24259
rect 12406 24256 12434 24296
rect 14016 24296 15209 24324
rect 12713 24259 12771 24265
rect 12713 24256 12725 24259
rect 12406 24228 12725 24256
rect 12161 24219 12219 24225
rect 12713 24225 12725 24228
rect 12759 24225 12771 24259
rect 13265 24259 13323 24265
rect 13265 24256 13277 24259
rect 12713 24219 12771 24225
rect 12820 24228 13277 24256
rect 11011 24160 11376 24188
rect 11011 24157 11023 24160
rect 10965 24151 11023 24157
rect 11422 24148 11428 24200
rect 11480 24148 11486 24200
rect 11514 24148 11520 24200
rect 11572 24188 11578 24200
rect 11572 24160 11617 24188
rect 11572 24148 11578 24160
rect 11790 24148 11796 24200
rect 11848 24148 11854 24200
rect 11931 24191 11989 24197
rect 11931 24157 11943 24191
rect 11977 24188 11989 24191
rect 12066 24188 12072 24200
rect 11977 24160 12072 24188
rect 11977 24157 11989 24160
rect 11931 24151 11989 24157
rect 12066 24148 12072 24160
rect 12124 24148 12130 24200
rect 12342 24148 12348 24200
rect 12400 24188 12406 24200
rect 12820 24188 12848 24228
rect 13265 24225 13277 24228
rect 13311 24225 13323 24259
rect 14016 24256 14044 24296
rect 15197 24293 15209 24296
rect 15243 24293 15255 24327
rect 15197 24287 15255 24293
rect 17862 24284 17868 24336
rect 17920 24324 17926 24336
rect 18785 24327 18843 24333
rect 18785 24324 18797 24327
rect 17920 24296 18797 24324
rect 17920 24284 17926 24296
rect 18785 24293 18797 24296
rect 18831 24293 18843 24327
rect 18785 24287 18843 24293
rect 21637 24327 21695 24333
rect 21637 24293 21649 24327
rect 21683 24324 21695 24327
rect 21683 24296 22508 24324
rect 21683 24293 21695 24296
rect 21637 24287 21695 24293
rect 13265 24219 13323 24225
rect 13464 24228 14044 24256
rect 15013 24259 15071 24265
rect 12400 24160 12848 24188
rect 12897 24191 12955 24197
rect 12400 24148 12406 24160
rect 12897 24157 12909 24191
rect 12943 24188 12955 24191
rect 13464 24188 13492 24228
rect 15013 24225 15025 24259
rect 15059 24256 15071 24259
rect 15102 24256 15108 24268
rect 15059 24228 15108 24256
rect 15059 24225 15071 24228
rect 15013 24219 15071 24225
rect 15102 24216 15108 24228
rect 15160 24216 15166 24268
rect 15286 24216 15292 24268
rect 15344 24256 15350 24268
rect 15838 24256 15844 24268
rect 15344 24228 15844 24256
rect 15344 24216 15350 24228
rect 15838 24216 15844 24228
rect 15896 24216 15902 24268
rect 16117 24259 16175 24265
rect 16117 24225 16129 24259
rect 16163 24256 16175 24259
rect 18417 24259 18475 24265
rect 18417 24256 18429 24259
rect 16163 24228 18000 24256
rect 16163 24225 16175 24228
rect 16117 24219 16175 24225
rect 17972 24200 18000 24228
rect 18064 24228 18429 24256
rect 12943 24160 13492 24188
rect 13541 24191 13599 24197
rect 12943 24157 12955 24160
rect 12897 24151 12955 24157
rect 13541 24157 13553 24191
rect 13587 24188 13599 24191
rect 13814 24188 13820 24200
rect 13587 24160 13820 24188
rect 13587 24157 13599 24160
rect 13541 24151 13599 24157
rect 13814 24148 13820 24160
rect 13872 24148 13878 24200
rect 13906 24148 13912 24200
rect 13964 24188 13970 24200
rect 14277 24191 14335 24197
rect 14277 24188 14289 24191
rect 13964 24160 14289 24188
rect 13964 24148 13970 24160
rect 14277 24157 14289 24160
rect 14323 24157 14335 24191
rect 14277 24151 14335 24157
rect 14458 24148 14464 24200
rect 14516 24148 14522 24200
rect 15657 24191 15715 24197
rect 15657 24188 15669 24191
rect 14568 24160 15669 24188
rect 11701 24123 11759 24129
rect 11701 24089 11713 24123
rect 11747 24089 11759 24123
rect 12986 24120 12992 24132
rect 11701 24083 11759 24089
rect 11992 24092 12992 24120
rect 7561 24055 7619 24061
rect 7561 24052 7573 24055
rect 7156 24024 7573 24052
rect 7156 24012 7162 24024
rect 7561 24021 7573 24024
rect 7607 24021 7619 24055
rect 7561 24015 7619 24021
rect 10597 24055 10655 24061
rect 10597 24021 10609 24055
rect 10643 24021 10655 24055
rect 11716 24052 11744 24083
rect 11992 24052 12020 24092
rect 12986 24080 12992 24092
rect 13044 24080 13050 24132
rect 14568 24120 14596 24160
rect 15657 24157 15669 24160
rect 15703 24157 15715 24191
rect 17862 24188 17868 24200
rect 17526 24160 17868 24188
rect 15657 24151 15715 24157
rect 17862 24148 17868 24160
rect 17920 24148 17926 24200
rect 17954 24148 17960 24200
rect 18012 24148 18018 24200
rect 18064 24120 18092 24228
rect 18417 24225 18429 24228
rect 18463 24225 18475 24259
rect 18417 24219 18475 24225
rect 18598 24216 18604 24268
rect 18656 24216 18662 24268
rect 20257 24259 20315 24265
rect 20257 24225 20269 24259
rect 20303 24256 20315 24259
rect 21085 24259 21143 24265
rect 21085 24256 21097 24259
rect 20303 24228 21097 24256
rect 20303 24225 20315 24228
rect 20257 24219 20315 24225
rect 21085 24225 21097 24228
rect 21131 24225 21143 24259
rect 21085 24219 21143 24225
rect 18690 24148 18696 24200
rect 18748 24188 18754 24200
rect 18969 24191 19027 24197
rect 18969 24188 18981 24191
rect 18748 24160 18981 24188
rect 18748 24148 18754 24160
rect 18969 24157 18981 24160
rect 19015 24157 19027 24191
rect 18969 24151 19027 24157
rect 19797 24191 19855 24197
rect 19797 24157 19809 24191
rect 19843 24157 19855 24191
rect 21100 24188 21128 24219
rect 21174 24216 21180 24268
rect 21232 24216 21238 24268
rect 22002 24216 22008 24268
rect 22060 24216 22066 24268
rect 22480 24265 22508 24296
rect 22465 24259 22523 24265
rect 22465 24225 22477 24259
rect 22511 24225 22523 24259
rect 22465 24219 22523 24225
rect 23109 24259 23167 24265
rect 23109 24225 23121 24259
rect 23155 24256 23167 24259
rect 23155 24228 23704 24256
rect 23155 24225 23167 24228
rect 23109 24219 23167 24225
rect 22020 24188 22048 24216
rect 21100 24160 22048 24188
rect 19797 24151 19855 24157
rect 13464 24092 14596 24120
rect 17788 24092 18092 24120
rect 18325 24123 18383 24129
rect 13464 24064 13492 24092
rect 11716 24024 12020 24052
rect 10597 24015 10655 24021
rect 12526 24012 12532 24064
rect 12584 24052 12590 24064
rect 13446 24052 13452 24064
rect 12584 24024 13452 24052
rect 12584 24012 12590 24024
rect 13446 24012 13452 24024
rect 13504 24012 13510 24064
rect 13906 24012 13912 24064
rect 13964 24012 13970 24064
rect 14090 24012 14096 24064
rect 14148 24012 14154 24064
rect 15562 24012 15568 24064
rect 15620 24012 15626 24064
rect 17310 24012 17316 24064
rect 17368 24052 17374 24064
rect 17788 24052 17816 24092
rect 18325 24089 18337 24123
rect 18371 24120 18383 24123
rect 19245 24123 19303 24129
rect 19245 24120 19257 24123
rect 18371 24092 19257 24120
rect 18371 24089 18383 24092
rect 18325 24083 18383 24089
rect 19245 24089 19257 24092
rect 19291 24089 19303 24123
rect 19245 24083 19303 24089
rect 17368 24024 17816 24052
rect 17865 24055 17923 24061
rect 17368 24012 17374 24024
rect 17865 24021 17877 24055
rect 17911 24052 17923 24055
rect 19334 24052 19340 24064
rect 17911 24024 19340 24052
rect 17911 24021 17923 24024
rect 17865 24015 17923 24021
rect 19334 24012 19340 24024
rect 19392 24052 19398 24064
rect 19812 24052 19840 24151
rect 22186 24148 22192 24200
rect 22244 24188 22250 24200
rect 22281 24191 22339 24197
rect 22281 24188 22293 24191
rect 22244 24160 22293 24188
rect 22244 24148 22250 24160
rect 22281 24157 22293 24160
rect 22327 24157 22339 24191
rect 22281 24151 22339 24157
rect 22922 24148 22928 24200
rect 22980 24188 22986 24200
rect 23676 24197 23704 24228
rect 23201 24191 23259 24197
rect 23201 24188 23213 24191
rect 22980 24160 23213 24188
rect 22980 24148 22986 24160
rect 23201 24157 23213 24160
rect 23247 24157 23259 24191
rect 23201 24151 23259 24157
rect 23661 24191 23719 24197
rect 23661 24157 23673 24191
rect 23707 24157 23719 24191
rect 23661 24151 23719 24157
rect 21269 24123 21327 24129
rect 21269 24089 21281 24123
rect 21315 24120 21327 24123
rect 22094 24120 22100 24132
rect 21315 24092 22100 24120
rect 21315 24089 21327 24092
rect 21269 24083 21327 24089
rect 22094 24080 22100 24092
rect 22152 24080 22158 24132
rect 19392 24024 19840 24052
rect 19392 24012 19398 24024
rect 20346 24012 20352 24064
rect 20404 24012 20410 24064
rect 20441 24055 20499 24061
rect 20441 24021 20453 24055
rect 20487 24052 20499 24055
rect 20622 24052 20628 24064
rect 20487 24024 20628 24052
rect 20487 24021 20499 24024
rect 20441 24015 20499 24021
rect 20622 24012 20628 24024
rect 20680 24012 20686 24064
rect 21726 24012 21732 24064
rect 21784 24012 21790 24064
rect 23385 24055 23443 24061
rect 23385 24021 23397 24055
rect 23431 24052 23443 24055
rect 23658 24052 23664 24064
rect 23431 24024 23664 24052
rect 23431 24021 23443 24024
rect 23385 24015 23443 24021
rect 23658 24012 23664 24024
rect 23716 24012 23722 24064
rect 1104 23962 26472 23984
rect 1104 23910 7252 23962
rect 7304 23910 7316 23962
rect 7368 23910 7380 23962
rect 7432 23910 7444 23962
rect 7496 23910 7508 23962
rect 7560 23910 13554 23962
rect 13606 23910 13618 23962
rect 13670 23910 13682 23962
rect 13734 23910 13746 23962
rect 13798 23910 13810 23962
rect 13862 23910 19856 23962
rect 19908 23910 19920 23962
rect 19972 23910 19984 23962
rect 20036 23910 20048 23962
rect 20100 23910 20112 23962
rect 20164 23910 26158 23962
rect 26210 23910 26222 23962
rect 26274 23910 26286 23962
rect 26338 23910 26350 23962
rect 26402 23910 26414 23962
rect 26466 23910 26472 23962
rect 1104 23888 26472 23910
rect 4706 23808 4712 23860
rect 4764 23848 4770 23860
rect 5261 23851 5319 23857
rect 5261 23848 5273 23851
rect 4764 23820 5273 23848
rect 4764 23808 4770 23820
rect 5261 23817 5273 23820
rect 5307 23817 5319 23851
rect 5261 23811 5319 23817
rect 7650 23808 7656 23860
rect 7708 23848 7714 23860
rect 7708 23820 7972 23848
rect 7708 23808 7714 23820
rect 5169 23783 5227 23789
rect 4724 23752 5120 23780
rect 4724 23656 4752 23752
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23712 4859 23715
rect 5092 23713 5120 23752
rect 5169 23749 5181 23783
rect 5215 23780 5227 23783
rect 6089 23783 6147 23789
rect 6089 23780 6101 23783
rect 5215 23752 6101 23780
rect 5215 23749 5227 23752
rect 5169 23743 5227 23749
rect 6089 23749 6101 23752
rect 6135 23749 6147 23783
rect 6089 23743 6147 23749
rect 5092 23712 5212 23713
rect 4847 23684 5028 23712
rect 5092 23685 5304 23712
rect 5184 23684 5304 23685
rect 4847 23681 4859 23684
rect 4801 23675 4859 23681
rect 5000 23656 5028 23684
rect 4706 23604 4712 23656
rect 4764 23604 4770 23656
rect 4982 23604 4988 23656
rect 5040 23604 5046 23656
rect 5077 23647 5135 23653
rect 5077 23613 5089 23647
rect 5123 23613 5135 23647
rect 5276 23644 5304 23684
rect 5350 23672 5356 23724
rect 5408 23712 5414 23724
rect 5997 23715 6055 23721
rect 5997 23712 6009 23715
rect 5408 23684 6009 23712
rect 5408 23672 5414 23684
rect 5997 23681 6009 23684
rect 6043 23681 6055 23715
rect 5997 23675 6055 23681
rect 6454 23672 6460 23724
rect 6512 23672 6518 23724
rect 7944 23698 7972 23820
rect 8294 23808 8300 23860
rect 8352 23808 8358 23860
rect 14090 23848 14096 23860
rect 13464 23820 14096 23848
rect 13464 23789 13492 23820
rect 14090 23808 14096 23820
rect 14148 23808 14154 23860
rect 14918 23808 14924 23860
rect 14976 23808 14982 23860
rect 15194 23808 15200 23860
rect 15252 23808 15258 23860
rect 15562 23808 15568 23860
rect 15620 23848 15626 23860
rect 15841 23851 15899 23857
rect 15841 23848 15853 23851
rect 15620 23820 15853 23848
rect 15620 23808 15626 23820
rect 15841 23817 15853 23820
rect 15887 23817 15899 23851
rect 17954 23848 17960 23860
rect 15841 23811 15899 23817
rect 16684 23820 17960 23848
rect 13449 23783 13507 23789
rect 13449 23749 13461 23783
rect 13495 23749 13507 23783
rect 15102 23780 15108 23792
rect 14674 23752 15108 23780
rect 13449 23743 13507 23749
rect 14936 23724 14964 23752
rect 15102 23740 15108 23752
rect 15160 23740 15166 23792
rect 9030 23672 9036 23724
rect 9088 23712 9094 23724
rect 9088 23684 9168 23712
rect 9088 23672 9094 23684
rect 5442 23644 5448 23656
rect 5276 23616 5448 23644
rect 5077 23607 5135 23613
rect 4522 23468 4528 23520
rect 4580 23468 4586 23520
rect 5092 23508 5120 23607
rect 5442 23604 5448 23616
rect 5500 23644 5506 23656
rect 5813 23647 5871 23653
rect 5813 23644 5825 23647
rect 5500 23616 5825 23644
rect 5500 23604 5506 23616
rect 5813 23613 5825 23616
rect 5859 23613 5871 23647
rect 6472 23644 6500 23672
rect 6549 23647 6607 23653
rect 6549 23644 6561 23647
rect 6472 23616 6561 23644
rect 5813 23607 5871 23613
rect 6549 23613 6561 23616
rect 6595 23613 6607 23647
rect 6549 23607 6607 23613
rect 6825 23647 6883 23653
rect 6825 23613 6837 23647
rect 6871 23644 6883 23647
rect 6914 23644 6920 23656
rect 6871 23616 6920 23644
rect 6871 23613 6883 23616
rect 6825 23607 6883 23613
rect 6914 23604 6920 23616
rect 6972 23604 6978 23656
rect 9140 23644 9168 23684
rect 9306 23672 9312 23724
rect 9364 23672 9370 23724
rect 10781 23715 10839 23721
rect 10781 23681 10793 23715
rect 10827 23712 10839 23715
rect 11514 23712 11520 23724
rect 10827 23684 11520 23712
rect 10827 23681 10839 23684
rect 10781 23675 10839 23681
rect 11514 23672 11520 23684
rect 11572 23672 11578 23724
rect 12897 23715 12955 23721
rect 12897 23681 12909 23715
rect 12943 23712 12955 23715
rect 13078 23712 13084 23724
rect 12943 23684 13084 23712
rect 12943 23681 12955 23684
rect 12897 23675 12955 23681
rect 13078 23672 13084 23684
rect 13136 23672 13142 23724
rect 13170 23672 13176 23724
rect 13228 23672 13234 23724
rect 14918 23672 14924 23724
rect 14976 23672 14982 23724
rect 15212 23721 15240 23808
rect 16684 23721 16712 23820
rect 17954 23808 17960 23820
rect 18012 23808 18018 23860
rect 18064 23820 18276 23848
rect 15197 23715 15255 23721
rect 15197 23681 15209 23715
rect 15243 23681 15255 23715
rect 15197 23675 15255 23681
rect 16669 23715 16727 23721
rect 16669 23681 16681 23715
rect 16715 23681 16727 23715
rect 16669 23675 16727 23681
rect 17954 23672 17960 23724
rect 18012 23712 18018 23724
rect 18064 23712 18092 23820
rect 18248 23792 18276 23820
rect 19702 23808 19708 23860
rect 19760 23848 19766 23860
rect 19981 23851 20039 23857
rect 19981 23848 19993 23851
rect 19760 23820 19993 23848
rect 19760 23808 19766 23820
rect 19981 23817 19993 23820
rect 20027 23817 20039 23851
rect 19981 23811 20039 23817
rect 20349 23851 20407 23857
rect 20349 23817 20361 23851
rect 20395 23848 20407 23851
rect 21269 23851 21327 23857
rect 21269 23848 21281 23851
rect 20395 23820 21281 23848
rect 20395 23817 20407 23820
rect 20349 23811 20407 23817
rect 21269 23817 21281 23820
rect 21315 23848 21327 23851
rect 21726 23848 21732 23860
rect 21315 23820 21732 23848
rect 21315 23817 21327 23820
rect 21269 23811 21327 23817
rect 21726 23808 21732 23820
rect 21784 23808 21790 23860
rect 22646 23808 22652 23860
rect 22704 23808 22710 23860
rect 23658 23808 23664 23860
rect 23716 23848 23722 23860
rect 23716 23820 23980 23848
rect 23716 23808 23722 23820
rect 18230 23740 18236 23792
rect 18288 23740 18294 23792
rect 19150 23740 19156 23792
rect 19208 23780 19214 23792
rect 19613 23783 19671 23789
rect 19613 23780 19625 23783
rect 19208 23752 19625 23780
rect 19208 23740 19214 23752
rect 19613 23749 19625 23752
rect 19659 23749 19671 23783
rect 19613 23743 19671 23749
rect 21177 23783 21235 23789
rect 21177 23749 21189 23783
rect 21223 23780 21235 23783
rect 22664 23780 22692 23808
rect 23952 23789 23980 23820
rect 21223 23752 22692 23780
rect 23937 23783 23995 23789
rect 21223 23749 21235 23752
rect 21177 23743 21235 23749
rect 23937 23749 23949 23783
rect 23983 23749 23995 23783
rect 23937 23743 23995 23749
rect 19061 23715 19119 23721
rect 19061 23712 19073 23715
rect 18012 23698 18092 23712
rect 18012 23684 18078 23698
rect 18432 23684 19073 23712
rect 18012 23672 18018 23684
rect 12526 23644 12532 23656
rect 9140 23616 12532 23644
rect 12526 23604 12532 23616
rect 12584 23604 12590 23656
rect 12618 23604 12624 23656
rect 12676 23604 12682 23656
rect 16945 23647 17003 23653
rect 16945 23613 16957 23647
rect 16991 23644 17003 23647
rect 17034 23644 17040 23656
rect 16991 23616 17040 23644
rect 16991 23613 17003 23616
rect 16945 23607 17003 23613
rect 17034 23604 17040 23616
rect 17092 23604 17098 23656
rect 17310 23604 17316 23656
rect 17368 23644 17374 23656
rect 18432 23653 18460 23684
rect 19061 23681 19073 23684
rect 19107 23681 19119 23715
rect 19061 23675 19119 23681
rect 19245 23715 19303 23721
rect 19245 23681 19257 23715
rect 19291 23681 19303 23715
rect 19245 23675 19303 23681
rect 18417 23647 18475 23653
rect 18417 23644 18429 23647
rect 17368 23616 18429 23644
rect 17368 23604 17374 23616
rect 18417 23613 18429 23616
rect 18463 23613 18475 23647
rect 18417 23607 18475 23613
rect 18966 23604 18972 23656
rect 19024 23644 19030 23656
rect 19260 23644 19288 23675
rect 19334 23672 19340 23724
rect 19392 23712 19398 23724
rect 19521 23715 19579 23721
rect 19392 23684 19437 23712
rect 19392 23672 19398 23684
rect 19521 23681 19533 23715
rect 19567 23681 19579 23715
rect 19710 23715 19768 23721
rect 19710 23712 19722 23715
rect 19521 23675 19579 23681
rect 19628 23684 19722 23712
rect 19024 23616 19288 23644
rect 19024 23604 19030 23616
rect 19536 23576 19564 23675
rect 18892 23548 19564 23576
rect 18892 23520 18920 23548
rect 6270 23508 6276 23520
rect 5092 23480 6276 23508
rect 6270 23468 6276 23480
rect 6328 23468 6334 23520
rect 8389 23511 8447 23517
rect 8389 23477 8401 23511
rect 8435 23508 8447 23511
rect 8478 23508 8484 23520
rect 8435 23480 8484 23508
rect 8435 23477 8447 23480
rect 8389 23471 8447 23477
rect 8478 23468 8484 23480
rect 8536 23468 8542 23520
rect 9122 23468 9128 23520
rect 9180 23468 9186 23520
rect 10318 23468 10324 23520
rect 10376 23508 10382 23520
rect 10597 23511 10655 23517
rect 10597 23508 10609 23511
rect 10376 23480 10609 23508
rect 10376 23468 10382 23480
rect 10597 23477 10609 23480
rect 10643 23477 10655 23511
rect 10597 23471 10655 23477
rect 11974 23468 11980 23520
rect 12032 23468 12038 23520
rect 12986 23468 12992 23520
rect 13044 23508 13050 23520
rect 13446 23508 13452 23520
rect 13044 23480 13452 23508
rect 13044 23468 13050 23480
rect 13446 23468 13452 23480
rect 13504 23468 13510 23520
rect 15930 23468 15936 23520
rect 15988 23508 15994 23520
rect 18138 23508 18144 23520
rect 15988 23480 18144 23508
rect 15988 23468 15994 23480
rect 18138 23468 18144 23480
rect 18196 23468 18202 23520
rect 18506 23468 18512 23520
rect 18564 23468 18570 23520
rect 18874 23468 18880 23520
rect 18932 23468 18938 23520
rect 19058 23468 19064 23520
rect 19116 23508 19122 23520
rect 19628 23508 19656 23684
rect 19710 23681 19722 23684
rect 19756 23681 19768 23715
rect 19710 23675 19768 23681
rect 20346 23672 20352 23724
rect 20404 23672 20410 23724
rect 20441 23715 20499 23721
rect 20441 23681 20453 23715
rect 20487 23712 20499 23715
rect 20806 23712 20812 23724
rect 20487 23684 20812 23712
rect 20487 23681 20499 23684
rect 20441 23675 20499 23681
rect 20806 23672 20812 23684
rect 20864 23672 20870 23724
rect 22094 23672 22100 23724
rect 22152 23712 22158 23724
rect 22152 23684 22324 23712
rect 22152 23672 22158 23684
rect 20364 23576 20392 23672
rect 20625 23647 20683 23653
rect 20625 23613 20637 23647
rect 20671 23644 20683 23647
rect 21453 23647 21511 23653
rect 21453 23644 21465 23647
rect 20671 23616 21465 23644
rect 20671 23613 20683 23616
rect 20625 23607 20683 23613
rect 21453 23613 21465 23616
rect 21499 23644 21511 23647
rect 22002 23644 22008 23656
rect 21499 23616 22008 23644
rect 21499 23613 21511 23616
rect 21453 23607 21511 23613
rect 22002 23604 22008 23616
rect 22060 23604 22066 23656
rect 22189 23647 22247 23653
rect 22189 23613 22201 23647
rect 22235 23613 22247 23647
rect 22296 23644 22324 23684
rect 22370 23672 22376 23724
rect 22428 23672 22434 23724
rect 22646 23672 22652 23724
rect 22704 23712 22710 23724
rect 22704 23684 22862 23712
rect 22704 23672 22710 23684
rect 22465 23647 22523 23653
rect 22465 23644 22477 23647
rect 22296 23616 22477 23644
rect 22189 23607 22247 23613
rect 22465 23613 22477 23616
rect 22511 23644 22523 23647
rect 22738 23644 22744 23656
rect 22511 23616 22744 23644
rect 22511 23613 22523 23616
rect 22465 23607 22523 23613
rect 22204 23576 22232 23607
rect 22738 23604 22744 23616
rect 22796 23604 22802 23656
rect 24213 23647 24271 23653
rect 24213 23613 24225 23647
rect 24259 23613 24271 23647
rect 24213 23607 24271 23613
rect 22646 23576 22652 23588
rect 20364 23548 22140 23576
rect 22204 23548 22652 23576
rect 19116 23480 19656 23508
rect 19116 23468 19122 23480
rect 19886 23468 19892 23520
rect 19944 23468 19950 23520
rect 20070 23468 20076 23520
rect 20128 23508 20134 23520
rect 20809 23511 20867 23517
rect 20809 23508 20821 23511
rect 20128 23480 20821 23508
rect 20128 23468 20134 23480
rect 20809 23477 20821 23480
rect 20855 23477 20867 23511
rect 20809 23471 20867 23477
rect 21910 23468 21916 23520
rect 21968 23468 21974 23520
rect 22112 23517 22140 23548
rect 22646 23536 22652 23548
rect 22704 23536 22710 23588
rect 22097 23511 22155 23517
rect 22097 23477 22109 23511
rect 22143 23508 22155 23511
rect 22554 23508 22560 23520
rect 22143 23480 22560 23508
rect 22143 23477 22155 23480
rect 22097 23471 22155 23477
rect 22554 23468 22560 23480
rect 22612 23468 22618 23520
rect 23382 23468 23388 23520
rect 23440 23508 23446 23520
rect 24228 23508 24256 23607
rect 23440 23480 24256 23508
rect 23440 23468 23446 23480
rect 1104 23418 26312 23440
rect 1104 23366 4101 23418
rect 4153 23366 4165 23418
rect 4217 23366 4229 23418
rect 4281 23366 4293 23418
rect 4345 23366 4357 23418
rect 4409 23366 10403 23418
rect 10455 23366 10467 23418
rect 10519 23366 10531 23418
rect 10583 23366 10595 23418
rect 10647 23366 10659 23418
rect 10711 23366 16705 23418
rect 16757 23366 16769 23418
rect 16821 23366 16833 23418
rect 16885 23366 16897 23418
rect 16949 23366 16961 23418
rect 17013 23366 23007 23418
rect 23059 23366 23071 23418
rect 23123 23366 23135 23418
rect 23187 23366 23199 23418
rect 23251 23366 23263 23418
rect 23315 23366 26312 23418
rect 1104 23344 26312 23366
rect 6454 23264 6460 23316
rect 6512 23304 6518 23316
rect 8757 23307 8815 23313
rect 6512 23276 7052 23304
rect 6512 23264 6518 23276
rect 6914 23196 6920 23248
rect 6972 23196 6978 23248
rect 4065 23171 4123 23177
rect 4065 23137 4077 23171
rect 4111 23168 4123 23171
rect 4430 23168 4436 23180
rect 4111 23140 4436 23168
rect 4111 23137 4123 23140
rect 4065 23131 4123 23137
rect 4430 23128 4436 23140
rect 4488 23128 4494 23180
rect 7024 23177 7052 23276
rect 8757 23273 8769 23307
rect 8803 23304 8815 23307
rect 9030 23304 9036 23316
rect 8803 23276 9036 23304
rect 8803 23273 8815 23276
rect 8757 23267 8815 23273
rect 9030 23264 9036 23276
rect 9088 23264 9094 23316
rect 10318 23264 10324 23316
rect 10376 23264 10382 23316
rect 12066 23264 12072 23316
rect 12124 23304 12130 23316
rect 12802 23304 12808 23316
rect 12124 23276 12808 23304
rect 12124 23264 12130 23276
rect 12802 23264 12808 23276
rect 12860 23304 12866 23316
rect 16022 23304 16028 23316
rect 12860 23276 16028 23304
rect 12860 23264 12866 23276
rect 16022 23264 16028 23276
rect 16080 23264 16086 23316
rect 16577 23307 16635 23313
rect 16577 23273 16589 23307
rect 16623 23304 16635 23307
rect 17034 23304 17040 23316
rect 16623 23276 17040 23304
rect 16623 23273 16635 23276
rect 16577 23267 16635 23273
rect 17034 23264 17040 23276
rect 17092 23264 17098 23316
rect 18049 23307 18107 23313
rect 18049 23273 18061 23307
rect 18095 23304 18107 23307
rect 18690 23304 18696 23316
rect 18095 23276 18696 23304
rect 18095 23273 18107 23276
rect 18049 23267 18107 23273
rect 18690 23264 18696 23276
rect 18748 23264 18754 23316
rect 20070 23304 20076 23316
rect 18892 23276 20076 23304
rect 7009 23171 7067 23177
rect 7009 23137 7021 23171
rect 7055 23168 7067 23171
rect 8294 23168 8300 23180
rect 7055 23140 8300 23168
rect 7055 23137 7067 23140
rect 7009 23131 7067 23137
rect 8294 23128 8300 23140
rect 8352 23168 8358 23180
rect 9033 23171 9091 23177
rect 9033 23168 9045 23171
rect 8352 23140 9045 23168
rect 8352 23128 8358 23140
rect 9033 23137 9045 23140
rect 9079 23137 9091 23171
rect 10336 23168 10364 23264
rect 10505 23171 10563 23177
rect 10505 23168 10517 23171
rect 10336 23140 10517 23168
rect 9033 23131 9091 23137
rect 10505 23137 10517 23140
rect 10551 23137 10563 23171
rect 10505 23131 10563 23137
rect 11977 23171 12035 23177
rect 11977 23137 11989 23171
rect 12023 23168 12035 23171
rect 12618 23168 12624 23180
rect 12023 23140 12624 23168
rect 12023 23137 12035 23140
rect 11977 23131 12035 23137
rect 12618 23128 12624 23140
rect 12676 23168 12682 23180
rect 13354 23168 13360 23180
rect 12676 23140 13360 23168
rect 12676 23128 12682 23140
rect 13354 23128 13360 23140
rect 13412 23128 13418 23180
rect 16206 23128 16212 23180
rect 16264 23128 16270 23180
rect 17310 23128 17316 23180
rect 17368 23128 17374 23180
rect 17402 23128 17408 23180
rect 17460 23128 17466 23180
rect 5442 23060 5448 23112
rect 5500 23100 5506 23112
rect 5994 23100 6000 23112
rect 5500 23072 6000 23100
rect 5500 23060 5506 23072
rect 5994 23060 6000 23072
rect 6052 23060 6058 23112
rect 6365 23103 6423 23109
rect 6365 23069 6377 23103
rect 6411 23069 6423 23103
rect 6365 23063 6423 23069
rect 6733 23103 6791 23109
rect 6733 23069 6745 23103
rect 6779 23100 6791 23103
rect 6914 23100 6920 23112
rect 6779 23072 6920 23100
rect 6779 23069 6791 23072
rect 6733 23063 6791 23069
rect 4341 23035 4399 23041
rect 4341 23001 4353 23035
rect 4387 23001 4399 23035
rect 4341 22995 4399 23001
rect 6089 23035 6147 23041
rect 6089 23001 6101 23035
rect 6135 23032 6147 23035
rect 6270 23032 6276 23044
rect 6135 23004 6276 23032
rect 6135 23001 6147 23004
rect 6089 22995 6147 23001
rect 4356 22964 4384 22995
rect 6270 22992 6276 23004
rect 6328 22992 6334 23044
rect 4522 22964 4528 22976
rect 4356 22936 4528 22964
rect 4522 22924 4528 22936
rect 4580 22924 4586 22976
rect 6380 22964 6408 23063
rect 6914 23060 6920 23072
rect 6972 23060 6978 23112
rect 10226 23060 10232 23112
rect 10284 23060 10290 23112
rect 12529 23103 12587 23109
rect 6546 22992 6552 23044
rect 6604 22992 6610 23044
rect 6641 23035 6699 23041
rect 6641 23001 6653 23035
rect 6687 23032 6699 23035
rect 7190 23032 7196 23044
rect 6687 23004 7196 23032
rect 6687 23001 6699 23004
rect 6641 22995 6699 23001
rect 7190 22992 7196 23004
rect 7248 22992 7254 23044
rect 7285 23035 7343 23041
rect 7285 23001 7297 23035
rect 7331 23001 7343 23035
rect 9861 23035 9919 23041
rect 7285 22995 7343 23001
rect 7668 23004 7774 23032
rect 6822 22964 6828 22976
rect 6380 22936 6828 22964
rect 6822 22924 6828 22936
rect 6880 22924 6886 22976
rect 7098 22924 7104 22976
rect 7156 22964 7162 22976
rect 7300 22964 7328 22995
rect 7668 22976 7696 23004
rect 9861 23001 9873 23035
rect 9907 23032 9919 23035
rect 10134 23032 10140 23044
rect 9907 23004 10140 23032
rect 9907 23001 9919 23004
rect 9861 22995 9919 23001
rect 10134 22992 10140 23004
rect 10192 22992 10198 23044
rect 7156 22936 7328 22964
rect 7156 22924 7162 22936
rect 7650 22924 7656 22976
rect 7708 22924 7714 22976
rect 10870 22924 10876 22976
rect 10928 22964 10934 22976
rect 11422 22964 11428 22976
rect 10928 22936 11428 22964
rect 10928 22924 10934 22936
rect 11422 22924 11428 22936
rect 11480 22964 11486 22976
rect 11624 22964 11652 23086
rect 12529 23069 12541 23103
rect 12575 23069 12587 23103
rect 12529 23063 12587 23069
rect 11480 22936 11652 22964
rect 12544 22964 12572 23063
rect 12802 23060 12808 23112
rect 12860 23060 12866 23112
rect 12894 23060 12900 23112
rect 12952 23060 12958 23112
rect 13078 23060 13084 23112
rect 13136 23060 13142 23112
rect 16025 23103 16083 23109
rect 16025 23069 16037 23103
rect 16071 23100 16083 23103
rect 16224 23100 16252 23128
rect 16071 23072 16252 23100
rect 16071 23069 16083 23072
rect 16025 23063 16083 23069
rect 16390 23060 16396 23112
rect 16448 23060 16454 23112
rect 17328 23100 17356 23128
rect 17589 23103 17647 23109
rect 17589 23100 17601 23103
rect 17328 23072 17601 23100
rect 17589 23069 17601 23072
rect 17635 23069 17647 23103
rect 17589 23063 17647 23069
rect 17681 23103 17739 23109
rect 17681 23069 17693 23103
rect 17727 23100 17739 23103
rect 17770 23100 17776 23112
rect 17727 23072 17776 23100
rect 17727 23069 17739 23072
rect 17681 23063 17739 23069
rect 17770 23060 17776 23072
rect 17828 23060 17834 23112
rect 18506 23060 18512 23112
rect 18564 23060 18570 23112
rect 18601 23103 18659 23109
rect 18601 23069 18613 23103
rect 18647 23100 18659 23103
rect 18782 23100 18788 23112
rect 18647 23072 18788 23100
rect 18647 23069 18659 23072
rect 18601 23063 18659 23069
rect 18782 23060 18788 23072
rect 18840 23060 18846 23112
rect 18892 23109 18920 23276
rect 20070 23264 20076 23276
rect 20128 23264 20134 23316
rect 22002 23264 22008 23316
rect 22060 23264 22066 23316
rect 22097 23307 22155 23313
rect 22097 23273 22109 23307
rect 22143 23273 22155 23307
rect 22097 23267 22155 23273
rect 22281 23307 22339 23313
rect 22281 23273 22293 23307
rect 22327 23304 22339 23307
rect 22370 23304 22376 23316
rect 22327 23276 22376 23304
rect 22327 23273 22339 23276
rect 22281 23267 22339 23273
rect 20622 23196 20628 23248
rect 20680 23236 20686 23248
rect 20680 23208 21956 23236
rect 20680 23196 20686 23208
rect 20254 23128 20260 23180
rect 20312 23168 20318 23180
rect 21928 23177 21956 23208
rect 20993 23171 21051 23177
rect 20312 23140 20760 23168
rect 20312 23128 20318 23140
rect 18877 23103 18935 23109
rect 18877 23069 18889 23103
rect 18923 23069 18935 23103
rect 18877 23063 18935 23069
rect 19242 23060 19248 23112
rect 19300 23060 19306 23112
rect 20732 23100 20760 23140
rect 20993 23137 21005 23171
rect 21039 23168 21051 23171
rect 21913 23171 21971 23177
rect 21039 23140 21772 23168
rect 21039 23137 21051 23140
rect 20993 23131 21051 23137
rect 21637 23103 21695 23109
rect 21637 23100 21649 23103
rect 20732 23072 21649 23100
rect 21637 23069 21649 23072
rect 21683 23069 21695 23103
rect 21744 23100 21772 23140
rect 21913 23137 21925 23171
rect 21959 23137 21971 23171
rect 22020 23168 22048 23264
rect 22112 23236 22140 23267
rect 22370 23264 22376 23276
rect 22428 23264 22434 23316
rect 22922 23264 22928 23316
rect 22980 23304 22986 23316
rect 23293 23307 23351 23313
rect 23293 23304 23305 23307
rect 22980 23276 23305 23304
rect 22980 23264 22986 23276
rect 23293 23273 23305 23276
rect 23339 23273 23351 23307
rect 23293 23267 23351 23273
rect 22554 23236 22560 23248
rect 22112 23208 22560 23236
rect 22554 23196 22560 23208
rect 22612 23236 22618 23248
rect 22612 23208 24164 23236
rect 22612 23196 22618 23208
rect 22649 23171 22707 23177
rect 22649 23168 22661 23171
rect 22020 23140 22661 23168
rect 21913 23131 21971 23137
rect 22649 23137 22661 23140
rect 22695 23137 22707 23171
rect 22649 23131 22707 23137
rect 22097 23103 22155 23109
rect 22097 23100 22109 23103
rect 21744 23072 22109 23100
rect 21637 23063 21695 23069
rect 22097 23069 22109 23072
rect 22143 23100 22155 23103
rect 22186 23100 22192 23112
rect 22143 23072 22192 23100
rect 22143 23069 22155 23072
rect 22097 23063 22155 23069
rect 22186 23060 22192 23072
rect 22244 23060 22250 23112
rect 12912 23032 12940 23060
rect 15930 23032 15936 23044
rect 12912 23004 15936 23032
rect 15930 22992 15936 23004
rect 15988 22992 15994 23044
rect 16209 23035 16267 23041
rect 16209 23001 16221 23035
rect 16255 23001 16267 23035
rect 16209 22995 16267 23001
rect 15470 22964 15476 22976
rect 12544 22936 15476 22964
rect 11480 22924 11486 22936
rect 15470 22924 15476 22936
rect 15528 22964 15534 22976
rect 15838 22964 15844 22976
rect 15528 22936 15844 22964
rect 15528 22924 15534 22936
rect 15838 22924 15844 22936
rect 15896 22924 15902 22976
rect 16224 22964 16252 22995
rect 16298 22992 16304 23044
rect 16356 22992 16362 23044
rect 18524 23032 18552 23060
rect 19521 23035 19579 23041
rect 19521 23032 19533 23035
rect 16408 23004 18552 23032
rect 19076 23004 19533 23032
rect 16408 22964 16436 23004
rect 16224 22936 16436 22964
rect 18782 22924 18788 22976
rect 18840 22924 18846 22976
rect 19076 22973 19104 23004
rect 19521 23001 19533 23004
rect 19567 23001 19579 23035
rect 20990 23032 20996 23044
rect 20746 23004 20996 23032
rect 19521 22995 19579 23001
rect 20990 22992 20996 23004
rect 21048 23032 21054 23044
rect 21048 23004 21220 23032
rect 21048 22992 21054 23004
rect 19061 22967 19119 22973
rect 19061 22933 19073 22967
rect 19107 22933 19119 22967
rect 19061 22927 19119 22933
rect 21082 22924 21088 22976
rect 21140 22924 21146 22976
rect 21192 22964 21220 23004
rect 21450 22992 21456 23044
rect 21508 23032 21514 23044
rect 21821 23035 21879 23041
rect 21821 23032 21833 23035
rect 21508 23004 21833 23032
rect 21508 22992 21514 23004
rect 21821 23001 21833 23004
rect 21867 23001 21879 23035
rect 21821 22995 21879 23001
rect 22462 22964 22468 22976
rect 21192 22936 22468 22964
rect 22462 22924 22468 22936
rect 22520 22924 22526 22976
rect 22664 22964 22692 23131
rect 22738 23128 22744 23180
rect 22796 23168 22802 23180
rect 24136 23177 24164 23208
rect 22833 23171 22891 23177
rect 22833 23168 22845 23171
rect 22796 23140 22845 23168
rect 22796 23128 22802 23140
rect 22833 23137 22845 23140
rect 22879 23137 22891 23171
rect 22833 23131 22891 23137
rect 24121 23171 24179 23177
rect 24121 23137 24133 23171
rect 24167 23137 24179 23171
rect 24121 23131 24179 23137
rect 22738 22964 22744 22976
rect 22664 22936 22744 22964
rect 22738 22924 22744 22936
rect 22796 22924 22802 22976
rect 22925 22967 22983 22973
rect 22925 22933 22937 22967
rect 22971 22964 22983 22967
rect 23569 22967 23627 22973
rect 23569 22964 23581 22967
rect 22971 22936 23581 22964
rect 22971 22933 22983 22936
rect 22925 22927 22983 22933
rect 23569 22933 23581 22936
rect 23615 22933 23627 22967
rect 23569 22927 23627 22933
rect 1104 22874 26472 22896
rect 1104 22822 7252 22874
rect 7304 22822 7316 22874
rect 7368 22822 7380 22874
rect 7432 22822 7444 22874
rect 7496 22822 7508 22874
rect 7560 22822 13554 22874
rect 13606 22822 13618 22874
rect 13670 22822 13682 22874
rect 13734 22822 13746 22874
rect 13798 22822 13810 22874
rect 13862 22822 19856 22874
rect 19908 22822 19920 22874
rect 19972 22822 19984 22874
rect 20036 22822 20048 22874
rect 20100 22822 20112 22874
rect 20164 22822 26158 22874
rect 26210 22822 26222 22874
rect 26274 22822 26286 22874
rect 26338 22822 26350 22874
rect 26402 22822 26414 22874
rect 26466 22822 26472 22874
rect 1104 22800 26472 22822
rect 3142 22720 3148 22772
rect 3200 22760 3206 22772
rect 4893 22763 4951 22769
rect 3200 22732 4292 22760
rect 3200 22720 3206 22732
rect 4264 22692 4292 22732
rect 4893 22729 4905 22763
rect 4939 22760 4951 22763
rect 5350 22760 5356 22772
rect 4939 22732 5356 22760
rect 4939 22729 4951 22732
rect 4893 22723 4951 22729
rect 5350 22720 5356 22732
rect 5408 22720 5414 22772
rect 7098 22720 7104 22772
rect 7156 22760 7162 22772
rect 7285 22763 7343 22769
rect 7285 22760 7297 22763
rect 7156 22732 7297 22760
rect 7156 22720 7162 22732
rect 7285 22729 7297 22732
rect 7331 22729 7343 22763
rect 7285 22723 7343 22729
rect 8294 22720 8300 22772
rect 8352 22720 8358 22772
rect 9122 22760 9128 22772
rect 8496 22732 9128 22760
rect 5442 22692 5448 22704
rect 4186 22664 5448 22692
rect 5442 22652 5448 22664
rect 5500 22652 5506 22704
rect 6178 22652 6184 22704
rect 6236 22692 6242 22704
rect 6917 22695 6975 22701
rect 6917 22692 6929 22695
rect 6236 22664 6929 22692
rect 6236 22652 6242 22664
rect 6917 22661 6929 22664
rect 6963 22661 6975 22695
rect 8312 22692 8340 22720
rect 8496 22701 8524 22732
rect 9122 22720 9128 22732
rect 9180 22720 9186 22772
rect 11514 22720 11520 22772
rect 11572 22720 11578 22772
rect 11885 22763 11943 22769
rect 11885 22729 11897 22763
rect 11931 22760 11943 22763
rect 11974 22760 11980 22772
rect 11931 22732 11980 22760
rect 11931 22729 11943 22732
rect 11885 22723 11943 22729
rect 11974 22720 11980 22732
rect 12032 22720 12038 22772
rect 14826 22720 14832 22772
rect 14884 22760 14890 22772
rect 16298 22760 16304 22772
rect 14884 22732 16304 22760
rect 14884 22720 14890 22732
rect 16298 22720 16304 22732
rect 16356 22720 16362 22772
rect 16390 22720 16396 22772
rect 16448 22720 16454 22772
rect 18782 22720 18788 22772
rect 18840 22760 18846 22772
rect 18840 22732 19380 22760
rect 18840 22720 18846 22732
rect 6917 22655 6975 22661
rect 8220 22664 8340 22692
rect 8481 22695 8539 22701
rect 4982 22584 4988 22636
rect 5040 22584 5046 22636
rect 5353 22627 5411 22633
rect 5353 22593 5365 22627
rect 5399 22593 5411 22627
rect 5353 22587 5411 22593
rect 2682 22516 2688 22568
rect 2740 22516 2746 22568
rect 2961 22559 3019 22565
rect 2961 22525 2973 22559
rect 3007 22556 3019 22559
rect 3510 22556 3516 22568
rect 3007 22528 3516 22556
rect 3007 22525 3019 22528
rect 2961 22519 3019 22525
rect 3510 22516 3516 22528
rect 3568 22516 3574 22568
rect 4433 22559 4491 22565
rect 4433 22525 4445 22559
rect 4479 22556 4491 22559
rect 4706 22556 4712 22568
rect 4479 22528 4712 22556
rect 4479 22525 4491 22528
rect 4433 22519 4491 22525
rect 4706 22516 4712 22528
rect 4764 22556 4770 22568
rect 5368 22556 5396 22587
rect 5810 22584 5816 22636
rect 5868 22584 5874 22636
rect 6733 22627 6791 22633
rect 6733 22593 6745 22627
rect 6779 22624 6791 22627
rect 6822 22624 6828 22636
rect 6779 22596 6828 22624
rect 6779 22593 6791 22596
rect 6733 22587 6791 22593
rect 6822 22584 6828 22596
rect 6880 22584 6886 22636
rect 7009 22627 7067 22633
rect 7009 22593 7021 22627
rect 7055 22593 7067 22627
rect 7009 22587 7067 22593
rect 4764 22528 5396 22556
rect 7024 22556 7052 22587
rect 7098 22584 7104 22636
rect 7156 22584 7162 22636
rect 8220 22633 8248 22664
rect 8481 22661 8493 22695
rect 8527 22661 8539 22695
rect 9858 22692 9864 22704
rect 9706 22664 9864 22692
rect 8481 22655 8539 22661
rect 9858 22652 9864 22664
rect 9916 22652 9922 22704
rect 11238 22652 11244 22704
rect 11296 22692 11302 22704
rect 15286 22692 15292 22704
rect 11296 22664 15292 22692
rect 11296 22652 11302 22664
rect 8205 22627 8263 22633
rect 8205 22593 8217 22627
rect 8251 22593 8263 22627
rect 8205 22587 8263 22593
rect 11146 22584 11152 22636
rect 11204 22584 11210 22636
rect 8478 22556 8484 22568
rect 7024 22528 8484 22556
rect 4764 22516 4770 22528
rect 8478 22516 8484 22528
rect 8536 22516 8542 22568
rect 9766 22516 9772 22568
rect 9824 22556 9830 22568
rect 10045 22559 10103 22565
rect 10045 22556 10057 22559
rect 9824 22528 10057 22556
rect 9824 22516 9830 22528
rect 10045 22525 10057 22528
rect 10091 22525 10103 22559
rect 10045 22519 10103 22525
rect 10318 22516 10324 22568
rect 10376 22556 10382 22568
rect 10597 22559 10655 22565
rect 10597 22556 10609 22559
rect 10376 22528 10609 22556
rect 10376 22516 10382 22528
rect 10597 22525 10609 22528
rect 10643 22525 10655 22559
rect 10597 22519 10655 22525
rect 11974 22516 11980 22568
rect 12032 22516 12038 22568
rect 12161 22559 12219 22565
rect 12161 22525 12173 22559
rect 12207 22556 12219 22559
rect 12360 22556 12388 22664
rect 15286 22652 15292 22664
rect 15344 22652 15350 22704
rect 14645 22627 14703 22633
rect 14645 22593 14657 22627
rect 14691 22624 14703 22627
rect 15562 22624 15568 22636
rect 14691 22596 15568 22624
rect 14691 22593 14703 22596
rect 14645 22587 14703 22593
rect 15562 22584 15568 22596
rect 15620 22584 15626 22636
rect 12207 22528 12388 22556
rect 12207 22525 12219 22528
rect 12161 22519 12219 22525
rect 12434 22516 12440 22568
rect 12492 22556 12498 22568
rect 12897 22559 12955 22565
rect 12897 22556 12909 22559
rect 12492 22528 12909 22556
rect 12492 22516 12498 22528
rect 12897 22525 12909 22528
rect 12943 22525 12955 22559
rect 12897 22519 12955 22525
rect 14734 22516 14740 22568
rect 14792 22516 14798 22568
rect 14921 22559 14979 22565
rect 14921 22525 14933 22559
rect 14967 22556 14979 22559
rect 15010 22556 15016 22568
rect 14967 22528 15016 22556
rect 14967 22525 14979 22528
rect 14921 22519 14979 22525
rect 15010 22516 15016 22528
rect 15068 22516 15074 22568
rect 16022 22516 16028 22568
rect 16080 22516 16086 22568
rect 16408 22488 16436 22720
rect 19242 22692 19248 22704
rect 19076 22664 19248 22692
rect 19076 22633 19104 22664
rect 19242 22652 19248 22664
rect 19300 22652 19306 22704
rect 19352 22701 19380 22732
rect 20806 22720 20812 22772
rect 20864 22760 20870 22772
rect 21450 22760 21456 22772
rect 20864 22732 21456 22760
rect 20864 22720 20870 22732
rect 21450 22720 21456 22732
rect 21508 22720 21514 22772
rect 23382 22760 23388 22772
rect 22296 22732 23388 22760
rect 19337 22695 19395 22701
rect 19337 22661 19349 22695
rect 19383 22661 19395 22695
rect 19337 22655 19395 22661
rect 19061 22627 19119 22633
rect 19061 22593 19073 22627
rect 19107 22593 19119 22627
rect 21266 22624 21272 22636
rect 20470 22596 21272 22624
rect 19061 22587 19119 22593
rect 21266 22584 21272 22596
rect 21324 22584 21330 22636
rect 21468 22633 21496 22720
rect 22186 22692 22192 22704
rect 22020 22664 22192 22692
rect 22020 22633 22048 22664
rect 22186 22652 22192 22664
rect 22244 22652 22250 22704
rect 21453 22627 21511 22633
rect 21453 22593 21465 22627
rect 21499 22593 21511 22627
rect 21453 22587 21511 22593
rect 22005 22627 22063 22633
rect 22005 22593 22017 22627
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 22094 22584 22100 22636
rect 22152 22624 22158 22636
rect 22296 22633 22324 22732
rect 23382 22720 23388 22732
rect 23440 22720 23446 22772
rect 22462 22652 22468 22704
rect 22520 22692 22526 22704
rect 22520 22664 23046 22692
rect 22520 22652 22526 22664
rect 22281 22627 22339 22633
rect 22281 22624 22293 22627
rect 22152 22596 22293 22624
rect 22152 22584 22158 22596
rect 22281 22593 22293 22596
rect 22327 22593 22339 22627
rect 22281 22587 22339 22593
rect 22557 22559 22615 22565
rect 22557 22556 22569 22559
rect 22204 22528 22569 22556
rect 22204 22497 22232 22528
rect 22557 22525 22569 22528
rect 22603 22525 22615 22559
rect 22557 22519 22615 22525
rect 9508 22460 16436 22488
rect 22189 22491 22247 22497
rect 5902 22380 5908 22432
rect 5960 22420 5966 22432
rect 6270 22420 6276 22432
rect 5960 22392 6276 22420
rect 5960 22380 5966 22392
rect 6270 22380 6276 22392
rect 6328 22420 6334 22432
rect 9508 22420 9536 22460
rect 22189 22457 22201 22491
rect 22235 22457 22247 22491
rect 22189 22451 22247 22457
rect 6328 22392 9536 22420
rect 6328 22380 6334 22392
rect 9950 22380 9956 22432
rect 10008 22380 10014 22432
rect 10962 22380 10968 22432
rect 11020 22380 11026 22432
rect 12342 22380 12348 22432
rect 12400 22380 12406 22432
rect 13998 22380 14004 22432
rect 14056 22420 14062 22432
rect 14277 22423 14335 22429
rect 14277 22420 14289 22423
rect 14056 22392 14289 22420
rect 14056 22380 14062 22392
rect 14277 22389 14289 22392
rect 14323 22389 14335 22423
rect 14277 22383 14335 22389
rect 15470 22380 15476 22432
rect 15528 22380 15534 22432
rect 15838 22380 15844 22432
rect 15896 22420 15902 22432
rect 16298 22420 16304 22432
rect 15896 22392 16304 22420
rect 15896 22380 15902 22392
rect 16298 22380 16304 22392
rect 16356 22380 16362 22432
rect 20898 22380 20904 22432
rect 20956 22380 20962 22432
rect 22554 22380 22560 22432
rect 22612 22420 22618 22432
rect 24029 22423 24087 22429
rect 24029 22420 24041 22423
rect 22612 22392 24041 22420
rect 22612 22380 22618 22392
rect 24029 22389 24041 22392
rect 24075 22389 24087 22423
rect 24029 22383 24087 22389
rect 1104 22330 26312 22352
rect 1104 22278 4101 22330
rect 4153 22278 4165 22330
rect 4217 22278 4229 22330
rect 4281 22278 4293 22330
rect 4345 22278 4357 22330
rect 4409 22278 10403 22330
rect 10455 22278 10467 22330
rect 10519 22278 10531 22330
rect 10583 22278 10595 22330
rect 10647 22278 10659 22330
rect 10711 22278 16705 22330
rect 16757 22278 16769 22330
rect 16821 22278 16833 22330
rect 16885 22278 16897 22330
rect 16949 22278 16961 22330
rect 17013 22278 23007 22330
rect 23059 22278 23071 22330
rect 23123 22278 23135 22330
rect 23187 22278 23199 22330
rect 23251 22278 23263 22330
rect 23315 22278 26312 22330
rect 1104 22256 26312 22278
rect 6914 22176 6920 22228
rect 6972 22216 6978 22228
rect 7650 22216 7656 22228
rect 6972 22188 7656 22216
rect 6972 22176 6978 22188
rect 7650 22176 7656 22188
rect 7708 22176 7714 22228
rect 9582 22176 9588 22228
rect 9640 22176 9646 22228
rect 12986 22216 12992 22228
rect 10152 22188 12992 22216
rect 9600 22148 9628 22176
rect 9600 22120 9674 22148
rect 6822 22040 6828 22092
rect 6880 22080 6886 22092
rect 9646 22080 9674 22120
rect 9769 22083 9827 22089
rect 9769 22080 9781 22083
rect 6880 22052 9260 22080
rect 9646 22052 9781 22080
rect 6880 22040 6886 22052
rect 5534 21972 5540 22024
rect 5592 21972 5598 22024
rect 6914 21972 6920 22024
rect 6972 21972 6978 22024
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 21981 9183 22015
rect 9232 22012 9260 22052
rect 9769 22049 9781 22052
rect 9815 22049 9827 22083
rect 10152 22080 10180 22188
rect 12986 22176 12992 22188
rect 13044 22216 13050 22228
rect 14826 22216 14832 22228
rect 13044 22188 14832 22216
rect 13044 22176 13050 22188
rect 14826 22176 14832 22188
rect 14884 22176 14890 22228
rect 15470 22216 15476 22228
rect 15212 22188 15476 22216
rect 14737 22151 14795 22157
rect 14737 22148 14749 22151
rect 14108 22120 14749 22148
rect 9769 22043 9827 22049
rect 9968 22052 10180 22080
rect 9968 22012 9996 22052
rect 10226 22040 10232 22092
rect 10284 22080 10290 22092
rect 10689 22083 10747 22089
rect 10689 22080 10701 22083
rect 10284 22052 10701 22080
rect 10284 22040 10290 22052
rect 10689 22049 10701 22052
rect 10735 22080 10747 22083
rect 13170 22080 13176 22092
rect 10735 22052 13176 22080
rect 10735 22049 10747 22052
rect 10689 22043 10747 22049
rect 13170 22040 13176 22052
rect 13228 22080 13234 22092
rect 13265 22083 13323 22089
rect 13265 22080 13277 22083
rect 13228 22052 13277 22080
rect 13228 22040 13234 22052
rect 13265 22049 13277 22052
rect 13311 22049 13323 22083
rect 13265 22043 13323 22049
rect 9232 21984 9996 22012
rect 9125 21975 9183 21981
rect 5810 21904 5816 21956
rect 5868 21904 5874 21956
rect 7285 21879 7343 21885
rect 7285 21845 7297 21879
rect 7331 21876 7343 21879
rect 8018 21876 8024 21888
rect 7331 21848 8024 21876
rect 7331 21845 7343 21848
rect 7285 21839 7343 21845
rect 8018 21836 8024 21848
rect 8076 21836 8082 21888
rect 8570 21836 8576 21888
rect 8628 21876 8634 21888
rect 8941 21879 8999 21885
rect 8941 21876 8953 21879
rect 8628 21848 8953 21876
rect 8628 21836 8634 21848
rect 8941 21845 8953 21848
rect 8987 21845 8999 21879
rect 9140 21876 9168 21975
rect 10042 21972 10048 22024
rect 10100 21972 10106 22024
rect 10413 22015 10471 22021
rect 10413 21981 10425 22015
rect 10459 22012 10471 22015
rect 10594 22012 10600 22024
rect 10459 21984 10600 22012
rect 10459 21981 10471 21984
rect 10413 21975 10471 21981
rect 10594 21972 10600 21984
rect 10652 21972 10658 22024
rect 12066 21972 12072 22024
rect 12124 21972 12130 22024
rect 13725 22015 13783 22021
rect 13725 21981 13737 22015
rect 13771 22012 13783 22015
rect 14108 22012 14136 22120
rect 14737 22117 14749 22120
rect 14783 22117 14795 22151
rect 14737 22111 14795 22117
rect 14844 22080 14872 22176
rect 15212 22089 15240 22188
rect 15470 22176 15476 22188
rect 15528 22176 15534 22228
rect 16114 22176 16120 22228
rect 16172 22216 16178 22228
rect 17862 22216 17868 22228
rect 16172 22188 17868 22216
rect 16172 22176 16178 22188
rect 17862 22176 17868 22188
rect 17920 22176 17926 22228
rect 22186 22176 22192 22228
rect 22244 22216 22250 22228
rect 22465 22219 22523 22225
rect 22465 22216 22477 22219
rect 22244 22188 22477 22216
rect 22244 22176 22250 22188
rect 22465 22185 22477 22188
rect 22511 22185 22523 22219
rect 22465 22179 22523 22185
rect 16132 22148 16160 22176
rect 15396 22120 16160 22148
rect 15396 22089 15424 22120
rect 22370 22108 22376 22160
rect 22428 22108 22434 22160
rect 14660 22052 14872 22080
rect 15197 22083 15255 22089
rect 14660 22021 14688 22052
rect 15197 22049 15209 22083
rect 15243 22049 15255 22083
rect 15197 22043 15255 22049
rect 15381 22083 15439 22089
rect 15381 22049 15393 22083
rect 15427 22049 15439 22083
rect 15381 22043 15439 22049
rect 15562 22040 15568 22092
rect 15620 22040 15626 22092
rect 17221 22083 17279 22089
rect 17221 22049 17233 22083
rect 17267 22080 17279 22083
rect 18506 22080 18512 22092
rect 17267 22052 18512 22080
rect 17267 22049 17279 22052
rect 17221 22043 17279 22049
rect 18506 22040 18512 22052
rect 18564 22040 18570 22092
rect 19242 22040 19248 22092
rect 19300 22080 19306 22092
rect 19337 22083 19395 22089
rect 19337 22080 19349 22083
rect 19300 22052 19349 22080
rect 19300 22040 19306 22052
rect 19337 22049 19349 22052
rect 19383 22049 19395 22083
rect 19337 22043 19395 22049
rect 20272 22052 21128 22080
rect 13771 21984 14136 22012
rect 14277 22015 14335 22021
rect 13771 21981 13783 21984
rect 13725 21975 13783 21981
rect 14277 21981 14289 22015
rect 14323 22012 14335 22015
rect 14645 22015 14703 22021
rect 14323 21984 14596 22012
rect 14323 21981 14335 21984
rect 14277 21975 14335 21981
rect 9677 21947 9735 21953
rect 9677 21913 9689 21947
rect 9723 21944 9735 21947
rect 9766 21944 9772 21956
rect 9723 21916 9772 21944
rect 9723 21913 9735 21916
rect 9677 21907 9735 21913
rect 9766 21904 9772 21916
rect 9824 21904 9830 21956
rect 10226 21904 10232 21956
rect 10284 21904 10290 21956
rect 10318 21904 10324 21956
rect 10376 21904 10382 21956
rect 10520 21916 10824 21944
rect 9217 21879 9275 21885
rect 9217 21876 9229 21879
rect 9140 21848 9229 21876
rect 8941 21839 8999 21845
rect 9217 21845 9229 21848
rect 9263 21845 9275 21879
rect 9217 21839 9275 21845
rect 9582 21836 9588 21888
rect 9640 21876 9646 21888
rect 9950 21876 9956 21888
rect 9640 21848 9956 21876
rect 9640 21836 9646 21848
rect 9950 21836 9956 21848
rect 10008 21876 10014 21888
rect 10520 21876 10548 21916
rect 10796 21888 10824 21916
rect 10962 21904 10968 21956
rect 11020 21904 11026 21956
rect 12526 21944 12532 21956
rect 12360 21916 12532 21944
rect 10008 21848 10548 21876
rect 10008 21836 10014 21848
rect 10594 21836 10600 21888
rect 10652 21836 10658 21888
rect 10778 21836 10784 21888
rect 10836 21836 10842 21888
rect 11054 21836 11060 21888
rect 11112 21876 11118 21888
rect 12360 21876 12388 21916
rect 12526 21904 12532 21916
rect 12584 21904 12590 21956
rect 14366 21904 14372 21956
rect 14424 21904 14430 21956
rect 14458 21904 14464 21956
rect 14516 21904 14522 21956
rect 14568 21944 14596 21984
rect 14645 21981 14657 22015
rect 14691 21981 14703 22015
rect 14645 21975 14703 21981
rect 14734 21972 14740 22024
rect 14792 22012 14798 22024
rect 15105 22015 15163 22021
rect 15105 22012 15117 22015
rect 14792 21984 15117 22012
rect 14792 21972 14798 21984
rect 15105 21981 15117 21984
rect 15151 21981 15163 22015
rect 15105 21975 15163 21981
rect 16114 21972 16120 22024
rect 16172 21972 16178 22024
rect 16206 21972 16212 22024
rect 16264 21972 16270 22024
rect 16301 22015 16359 22021
rect 16301 21981 16313 22015
rect 16347 21981 16359 22015
rect 16301 21975 16359 21981
rect 15194 21944 15200 21956
rect 14568 21916 15200 21944
rect 15194 21904 15200 21916
rect 15252 21944 15258 21956
rect 16224 21944 16252 21972
rect 15252 21916 16252 21944
rect 16316 21944 16344 21975
rect 17494 21972 17500 22024
rect 17552 22012 17558 22024
rect 17589 22015 17647 22021
rect 17589 22012 17601 22015
rect 17552 21984 17601 22012
rect 17552 21972 17558 21984
rect 17589 21981 17601 21984
rect 17635 21981 17647 22015
rect 17589 21975 17647 21981
rect 18417 22015 18475 22021
rect 18417 21981 18429 22015
rect 18463 22012 18475 22015
rect 18690 22012 18696 22024
rect 18463 21984 18696 22012
rect 18463 21981 18475 21984
rect 18417 21975 18475 21981
rect 18690 21972 18696 21984
rect 18748 21972 18754 22024
rect 20272 22021 20300 22052
rect 20257 22015 20315 22021
rect 20257 21981 20269 22015
rect 20303 21981 20315 22015
rect 20257 21975 20315 21981
rect 20441 22015 20499 22021
rect 20441 21981 20453 22015
rect 20487 22012 20499 22015
rect 20625 22015 20683 22021
rect 20625 22012 20637 22015
rect 20487 21984 20637 22012
rect 20487 21981 20499 21984
rect 20441 21975 20499 21981
rect 20625 21981 20637 21984
rect 20671 21981 20683 22015
rect 20625 21975 20683 21981
rect 20714 21972 20720 22024
rect 20772 21972 20778 22024
rect 21100 22021 21128 22052
rect 22554 22040 22560 22092
rect 22612 22080 22618 22092
rect 22925 22083 22983 22089
rect 22925 22080 22937 22083
rect 22612 22052 22937 22080
rect 22612 22040 22618 22052
rect 22925 22049 22937 22052
rect 22971 22049 22983 22083
rect 22925 22043 22983 22049
rect 23017 22083 23075 22089
rect 23017 22049 23029 22083
rect 23063 22049 23075 22083
rect 23017 22043 23075 22049
rect 21085 22015 21143 22021
rect 21085 21981 21097 22015
rect 21131 22012 21143 22015
rect 21131 21984 21680 22012
rect 21131 21981 21143 21984
rect 21085 21975 21143 21981
rect 16945 21947 17003 21953
rect 16316 21916 16620 21944
rect 15252 21904 15258 21916
rect 11112 21848 12388 21876
rect 11112 21836 11118 21848
rect 12434 21836 12440 21888
rect 12492 21836 12498 21888
rect 13906 21836 13912 21888
rect 13964 21836 13970 21888
rect 14090 21836 14096 21888
rect 14148 21836 14154 21888
rect 16482 21836 16488 21888
rect 16540 21836 16546 21888
rect 16592 21885 16620 21916
rect 16945 21913 16957 21947
rect 16991 21944 17003 21947
rect 17773 21947 17831 21953
rect 17773 21944 17785 21947
rect 16991 21916 17785 21944
rect 16991 21913 17003 21916
rect 16945 21907 17003 21913
rect 17773 21913 17785 21916
rect 17819 21913 17831 21947
rect 17773 21907 17831 21913
rect 19334 21904 19340 21956
rect 19392 21944 19398 21956
rect 20165 21947 20223 21953
rect 20165 21944 20177 21947
rect 19392 21916 20177 21944
rect 19392 21904 19398 21916
rect 20165 21913 20177 21916
rect 20211 21913 20223 21947
rect 20165 21907 20223 21913
rect 21542 21904 21548 21956
rect 21600 21904 21606 21956
rect 21652 21944 21680 21984
rect 21910 21972 21916 22024
rect 21968 21972 21974 22024
rect 23032 22012 23060 22043
rect 22756 21984 23060 22012
rect 22756 21956 22784 21984
rect 22554 21944 22560 21956
rect 21652 21916 22560 21944
rect 22554 21904 22560 21916
rect 22612 21944 22618 21956
rect 22738 21944 22744 21956
rect 22612 21916 22744 21944
rect 22612 21904 22618 21916
rect 22738 21904 22744 21916
rect 22796 21904 22802 21956
rect 16577 21879 16635 21885
rect 16577 21845 16589 21879
rect 16623 21845 16635 21879
rect 16577 21839 16635 21845
rect 17034 21836 17040 21888
rect 17092 21836 17098 21888
rect 17402 21836 17408 21888
rect 17460 21836 17466 21888
rect 20346 21836 20352 21888
rect 20404 21836 20410 21888
rect 22830 21836 22836 21888
rect 22888 21836 22894 21888
rect 1104 21786 26472 21808
rect 1104 21734 7252 21786
rect 7304 21734 7316 21786
rect 7368 21734 7380 21786
rect 7432 21734 7444 21786
rect 7496 21734 7508 21786
rect 7560 21734 13554 21786
rect 13606 21734 13618 21786
rect 13670 21734 13682 21786
rect 13734 21734 13746 21786
rect 13798 21734 13810 21786
rect 13862 21734 19856 21786
rect 19908 21734 19920 21786
rect 19972 21734 19984 21786
rect 20036 21734 20048 21786
rect 20100 21734 20112 21786
rect 20164 21734 26158 21786
rect 26210 21734 26222 21786
rect 26274 21734 26286 21786
rect 26338 21734 26350 21786
rect 26402 21734 26414 21786
rect 26466 21734 26472 21786
rect 1104 21712 26472 21734
rect 5534 21672 5540 21684
rect 2792 21644 5540 21672
rect 2682 21564 2688 21616
rect 2740 21604 2746 21616
rect 2792 21604 2820 21644
rect 5534 21632 5540 21644
rect 5592 21632 5598 21684
rect 10134 21672 10140 21684
rect 6380 21644 10140 21672
rect 2740 21576 2820 21604
rect 2740 21564 2746 21576
rect 1765 21539 1823 21545
rect 1765 21505 1777 21539
rect 1811 21536 1823 21539
rect 1946 21536 1952 21548
rect 1811 21508 1952 21536
rect 1811 21505 1823 21508
rect 1765 21499 1823 21505
rect 1946 21496 1952 21508
rect 2004 21496 2010 21548
rect 2792 21545 2820 21576
rect 3142 21564 3148 21616
rect 3200 21604 3206 21616
rect 3200 21576 3542 21604
rect 3200 21564 3206 21576
rect 2777 21539 2835 21545
rect 2777 21505 2789 21539
rect 2823 21505 2835 21539
rect 5552 21536 5580 21632
rect 6380 21613 6408 21644
rect 10134 21632 10140 21644
rect 10192 21672 10198 21684
rect 11054 21672 11060 21684
rect 10192 21644 11060 21672
rect 10192 21632 10198 21644
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 11146 21632 11152 21684
rect 11204 21672 11210 21684
rect 11517 21675 11575 21681
rect 11517 21672 11529 21675
rect 11204 21644 11529 21672
rect 11204 21632 11210 21644
rect 11517 21641 11529 21644
rect 11563 21641 11575 21675
rect 11517 21635 11575 21641
rect 11885 21675 11943 21681
rect 11885 21641 11897 21675
rect 11931 21672 11943 21675
rect 12342 21672 12348 21684
rect 11931 21644 12348 21672
rect 11931 21641 11943 21644
rect 11885 21635 11943 21641
rect 12342 21632 12348 21644
rect 12400 21632 12406 21684
rect 12434 21632 12440 21684
rect 12492 21672 12498 21684
rect 12492 21644 13676 21672
rect 12492 21632 12498 21644
rect 6365 21607 6423 21613
rect 6365 21573 6377 21607
rect 6411 21573 6423 21607
rect 6365 21567 6423 21573
rect 8570 21564 8576 21616
rect 8628 21564 8634 21616
rect 10042 21564 10048 21616
rect 10100 21564 10106 21616
rect 10594 21564 10600 21616
rect 10652 21604 10658 21616
rect 10652 21576 12434 21604
rect 10652 21564 10658 21576
rect 6270 21536 6276 21548
rect 5552 21508 6276 21536
rect 2777 21499 2835 21505
rect 6270 21496 6276 21508
rect 6328 21536 6334 21548
rect 7101 21539 7159 21545
rect 7101 21536 7113 21539
rect 6328 21508 7113 21536
rect 6328 21496 6334 21508
rect 7101 21505 7113 21508
rect 7147 21536 7159 21539
rect 8294 21536 8300 21548
rect 7147 21508 8300 21536
rect 7147 21505 7159 21508
rect 7101 21499 7159 21505
rect 8294 21496 8300 21508
rect 8352 21496 8358 21548
rect 9582 21496 9588 21548
rect 9640 21496 9646 21548
rect 9858 21536 9864 21548
rect 9706 21508 9864 21536
rect 9858 21496 9864 21508
rect 9916 21496 9922 21548
rect 10060 21536 10088 21564
rect 10689 21539 10747 21545
rect 10689 21536 10701 21539
rect 10060 21508 10701 21536
rect 10689 21505 10701 21508
rect 10735 21505 10747 21539
rect 10689 21499 10747 21505
rect 10778 21496 10784 21548
rect 10836 21536 10842 21548
rect 11974 21536 11980 21548
rect 10836 21508 11980 21536
rect 10836 21496 10842 21508
rect 11974 21496 11980 21508
rect 12032 21496 12038 21548
rect 12406 21536 12434 21576
rect 12802 21564 12808 21616
rect 12860 21604 12866 21616
rect 12860 21576 13492 21604
rect 12860 21564 12866 21576
rect 13265 21539 13323 21545
rect 13265 21536 13277 21539
rect 12406 21508 13277 21536
rect 13265 21505 13277 21508
rect 13311 21505 13323 21539
rect 13265 21499 13323 21505
rect 13354 21496 13360 21548
rect 13412 21496 13418 21548
rect 13464 21536 13492 21576
rect 13538 21564 13544 21616
rect 13596 21564 13602 21616
rect 13648 21613 13676 21644
rect 14366 21632 14372 21684
rect 14424 21672 14430 21684
rect 15841 21675 15899 21681
rect 15841 21672 15853 21675
rect 14424 21644 15853 21672
rect 14424 21632 14430 21644
rect 15841 21641 15853 21644
rect 15887 21641 15899 21675
rect 15841 21635 15899 21641
rect 16206 21632 16212 21684
rect 16264 21672 16270 21684
rect 20346 21672 20352 21684
rect 16264 21644 18552 21672
rect 16264 21632 16270 21644
rect 13633 21607 13691 21613
rect 13633 21573 13645 21607
rect 13679 21573 13691 21607
rect 13633 21567 13691 21573
rect 13906 21564 13912 21616
rect 13964 21604 13970 21616
rect 14277 21607 14335 21613
rect 14277 21604 14289 21607
rect 13964 21576 14289 21604
rect 13964 21564 13970 21576
rect 14277 21573 14289 21576
rect 14323 21573 14335 21607
rect 14277 21567 14335 21573
rect 14918 21564 14924 21616
rect 14976 21564 14982 21616
rect 16482 21564 16488 21616
rect 16540 21604 16546 21616
rect 16945 21607 17003 21613
rect 16945 21604 16957 21607
rect 16540 21576 16957 21604
rect 16540 21564 16546 21576
rect 16945 21573 16957 21576
rect 16991 21573 17003 21607
rect 16945 21567 17003 21573
rect 17954 21564 17960 21616
rect 18012 21564 18018 21616
rect 13730 21539 13788 21545
rect 13730 21536 13742 21539
rect 13464 21508 13742 21536
rect 13730 21505 13742 21508
rect 13776 21505 13788 21539
rect 16393 21539 16451 21545
rect 16393 21536 16405 21539
rect 13730 21499 13788 21505
rect 15672 21508 16405 21536
rect 3050 21428 3056 21480
rect 3108 21428 3114 21480
rect 4798 21428 4804 21480
rect 4856 21468 4862 21480
rect 6362 21468 6368 21480
rect 4856 21440 6368 21468
rect 4856 21428 4862 21440
rect 6362 21428 6368 21440
rect 6420 21468 6426 21480
rect 7466 21468 7472 21480
rect 6420 21440 7472 21468
rect 6420 21428 6426 21440
rect 7466 21428 7472 21440
rect 7524 21428 7530 21480
rect 8018 21428 8024 21480
rect 8076 21468 8082 21480
rect 9600 21468 9628 21496
rect 8076 21440 9628 21468
rect 10045 21471 10103 21477
rect 8076 21428 8082 21440
rect 10045 21437 10057 21471
rect 10091 21468 10103 21471
rect 10318 21468 10324 21480
rect 10091 21440 10324 21468
rect 10091 21437 10103 21440
rect 10045 21431 10103 21437
rect 10318 21428 10324 21440
rect 10376 21428 10382 21480
rect 11422 21428 11428 21480
rect 11480 21468 11486 21480
rect 12066 21468 12072 21480
rect 11480 21440 12072 21468
rect 11480 21428 11486 21440
rect 12066 21428 12072 21440
rect 12124 21428 12130 21480
rect 12161 21471 12219 21477
rect 12161 21437 12173 21471
rect 12207 21468 12219 21471
rect 12250 21468 12256 21480
rect 12207 21440 12256 21468
rect 12207 21437 12219 21440
rect 12161 21431 12219 21437
rect 12250 21428 12256 21440
rect 12308 21428 12314 21480
rect 12802 21428 12808 21480
rect 12860 21468 12866 21480
rect 13081 21471 13139 21477
rect 13081 21468 13093 21471
rect 12860 21440 13093 21468
rect 12860 21428 12866 21440
rect 13081 21437 13093 21440
rect 13127 21437 13139 21471
rect 13081 21431 13139 21437
rect 13170 21428 13176 21480
rect 13228 21468 13234 21480
rect 14001 21471 14059 21477
rect 14001 21468 14013 21471
rect 13228 21440 14013 21468
rect 13228 21428 13234 21440
rect 14001 21437 14013 21440
rect 14047 21437 14059 21471
rect 14001 21431 14059 21437
rect 14734 21428 14740 21480
rect 14792 21468 14798 21480
rect 15672 21468 15700 21508
rect 16393 21505 16405 21508
rect 16439 21505 16451 21539
rect 16393 21499 16451 21505
rect 14792 21440 15700 21468
rect 15749 21471 15807 21477
rect 14792 21428 14798 21440
rect 15749 21437 15761 21471
rect 15795 21468 15807 21471
rect 16022 21468 16028 21480
rect 15795 21440 16028 21468
rect 15795 21437 15807 21440
rect 15749 21431 15807 21437
rect 16022 21428 16028 21440
rect 16080 21428 16086 21480
rect 16408 21468 16436 21499
rect 16574 21496 16580 21548
rect 16632 21536 16638 21548
rect 16669 21539 16727 21545
rect 16669 21536 16681 21539
rect 16632 21508 16681 21536
rect 16632 21496 16638 21508
rect 16669 21505 16681 21508
rect 16715 21505 16727 21539
rect 16669 21499 16727 21505
rect 17034 21468 17040 21480
rect 16408 21440 17040 21468
rect 17034 21428 17040 21440
rect 17092 21428 17098 21480
rect 18524 21468 18552 21644
rect 19720 21644 20352 21672
rect 19720 21613 19748 21644
rect 20346 21632 20352 21644
rect 20404 21632 20410 21684
rect 22830 21632 22836 21684
rect 22888 21672 22894 21684
rect 23201 21675 23259 21681
rect 23201 21672 23213 21675
rect 22888 21644 23213 21672
rect 22888 21632 22894 21644
rect 23201 21641 23213 21644
rect 23247 21641 23259 21675
rect 23201 21635 23259 21641
rect 19705 21607 19763 21613
rect 19705 21573 19717 21607
rect 19751 21573 19763 21607
rect 19705 21567 19763 21573
rect 20990 21564 20996 21616
rect 21048 21604 21054 21616
rect 22281 21607 22339 21613
rect 22281 21604 22293 21607
rect 21048 21576 22293 21604
rect 21048 21564 21054 21576
rect 22281 21573 22293 21576
rect 22327 21573 22339 21607
rect 22281 21567 22339 21573
rect 19242 21496 19248 21548
rect 19300 21536 19306 21548
rect 19429 21539 19487 21545
rect 19429 21536 19441 21539
rect 19300 21508 19441 21536
rect 19300 21496 19306 21508
rect 19429 21505 19441 21508
rect 19475 21505 19487 21539
rect 21266 21536 21272 21548
rect 20838 21508 21272 21536
rect 19429 21499 19487 21505
rect 21266 21496 21272 21508
rect 21324 21496 21330 21548
rect 21913 21539 21971 21545
rect 21913 21505 21925 21539
rect 21959 21505 21971 21539
rect 21913 21499 21971 21505
rect 20898 21468 20904 21480
rect 18524 21440 20904 21468
rect 20898 21428 20904 21440
rect 20956 21428 20962 21480
rect 21177 21471 21235 21477
rect 21177 21437 21189 21471
rect 21223 21468 21235 21471
rect 21928 21468 21956 21499
rect 22646 21496 22652 21548
rect 22704 21536 22710 21548
rect 23382 21536 23388 21548
rect 22704 21508 23388 21536
rect 22704 21496 22710 21508
rect 23382 21496 23388 21508
rect 23440 21536 23446 21548
rect 23753 21539 23811 21545
rect 23753 21536 23765 21539
rect 23440 21508 23765 21536
rect 23440 21496 23446 21508
rect 23753 21505 23765 21508
rect 23799 21505 23811 21539
rect 23753 21499 23811 21505
rect 25682 21496 25688 21548
rect 25740 21496 25746 21548
rect 21223 21440 21956 21468
rect 21223 21437 21235 21440
rect 21177 21431 21235 21437
rect 934 21292 940 21344
rect 992 21332 998 21344
rect 1489 21335 1547 21341
rect 1489 21332 1501 21335
rect 992 21304 1501 21332
rect 992 21292 998 21304
rect 1489 21301 1501 21304
rect 1535 21301 1547 21335
rect 1489 21295 1547 21301
rect 5994 21292 6000 21344
rect 6052 21332 6058 21344
rect 7282 21332 7288 21344
rect 6052 21304 7288 21332
rect 6052 21292 6058 21304
rect 7282 21292 7288 21304
rect 7340 21292 7346 21344
rect 7374 21292 7380 21344
rect 7432 21292 7438 21344
rect 10134 21292 10140 21344
rect 10192 21292 10198 21344
rect 12434 21292 12440 21344
rect 12492 21332 12498 21344
rect 12529 21335 12587 21341
rect 12529 21332 12541 21335
rect 12492 21304 12541 21332
rect 12492 21292 12498 21304
rect 12529 21301 12541 21304
rect 12575 21301 12587 21335
rect 12529 21295 12587 21301
rect 13906 21292 13912 21344
rect 13964 21292 13970 21344
rect 18417 21335 18475 21341
rect 18417 21301 18429 21335
rect 18463 21332 18475 21335
rect 18690 21332 18696 21344
rect 18463 21304 18696 21332
rect 18463 21301 18475 21304
rect 18417 21295 18475 21301
rect 18690 21292 18696 21304
rect 18748 21292 18754 21344
rect 25866 21292 25872 21344
rect 25924 21292 25930 21344
rect 1104 21242 26312 21264
rect 1104 21190 4101 21242
rect 4153 21190 4165 21242
rect 4217 21190 4229 21242
rect 4281 21190 4293 21242
rect 4345 21190 4357 21242
rect 4409 21190 10403 21242
rect 10455 21190 10467 21242
rect 10519 21190 10531 21242
rect 10583 21190 10595 21242
rect 10647 21190 10659 21242
rect 10711 21190 16705 21242
rect 16757 21190 16769 21242
rect 16821 21190 16833 21242
rect 16885 21190 16897 21242
rect 16949 21190 16961 21242
rect 17013 21190 23007 21242
rect 23059 21190 23071 21242
rect 23123 21190 23135 21242
rect 23187 21190 23199 21242
rect 23251 21190 23263 21242
rect 23315 21190 26312 21242
rect 1104 21168 26312 21190
rect 3050 21088 3056 21140
rect 3108 21128 3114 21140
rect 3145 21131 3203 21137
rect 3145 21128 3157 21131
rect 3108 21100 3157 21128
rect 3108 21088 3114 21100
rect 3145 21097 3157 21100
rect 3191 21097 3203 21131
rect 3145 21091 3203 21097
rect 5810 21088 5816 21140
rect 5868 21088 5874 21140
rect 6181 21131 6239 21137
rect 6181 21097 6193 21131
rect 6227 21128 6239 21131
rect 6546 21128 6552 21140
rect 6227 21100 6552 21128
rect 6227 21097 6239 21100
rect 6181 21091 6239 21097
rect 6546 21088 6552 21100
rect 6604 21088 6610 21140
rect 6730 21088 6736 21140
rect 6788 21128 6794 21140
rect 9125 21131 9183 21137
rect 6788 21100 7236 21128
rect 6788 21088 6794 21100
rect 5828 21060 5856 21088
rect 6365 21063 6423 21069
rect 6365 21060 6377 21063
rect 5828 21032 6377 21060
rect 6365 21029 6377 21032
rect 6411 21029 6423 21063
rect 7101 21063 7159 21069
rect 7101 21060 7113 21063
rect 6365 21023 6423 21029
rect 6564 21032 7113 21060
rect 4154 20952 4160 21004
rect 4212 20992 4218 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 4212 20964 4445 20992
rect 4212 20952 4218 20964
rect 4433 20961 4445 20964
rect 4479 20992 4491 20995
rect 5258 20992 5264 21004
rect 4479 20964 5264 20992
rect 4479 20961 4491 20964
rect 4433 20955 4491 20961
rect 5258 20952 5264 20964
rect 5316 20952 5322 21004
rect 5828 20964 6224 20992
rect 3329 20927 3387 20933
rect 3329 20893 3341 20927
rect 3375 20924 3387 20927
rect 3375 20896 3832 20924
rect 3375 20893 3387 20896
rect 3329 20887 3387 20893
rect 3804 20797 3832 20896
rect 4798 20884 4804 20936
rect 4856 20884 4862 20936
rect 5828 20933 5856 20964
rect 6196 20936 6224 20964
rect 5537 20927 5595 20933
rect 5537 20924 5549 20927
rect 4908 20896 5549 20924
rect 4157 20859 4215 20865
rect 4157 20825 4169 20859
rect 4203 20856 4215 20859
rect 4816 20856 4844 20884
rect 4203 20828 4844 20856
rect 4203 20825 4215 20828
rect 4157 20819 4215 20825
rect 3789 20791 3847 20797
rect 3789 20757 3801 20791
rect 3835 20757 3847 20791
rect 3789 20751 3847 20757
rect 4249 20791 4307 20797
rect 4249 20757 4261 20791
rect 4295 20788 4307 20791
rect 4798 20788 4804 20800
rect 4295 20760 4804 20788
rect 4295 20757 4307 20760
rect 4249 20751 4307 20757
rect 4798 20748 4804 20760
rect 4856 20788 4862 20800
rect 4908 20788 4936 20896
rect 5537 20893 5549 20896
rect 5583 20893 5595 20927
rect 5537 20887 5595 20893
rect 5813 20927 5871 20933
rect 5813 20893 5825 20927
rect 5859 20893 5871 20927
rect 5813 20887 5871 20893
rect 5997 20927 6055 20933
rect 5997 20893 6009 20927
rect 6043 20893 6055 20927
rect 5997 20887 6055 20893
rect 5258 20816 5264 20868
rect 5316 20856 5322 20868
rect 5675 20859 5733 20865
rect 5675 20856 5687 20859
rect 5316 20828 5687 20856
rect 5316 20816 5322 20828
rect 5675 20825 5687 20828
rect 5721 20825 5733 20859
rect 5675 20819 5733 20825
rect 5905 20859 5963 20865
rect 5905 20825 5917 20859
rect 5951 20825 5963 20859
rect 6012 20856 6040 20887
rect 6178 20884 6184 20936
rect 6236 20884 6242 20936
rect 6564 20933 6592 21032
rect 7101 21029 7113 21032
rect 7147 21029 7159 21063
rect 7208 21060 7236 21100
rect 9125 21097 9137 21131
rect 9171 21128 9183 21131
rect 9306 21128 9312 21140
rect 9171 21100 9312 21128
rect 9171 21097 9183 21100
rect 9125 21091 9183 21097
rect 9306 21088 9312 21100
rect 9364 21088 9370 21140
rect 10134 21088 10140 21140
rect 10192 21088 10198 21140
rect 15102 21128 15108 21140
rect 12406 21100 15108 21128
rect 7653 21063 7711 21069
rect 7653 21060 7665 21063
rect 7208 21032 7665 21060
rect 7101 21023 7159 21029
rect 7653 21029 7665 21032
rect 7699 21029 7711 21063
rect 7653 21023 7711 21029
rect 6638 20952 6644 21004
rect 6696 20952 6702 21004
rect 7374 20992 7380 21004
rect 6886 20964 7380 20992
rect 6549 20927 6607 20933
rect 6549 20893 6561 20927
rect 6595 20893 6607 20927
rect 6656 20924 6684 20952
rect 6886 20933 6914 20964
rect 7374 20952 7380 20964
rect 7432 20952 7438 21004
rect 7837 20995 7895 21001
rect 7837 20992 7849 20995
rect 7668 20964 7849 20992
rect 6733 20927 6791 20933
rect 6733 20924 6745 20927
rect 6656 20896 6745 20924
rect 6549 20887 6607 20893
rect 6733 20893 6745 20896
rect 6779 20893 6791 20927
rect 6733 20887 6791 20893
rect 6871 20927 6929 20933
rect 6871 20893 6883 20927
rect 6917 20893 6929 20927
rect 6871 20887 6929 20893
rect 7009 20927 7067 20933
rect 7009 20893 7021 20927
rect 7055 20893 7067 20927
rect 7009 20887 7067 20893
rect 6641 20859 6699 20865
rect 6012 20828 6592 20856
rect 5905 20819 5963 20825
rect 4856 20760 4936 20788
rect 5920 20788 5948 20819
rect 6564 20800 6592 20828
rect 6641 20825 6653 20859
rect 6687 20825 6699 20859
rect 7024 20856 7052 20887
rect 7098 20884 7104 20936
rect 7156 20924 7162 20936
rect 7561 20927 7619 20933
rect 7561 20924 7573 20927
rect 7156 20896 7573 20924
rect 7156 20884 7162 20896
rect 7561 20893 7573 20896
rect 7607 20893 7619 20927
rect 7561 20887 7619 20893
rect 7190 20856 7196 20868
rect 7024 20828 7196 20856
rect 6641 20819 6699 20825
rect 6178 20788 6184 20800
rect 5920 20760 6184 20788
rect 4856 20748 4862 20760
rect 6178 20748 6184 20760
rect 6236 20748 6242 20800
rect 6546 20748 6552 20800
rect 6604 20748 6610 20800
rect 6656 20788 6684 20819
rect 7190 20816 7196 20828
rect 7248 20816 7254 20868
rect 7282 20816 7288 20868
rect 7340 20816 7346 20868
rect 7466 20816 7472 20868
rect 7524 20856 7530 20868
rect 7668 20856 7696 20964
rect 7837 20961 7849 20964
rect 7883 20961 7895 20995
rect 7837 20955 7895 20961
rect 9398 20952 9404 21004
rect 9456 20992 9462 21004
rect 9677 20995 9735 21001
rect 9677 20992 9689 20995
rect 9456 20964 9689 20992
rect 9456 20952 9462 20964
rect 9677 20961 9689 20964
rect 9723 20961 9735 20995
rect 9677 20955 9735 20961
rect 9493 20927 9551 20933
rect 9493 20893 9505 20927
rect 9539 20924 9551 20927
rect 10152 20924 10180 21088
rect 9539 20896 10180 20924
rect 9539 20893 9551 20896
rect 9493 20887 9551 20893
rect 7524 20828 7696 20856
rect 7524 20816 7530 20828
rect 8110 20816 8116 20868
rect 8168 20856 8174 20868
rect 12406 20856 12434 21100
rect 15102 21088 15108 21100
rect 15160 21088 15166 21140
rect 15841 21131 15899 21137
rect 15841 21097 15853 21131
rect 15887 21128 15899 21131
rect 16114 21128 16120 21140
rect 15887 21100 16120 21128
rect 15887 21097 15899 21100
rect 15841 21091 15899 21097
rect 16114 21088 16120 21100
rect 16172 21088 16178 21140
rect 16390 21088 16396 21140
rect 16448 21128 16454 21140
rect 20990 21128 20996 21140
rect 16448 21100 20996 21128
rect 16448 21088 16454 21100
rect 20990 21088 20996 21100
rect 21048 21088 21054 21140
rect 21637 21131 21695 21137
rect 21637 21097 21649 21131
rect 21683 21128 21695 21131
rect 21986 21131 22044 21137
rect 21986 21128 21998 21131
rect 21683 21100 21998 21128
rect 21683 21097 21695 21100
rect 21637 21091 21695 21097
rect 21986 21097 21998 21100
rect 22032 21097 22044 21131
rect 21986 21091 22044 21097
rect 23382 21088 23388 21140
rect 23440 21128 23446 21140
rect 23477 21131 23535 21137
rect 23477 21128 23489 21131
rect 23440 21100 23489 21128
rect 23440 21088 23446 21100
rect 23477 21097 23489 21100
rect 23523 21097 23535 21131
rect 23477 21091 23535 21097
rect 17954 21020 17960 21072
rect 18012 21020 18018 21072
rect 16390 20992 16396 21004
rect 12544 20964 16396 20992
rect 12544 20936 12572 20964
rect 16390 20952 16396 20964
rect 16448 20952 16454 21004
rect 16482 20952 16488 21004
rect 16540 20952 16546 21004
rect 16761 20995 16819 21001
rect 16761 20961 16773 20995
rect 16807 20992 16819 20995
rect 17402 20992 17408 21004
rect 16807 20964 17408 20992
rect 16807 20961 16819 20964
rect 16761 20955 16819 20961
rect 17402 20952 17408 20964
rect 17460 20952 17466 21004
rect 12526 20884 12532 20936
rect 12584 20884 12590 20936
rect 13725 20927 13783 20933
rect 13725 20893 13737 20927
rect 13771 20924 13783 20927
rect 13998 20924 14004 20936
rect 13771 20896 14004 20924
rect 13771 20893 13783 20896
rect 13725 20887 13783 20893
rect 13998 20884 14004 20896
rect 14056 20884 14062 20936
rect 14093 20927 14151 20933
rect 14093 20893 14105 20927
rect 14139 20893 14151 20927
rect 14093 20887 14151 20893
rect 8168 20828 12434 20856
rect 8168 20816 8174 20828
rect 13078 20816 13084 20868
rect 13136 20856 13142 20868
rect 13265 20859 13323 20865
rect 13265 20856 13277 20859
rect 13136 20828 13277 20856
rect 13136 20816 13142 20828
rect 13265 20825 13277 20828
rect 13311 20856 13323 20859
rect 14108 20856 14136 20887
rect 17770 20884 17776 20936
rect 17828 20924 17834 20936
rect 17972 20924 18000 21020
rect 18233 20995 18291 21001
rect 18233 20961 18245 20995
rect 18279 20992 18291 20995
rect 18877 20995 18935 21001
rect 18877 20992 18889 20995
rect 18279 20964 18889 20992
rect 18279 20961 18291 20964
rect 18233 20955 18291 20961
rect 18877 20961 18889 20964
rect 18923 20992 18935 20995
rect 18966 20992 18972 21004
rect 18923 20964 18972 20992
rect 18923 20961 18935 20964
rect 18877 20955 18935 20961
rect 18966 20952 18972 20964
rect 19024 20952 19030 21004
rect 19521 20995 19579 21001
rect 19521 20961 19533 20995
rect 19567 20992 19579 20995
rect 21082 20992 21088 21004
rect 19567 20964 21088 20992
rect 19567 20961 19579 20964
rect 19521 20955 19579 20961
rect 21082 20952 21088 20964
rect 21140 20952 21146 21004
rect 21729 20995 21787 21001
rect 21729 20961 21741 20995
rect 21775 20992 21787 20995
rect 22094 20992 22100 21004
rect 21775 20964 22100 20992
rect 21775 20961 21787 20964
rect 21729 20955 21787 20961
rect 22094 20952 22100 20964
rect 22152 20952 22158 21004
rect 17828 20896 18000 20924
rect 17828 20884 17834 20896
rect 18414 20884 18420 20936
rect 18472 20924 18478 20936
rect 19245 20927 19303 20933
rect 19245 20924 19257 20927
rect 18472 20896 19257 20924
rect 18472 20884 18478 20896
rect 19245 20893 19257 20896
rect 19291 20893 19303 20927
rect 19245 20887 19303 20893
rect 21450 20884 21456 20936
rect 21508 20884 21514 20936
rect 13311 20828 14136 20856
rect 14369 20859 14427 20865
rect 13311 20825 13323 20828
rect 13265 20819 13323 20825
rect 14369 20825 14381 20859
rect 14415 20825 14427 20859
rect 15838 20856 15844 20868
rect 15594 20828 15844 20856
rect 14369 20819 14427 20825
rect 7837 20791 7895 20797
rect 7837 20788 7849 20791
rect 6656 20760 7849 20788
rect 7837 20757 7849 20760
rect 7883 20757 7895 20791
rect 7837 20751 7895 20757
rect 9585 20791 9643 20797
rect 9585 20757 9597 20791
rect 9631 20788 9643 20791
rect 9950 20788 9956 20800
rect 9631 20760 9956 20788
rect 9631 20757 9643 20760
rect 9585 20751 9643 20757
rect 9950 20748 9956 20760
rect 10008 20748 10014 20800
rect 13909 20791 13967 20797
rect 13909 20757 13921 20791
rect 13955 20788 13967 20791
rect 14384 20788 14412 20819
rect 13955 20760 14412 20788
rect 13955 20757 13967 20760
rect 13909 20751 13967 20757
rect 14550 20748 14556 20800
rect 14608 20788 14614 20800
rect 15672 20788 15700 20828
rect 15838 20816 15844 20828
rect 15896 20816 15902 20868
rect 18046 20816 18052 20868
rect 18104 20856 18110 20868
rect 18325 20859 18383 20865
rect 18325 20856 18337 20859
rect 18104 20828 18337 20856
rect 18104 20816 18110 20828
rect 18325 20825 18337 20828
rect 18371 20825 18383 20859
rect 21266 20856 21272 20868
rect 20746 20828 21272 20856
rect 18325 20819 18383 20825
rect 21266 20816 21272 20828
rect 21324 20816 21330 20868
rect 22112 20828 22494 20856
rect 14608 20760 15700 20788
rect 14608 20748 14614 20760
rect 20990 20748 20996 20800
rect 21048 20748 21054 20800
rect 21284 20788 21312 20816
rect 22112 20788 22140 20828
rect 21284 20760 22140 20788
rect 1104 20698 26472 20720
rect 1104 20646 7252 20698
rect 7304 20646 7316 20698
rect 7368 20646 7380 20698
rect 7432 20646 7444 20698
rect 7496 20646 7508 20698
rect 7560 20646 13554 20698
rect 13606 20646 13618 20698
rect 13670 20646 13682 20698
rect 13734 20646 13746 20698
rect 13798 20646 13810 20698
rect 13862 20646 19856 20698
rect 19908 20646 19920 20698
rect 19972 20646 19984 20698
rect 20036 20646 20048 20698
rect 20100 20646 20112 20698
rect 20164 20646 26158 20698
rect 26210 20646 26222 20698
rect 26274 20646 26286 20698
rect 26338 20646 26350 20698
rect 26402 20646 26414 20698
rect 26466 20646 26472 20698
rect 1104 20624 26472 20646
rect 5350 20544 5356 20596
rect 5408 20584 5414 20596
rect 6638 20584 6644 20596
rect 5408 20556 6644 20584
rect 5408 20544 5414 20556
rect 6638 20544 6644 20556
rect 6696 20544 6702 20596
rect 6730 20544 6736 20596
rect 6788 20544 6794 20596
rect 6917 20587 6975 20593
rect 6917 20553 6929 20587
rect 6963 20584 6975 20587
rect 7098 20584 7104 20596
rect 6963 20556 7104 20584
rect 6963 20553 6975 20556
rect 6917 20547 6975 20553
rect 4890 20476 4896 20528
rect 4948 20516 4954 20528
rect 6365 20519 6423 20525
rect 6365 20516 6377 20519
rect 4948 20488 6377 20516
rect 4948 20476 4954 20488
rect 6365 20485 6377 20488
rect 6411 20485 6423 20519
rect 6932 20516 6960 20547
rect 7098 20544 7104 20556
rect 7156 20544 7162 20596
rect 9401 20587 9459 20593
rect 9401 20553 9413 20587
rect 9447 20553 9459 20587
rect 9401 20547 9459 20553
rect 11977 20587 12035 20593
rect 11977 20553 11989 20587
rect 12023 20584 12035 20587
rect 12434 20584 12440 20596
rect 12023 20556 12440 20584
rect 12023 20553 12035 20556
rect 11977 20547 12035 20553
rect 6365 20479 6423 20485
rect 6472 20488 6960 20516
rect 2317 20451 2375 20457
rect 2317 20417 2329 20451
rect 2363 20417 2375 20451
rect 2317 20411 2375 20417
rect 2593 20451 2651 20457
rect 2593 20417 2605 20451
rect 2639 20448 2651 20451
rect 3237 20451 3295 20457
rect 2639 20420 2912 20448
rect 2639 20417 2651 20420
rect 2593 20411 2651 20417
rect 2332 20380 2360 20411
rect 2774 20380 2780 20392
rect 2332 20352 2780 20380
rect 2774 20340 2780 20352
rect 2832 20340 2838 20392
rect 2884 20321 2912 20420
rect 3237 20417 3249 20451
rect 3283 20448 3295 20451
rect 4798 20448 4804 20460
rect 3283 20420 4804 20448
rect 3283 20417 3295 20420
rect 3237 20411 3295 20417
rect 4798 20408 4804 20420
rect 4856 20448 4862 20460
rect 5077 20451 5135 20457
rect 5077 20448 5089 20451
rect 4856 20420 5089 20448
rect 4856 20408 4862 20420
rect 5077 20417 5089 20420
rect 5123 20417 5135 20451
rect 5077 20411 5135 20417
rect 5442 20408 5448 20460
rect 5500 20448 5506 20460
rect 5905 20451 5963 20457
rect 5905 20448 5917 20451
rect 5500 20420 5917 20448
rect 5500 20408 5506 20420
rect 5905 20417 5917 20420
rect 5951 20417 5963 20451
rect 5905 20411 5963 20417
rect 5994 20408 6000 20460
rect 6052 20448 6058 20460
rect 6089 20451 6147 20457
rect 6089 20448 6101 20451
rect 6052 20420 6101 20448
rect 6052 20408 6058 20420
rect 6089 20417 6101 20420
rect 6135 20417 6147 20451
rect 6089 20411 6147 20417
rect 6178 20408 6184 20460
rect 6236 20448 6242 20460
rect 6472 20448 6500 20488
rect 6236 20420 6500 20448
rect 6549 20451 6607 20457
rect 6236 20408 6242 20420
rect 6549 20417 6561 20451
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 3326 20340 3332 20392
rect 3384 20340 3390 20392
rect 3513 20383 3571 20389
rect 3513 20349 3525 20383
rect 3559 20380 3571 20383
rect 3970 20380 3976 20392
rect 3559 20352 3976 20380
rect 3559 20349 3571 20352
rect 3513 20343 3571 20349
rect 3970 20340 3976 20352
rect 4028 20380 4034 20392
rect 4154 20380 4160 20392
rect 4028 20352 4160 20380
rect 4028 20340 4034 20352
rect 4154 20340 4160 20352
rect 4212 20340 4218 20392
rect 4430 20340 4436 20392
rect 4488 20380 4494 20392
rect 5169 20383 5227 20389
rect 5169 20380 5181 20383
rect 4488 20352 5181 20380
rect 4488 20340 4494 20352
rect 5169 20349 5181 20352
rect 5215 20380 5227 20383
rect 6564 20380 6592 20411
rect 6638 20408 6644 20460
rect 6696 20448 6702 20460
rect 6825 20451 6883 20457
rect 6825 20448 6837 20451
rect 6696 20420 6837 20448
rect 6696 20408 6702 20420
rect 6825 20417 6837 20420
rect 6871 20417 6883 20451
rect 6825 20411 6883 20417
rect 7009 20451 7067 20457
rect 7009 20417 7021 20451
rect 7055 20417 7067 20451
rect 7009 20411 7067 20417
rect 9309 20451 9367 20457
rect 9309 20417 9321 20451
rect 9355 20448 9367 20451
rect 9416 20448 9444 20547
rect 12434 20544 12440 20556
rect 12492 20544 12498 20596
rect 14734 20544 14740 20596
rect 14792 20584 14798 20596
rect 14829 20587 14887 20593
rect 14829 20584 14841 20587
rect 14792 20556 14841 20584
rect 14792 20544 14798 20556
rect 14829 20553 14841 20556
rect 14875 20553 14887 20587
rect 16114 20584 16120 20596
rect 14829 20547 14887 20553
rect 15856 20556 16120 20584
rect 9769 20519 9827 20525
rect 9769 20485 9781 20519
rect 9815 20516 9827 20519
rect 9950 20516 9956 20528
rect 9815 20488 9956 20516
rect 9815 20485 9827 20488
rect 9769 20479 9827 20485
rect 9950 20476 9956 20488
rect 10008 20516 10014 20528
rect 14918 20516 14924 20528
rect 10008 20488 12112 20516
rect 14582 20488 14924 20516
rect 10008 20476 10014 20488
rect 12084 20457 12112 20488
rect 14918 20476 14924 20488
rect 14976 20516 14982 20528
rect 15470 20516 15476 20528
rect 14976 20488 15476 20516
rect 14976 20476 14982 20488
rect 15470 20476 15476 20488
rect 15528 20476 15534 20528
rect 9355 20420 9444 20448
rect 9861 20451 9919 20457
rect 9355 20417 9367 20420
rect 9309 20411 9367 20417
rect 9861 20417 9873 20451
rect 9907 20448 9919 20451
rect 10321 20451 10379 20457
rect 10321 20448 10333 20451
rect 9907 20420 10333 20448
rect 9907 20417 9919 20420
rect 9861 20411 9919 20417
rect 10321 20417 10333 20420
rect 10367 20417 10379 20451
rect 10321 20411 10379 20417
rect 12069 20451 12127 20457
rect 12069 20417 12081 20451
rect 12115 20448 12127 20451
rect 12894 20448 12900 20460
rect 12115 20420 12900 20448
rect 12115 20417 12127 20420
rect 12069 20411 12127 20417
rect 5215 20352 6592 20380
rect 5215 20349 5227 20352
rect 5169 20343 5227 20349
rect 2869 20315 2927 20321
rect 2869 20281 2881 20315
rect 2915 20281 2927 20315
rect 2869 20275 2927 20281
rect 5445 20315 5503 20321
rect 5445 20281 5457 20315
rect 5491 20312 5503 20315
rect 5626 20312 5632 20324
rect 5491 20284 5632 20312
rect 5491 20281 5503 20284
rect 5445 20275 5503 20281
rect 5626 20272 5632 20284
rect 5684 20272 5690 20324
rect 5718 20272 5724 20324
rect 5776 20272 5782 20324
rect 5810 20272 5816 20324
rect 5868 20312 5874 20324
rect 7024 20312 7052 20411
rect 12894 20408 12900 20420
rect 12952 20408 12958 20460
rect 15856 20457 15884 20556
rect 16114 20544 16120 20556
rect 16172 20544 16178 20596
rect 17034 20544 17040 20596
rect 17092 20544 17098 20596
rect 17494 20544 17500 20596
rect 17552 20544 17558 20596
rect 19334 20584 19340 20596
rect 17604 20556 19340 20584
rect 15930 20476 15936 20528
rect 15988 20516 15994 20528
rect 16025 20519 16083 20525
rect 16025 20516 16037 20519
rect 15988 20488 16037 20516
rect 15988 20476 15994 20488
rect 16025 20485 16037 20488
rect 16071 20485 16083 20519
rect 16025 20479 16083 20485
rect 16390 20476 16396 20528
rect 16448 20516 16454 20528
rect 17604 20516 17632 20556
rect 19334 20544 19340 20556
rect 19392 20584 19398 20596
rect 19392 20556 22784 20584
rect 19392 20544 19398 20556
rect 18325 20519 18383 20525
rect 18325 20516 18337 20519
rect 16448 20488 17264 20516
rect 16448 20476 16454 20488
rect 15841 20451 15899 20457
rect 15841 20417 15853 20451
rect 15887 20417 15899 20451
rect 15841 20411 15899 20417
rect 16114 20408 16120 20460
rect 16172 20408 16178 20460
rect 16206 20408 16212 20460
rect 16264 20408 16270 20460
rect 17129 20451 17187 20457
rect 17129 20417 17141 20451
rect 17175 20417 17187 20451
rect 17236 20448 17264 20488
rect 17512 20488 17632 20516
rect 17696 20488 18337 20516
rect 17512 20448 17540 20488
rect 17696 20460 17724 20488
rect 18325 20485 18337 20488
rect 18371 20516 18383 20519
rect 18414 20516 18420 20528
rect 18371 20488 18420 20516
rect 18371 20485 18383 20488
rect 18325 20479 18383 20485
rect 18414 20476 18420 20488
rect 18472 20476 18478 20528
rect 22005 20519 22063 20525
rect 22005 20485 22017 20519
rect 22051 20516 22063 20519
rect 22094 20516 22100 20528
rect 22051 20488 22100 20516
rect 22051 20485 22063 20488
rect 22005 20479 22063 20485
rect 22094 20476 22100 20488
rect 22152 20476 22158 20528
rect 22756 20525 22784 20556
rect 23290 20544 23296 20596
rect 23348 20544 23354 20596
rect 25225 20587 25283 20593
rect 25225 20553 25237 20587
rect 25271 20584 25283 20587
rect 25682 20584 25688 20596
rect 25271 20556 25688 20584
rect 25271 20553 25283 20556
rect 25225 20547 25283 20553
rect 25682 20544 25688 20556
rect 25740 20544 25746 20596
rect 22741 20519 22799 20525
rect 22741 20485 22753 20519
rect 22787 20516 22799 20519
rect 23201 20519 23259 20525
rect 22787 20488 22876 20516
rect 22787 20485 22799 20488
rect 22741 20479 22799 20485
rect 22848 20460 22876 20488
rect 23201 20485 23213 20519
rect 23247 20516 23259 20519
rect 23382 20516 23388 20528
rect 23247 20488 23388 20516
rect 23247 20485 23259 20488
rect 23201 20479 23259 20485
rect 23382 20476 23388 20488
rect 23440 20476 23446 20528
rect 17586 20448 17592 20460
rect 17236 20420 17592 20448
rect 17129 20411 17187 20417
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 9953 20383 10011 20389
rect 9953 20380 9965 20383
rect 9732 20352 9965 20380
rect 9732 20340 9738 20352
rect 9953 20349 9965 20352
rect 9999 20349 10011 20383
rect 9953 20343 10011 20349
rect 10778 20340 10784 20392
rect 10836 20380 10842 20392
rect 10873 20383 10931 20389
rect 10873 20380 10885 20383
rect 10836 20352 10885 20380
rect 10836 20340 10842 20352
rect 10873 20349 10885 20352
rect 10919 20349 10931 20383
rect 10873 20343 10931 20349
rect 12250 20340 12256 20392
rect 12308 20340 12314 20392
rect 12434 20340 12440 20392
rect 12492 20380 12498 20392
rect 13078 20380 13084 20392
rect 12492 20352 13084 20380
rect 12492 20340 12498 20352
rect 13078 20340 13084 20352
rect 13136 20340 13142 20392
rect 13357 20383 13415 20389
rect 13357 20349 13369 20383
rect 13403 20380 13415 20383
rect 14090 20380 14096 20392
rect 13403 20352 14096 20380
rect 13403 20349 13415 20352
rect 13357 20343 13415 20349
rect 14090 20340 14096 20352
rect 14148 20340 14154 20392
rect 16945 20383 17003 20389
rect 16945 20349 16957 20383
rect 16991 20380 17003 20383
rect 17034 20380 17040 20392
rect 16991 20352 17040 20380
rect 16991 20349 17003 20352
rect 16945 20343 17003 20349
rect 17034 20340 17040 20352
rect 17092 20340 17098 20392
rect 17144 20380 17172 20411
rect 17586 20408 17592 20420
rect 17644 20408 17650 20460
rect 17678 20408 17684 20460
rect 17736 20408 17742 20460
rect 18046 20408 18052 20460
rect 18104 20408 18110 20460
rect 18601 20451 18659 20457
rect 18601 20448 18613 20451
rect 18156 20420 18613 20448
rect 18064 20380 18092 20408
rect 17144 20352 18092 20380
rect 5868 20284 7052 20312
rect 5868 20272 5874 20284
rect 9858 20272 9864 20324
rect 9916 20312 9922 20324
rect 10962 20312 10968 20324
rect 9916 20284 10968 20312
rect 9916 20272 9922 20284
rect 10962 20272 10968 20284
rect 11020 20312 11026 20324
rect 12066 20312 12072 20324
rect 11020 20284 12072 20312
rect 11020 20272 11026 20284
rect 12066 20272 12072 20284
rect 12124 20312 12130 20324
rect 12526 20312 12532 20324
rect 12124 20284 12532 20312
rect 12124 20272 12130 20284
rect 12526 20272 12532 20284
rect 12584 20272 12590 20324
rect 16393 20315 16451 20321
rect 16393 20281 16405 20315
rect 16439 20312 16451 20315
rect 18156 20312 18184 20420
rect 18601 20417 18613 20420
rect 18647 20417 18659 20451
rect 18601 20411 18659 20417
rect 18690 20408 18696 20460
rect 18748 20408 18754 20460
rect 18874 20408 18880 20460
rect 18932 20408 18938 20460
rect 18966 20408 18972 20460
rect 19024 20408 19030 20460
rect 19058 20408 19064 20460
rect 19116 20457 19122 20460
rect 19116 20451 19143 20457
rect 19131 20417 19143 20451
rect 19116 20411 19143 20417
rect 19116 20408 19122 20411
rect 20254 20408 20260 20460
rect 20312 20448 20318 20460
rect 20625 20451 20683 20457
rect 20625 20448 20637 20451
rect 20312 20420 20637 20448
rect 20312 20408 20318 20420
rect 20625 20417 20637 20420
rect 20671 20417 20683 20451
rect 20625 20411 20683 20417
rect 22830 20408 22836 20460
rect 22888 20408 22894 20460
rect 23842 20408 23848 20460
rect 23900 20408 23906 20460
rect 23934 20408 23940 20460
rect 23992 20408 23998 20460
rect 24026 20408 24032 20460
rect 24084 20408 24090 20460
rect 24213 20451 24271 20457
rect 24213 20417 24225 20451
rect 24259 20417 24271 20451
rect 24213 20411 24271 20417
rect 25041 20451 25099 20457
rect 25041 20417 25053 20451
rect 25087 20448 25099 20451
rect 25130 20448 25136 20460
rect 25087 20420 25136 20448
rect 25087 20417 25099 20420
rect 25041 20411 25099 20417
rect 18322 20340 18328 20392
rect 18380 20380 18386 20392
rect 18892 20380 18920 20408
rect 18380 20352 18920 20380
rect 18380 20340 18386 20352
rect 22646 20340 22652 20392
rect 22704 20380 22710 20392
rect 23385 20383 23443 20389
rect 23385 20380 23397 20383
rect 22704 20352 23397 20380
rect 22704 20340 22710 20352
rect 23385 20349 23397 20352
rect 23431 20349 23443 20383
rect 23385 20343 23443 20349
rect 24228 20312 24256 20411
rect 25130 20408 25136 20420
rect 25188 20408 25194 20460
rect 16439 20284 18184 20312
rect 21376 20284 24256 20312
rect 16439 20281 16451 20284
rect 16393 20275 16451 20281
rect 21376 20256 21404 20284
rect 2130 20204 2136 20256
rect 2188 20204 2194 20256
rect 2406 20204 2412 20256
rect 2464 20204 2470 20256
rect 9125 20247 9183 20253
rect 9125 20213 9137 20247
rect 9171 20244 9183 20247
rect 9214 20244 9220 20256
rect 9171 20216 9220 20244
rect 9171 20213 9183 20216
rect 9125 20207 9183 20213
rect 9214 20204 9220 20216
rect 9272 20204 9278 20256
rect 11606 20204 11612 20256
rect 11664 20204 11670 20256
rect 16574 20204 16580 20256
rect 16632 20244 16638 20256
rect 17678 20244 17684 20256
rect 16632 20216 17684 20244
rect 16632 20204 16638 20216
rect 17678 20204 17684 20216
rect 17736 20204 17742 20256
rect 18966 20204 18972 20256
rect 19024 20244 19030 20256
rect 19245 20247 19303 20253
rect 19245 20244 19257 20247
rect 19024 20216 19257 20244
rect 19024 20204 19030 20216
rect 19245 20213 19257 20216
rect 19291 20213 19303 20247
rect 19245 20207 19303 20213
rect 20901 20247 20959 20253
rect 20901 20213 20913 20247
rect 20947 20244 20959 20247
rect 20990 20244 20996 20256
rect 20947 20216 20996 20244
rect 20947 20213 20959 20216
rect 20901 20207 20959 20213
rect 20990 20204 20996 20216
rect 21048 20204 21054 20256
rect 21085 20247 21143 20253
rect 21085 20213 21097 20247
rect 21131 20244 21143 20247
rect 21358 20244 21364 20256
rect 21131 20216 21364 20244
rect 21131 20213 21143 20216
rect 21085 20207 21143 20213
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 21450 20204 21456 20256
rect 21508 20244 21514 20256
rect 22833 20247 22891 20253
rect 22833 20244 22845 20247
rect 21508 20216 22845 20244
rect 21508 20204 21514 20216
rect 22833 20213 22845 20216
rect 22879 20213 22891 20247
rect 22833 20207 22891 20213
rect 23658 20204 23664 20256
rect 23716 20204 23722 20256
rect 1104 20154 26312 20176
rect 1104 20102 4101 20154
rect 4153 20102 4165 20154
rect 4217 20102 4229 20154
rect 4281 20102 4293 20154
rect 4345 20102 4357 20154
rect 4409 20102 10403 20154
rect 10455 20102 10467 20154
rect 10519 20102 10531 20154
rect 10583 20102 10595 20154
rect 10647 20102 10659 20154
rect 10711 20102 16705 20154
rect 16757 20102 16769 20154
rect 16821 20102 16833 20154
rect 16885 20102 16897 20154
rect 16949 20102 16961 20154
rect 17013 20102 23007 20154
rect 23059 20102 23071 20154
rect 23123 20102 23135 20154
rect 23187 20102 23199 20154
rect 23251 20102 23263 20154
rect 23315 20102 26312 20154
rect 1104 20080 26312 20102
rect 4430 20000 4436 20052
rect 4488 20000 4494 20052
rect 4890 20000 4896 20052
rect 4948 20000 4954 20052
rect 4985 20043 5043 20049
rect 4985 20009 4997 20043
rect 5031 20040 5043 20043
rect 5442 20040 5448 20052
rect 5031 20012 5448 20040
rect 5031 20009 5043 20012
rect 4985 20003 5043 20009
rect 5442 20000 5448 20012
rect 5500 20000 5506 20052
rect 5994 20040 6000 20052
rect 5644 20012 6000 20040
rect 1857 19907 1915 19913
rect 1857 19873 1869 19907
rect 1903 19904 1915 19907
rect 2406 19904 2412 19916
rect 1903 19876 2412 19904
rect 1903 19873 1915 19876
rect 1857 19867 1915 19873
rect 2406 19864 2412 19876
rect 2464 19864 2470 19916
rect 4525 19907 4583 19913
rect 4525 19904 4537 19907
rect 4264 19876 4537 19904
rect 1578 19796 1584 19848
rect 1636 19796 1642 19848
rect 4264 19845 4292 19876
rect 4525 19873 4537 19876
rect 4571 19904 4583 19907
rect 4614 19904 4620 19916
rect 4571 19876 4620 19904
rect 4571 19873 4583 19876
rect 4525 19867 4583 19873
rect 4614 19864 4620 19876
rect 4672 19904 4678 19916
rect 5644 19904 5672 20012
rect 5994 20000 6000 20012
rect 6052 20000 6058 20052
rect 6178 20000 6184 20052
rect 6236 20040 6242 20052
rect 6914 20040 6920 20052
rect 6236 20012 6920 20040
rect 6236 20000 6242 20012
rect 6914 20000 6920 20012
rect 6972 20040 6978 20052
rect 6972 20012 7604 20040
rect 6972 20000 6978 20012
rect 4672 19876 5672 19904
rect 5920 19944 6408 19972
rect 4672 19864 4678 19876
rect 4249 19839 4307 19845
rect 4249 19805 4261 19839
rect 4295 19805 4307 19839
rect 4249 19799 4307 19805
rect 4433 19839 4491 19845
rect 4433 19805 4445 19839
rect 4479 19805 4491 19839
rect 4433 19799 4491 19805
rect 4709 19839 4767 19845
rect 4709 19805 4721 19839
rect 4755 19805 4767 19839
rect 4709 19799 4767 19805
rect 5169 19839 5227 19845
rect 5169 19805 5181 19839
rect 5215 19836 5227 19839
rect 5258 19836 5264 19848
rect 5215 19808 5264 19836
rect 5215 19805 5227 19808
rect 5169 19799 5227 19805
rect 3142 19768 3148 19780
rect 3082 19740 3148 19768
rect 3142 19728 3148 19740
rect 3200 19728 3206 19780
rect 3605 19771 3663 19777
rect 3605 19737 3617 19771
rect 3651 19737 3663 19771
rect 4448 19768 4476 19799
rect 4724 19768 4752 19799
rect 5258 19796 5264 19808
rect 5316 19796 5322 19848
rect 5350 19796 5356 19848
rect 5408 19796 5414 19848
rect 5445 19839 5503 19845
rect 5445 19805 5457 19839
rect 5491 19836 5503 19839
rect 5626 19836 5632 19848
rect 5491 19808 5632 19836
rect 5491 19805 5503 19808
rect 5445 19799 5503 19805
rect 5626 19796 5632 19808
rect 5684 19796 5690 19848
rect 5718 19796 5724 19848
rect 5776 19796 5782 19848
rect 5920 19845 5948 19944
rect 6178 19864 6184 19916
rect 6236 19864 6242 19916
rect 6270 19864 6276 19916
rect 6328 19864 6334 19916
rect 6380 19904 6408 19944
rect 6546 19904 6552 19916
rect 6380 19876 6552 19904
rect 6546 19864 6552 19876
rect 6604 19864 6610 19916
rect 7576 19904 7604 20012
rect 8018 20000 8024 20052
rect 8076 20040 8082 20052
rect 9950 20040 9956 20052
rect 8076 20012 9956 20040
rect 8076 20000 8082 20012
rect 9950 20000 9956 20012
rect 10008 20000 10014 20052
rect 10689 20043 10747 20049
rect 10689 20009 10701 20043
rect 10735 20040 10747 20043
rect 10778 20040 10784 20052
rect 10735 20012 10784 20040
rect 10735 20009 10747 20012
rect 10689 20003 10747 20009
rect 10778 20000 10784 20012
rect 10836 20000 10842 20052
rect 11606 20040 11612 20052
rect 10888 20012 11612 20040
rect 7576 19876 8156 19904
rect 8128 19848 8156 19876
rect 8294 19864 8300 19916
rect 8352 19904 8358 19916
rect 8941 19907 8999 19913
rect 8941 19904 8953 19907
rect 8352 19876 8953 19904
rect 8352 19864 8358 19876
rect 8941 19873 8953 19876
rect 8987 19873 8999 19907
rect 8941 19867 8999 19873
rect 9214 19864 9220 19916
rect 9272 19864 9278 19916
rect 5905 19839 5963 19845
rect 5905 19805 5917 19839
rect 5951 19805 5963 19839
rect 5905 19799 5963 19805
rect 8110 19796 8116 19848
rect 8168 19796 8174 19848
rect 8754 19796 8760 19848
rect 8812 19796 8818 19848
rect 10888 19845 10916 20012
rect 11606 20000 11612 20012
rect 11664 20000 11670 20052
rect 12894 20000 12900 20052
rect 12952 20000 12958 20052
rect 15838 20000 15844 20052
rect 15896 20040 15902 20052
rect 18598 20040 18604 20052
rect 15896 20012 18604 20040
rect 15896 20000 15902 20012
rect 18598 20000 18604 20012
rect 18656 20000 18662 20052
rect 23293 20043 23351 20049
rect 23293 20009 23305 20043
rect 23339 20040 23351 20043
rect 23382 20040 23388 20052
rect 23339 20012 23388 20040
rect 23339 20009 23351 20012
rect 23293 20003 23351 20009
rect 23382 20000 23388 20012
rect 23440 20000 23446 20052
rect 24486 20000 24492 20052
rect 24544 20040 24550 20052
rect 24949 20043 25007 20049
rect 24949 20040 24961 20043
rect 24544 20012 24961 20040
rect 24544 20000 24550 20012
rect 24949 20009 24961 20012
rect 24995 20009 25007 20043
rect 24949 20003 25007 20009
rect 11149 19907 11207 19913
rect 11149 19873 11161 19907
rect 11195 19904 11207 19907
rect 12434 19904 12440 19916
rect 11195 19876 12440 19904
rect 11195 19873 11207 19876
rect 11149 19867 11207 19873
rect 12434 19864 12440 19876
rect 12492 19864 12498 19916
rect 12912 19904 12940 20000
rect 13354 19932 13360 19984
rect 13412 19972 13418 19984
rect 21821 19975 21879 19981
rect 13412 19944 13584 19972
rect 13412 19932 13418 19944
rect 13556 19913 13584 19944
rect 21821 19941 21833 19975
rect 21867 19941 21879 19975
rect 21821 19935 21879 19941
rect 13449 19907 13507 19913
rect 13449 19904 13461 19907
rect 12912 19876 13461 19904
rect 13449 19873 13461 19876
rect 13495 19873 13507 19907
rect 13449 19867 13507 19873
rect 13541 19907 13599 19913
rect 13541 19873 13553 19907
rect 13587 19873 13599 19907
rect 13541 19867 13599 19873
rect 17862 19864 17868 19916
rect 17920 19864 17926 19916
rect 10873 19839 10931 19845
rect 10873 19805 10885 19839
rect 10919 19805 10931 19839
rect 10873 19799 10931 19805
rect 10962 19796 10968 19848
rect 11020 19796 11026 19848
rect 12526 19796 12532 19848
rect 12584 19836 12590 19848
rect 12894 19836 12900 19848
rect 12584 19808 12900 19836
rect 12584 19796 12590 19808
rect 12894 19796 12900 19808
rect 12952 19796 12958 19848
rect 13262 19796 13268 19848
rect 13320 19836 13326 19848
rect 14645 19839 14703 19845
rect 14645 19836 14657 19839
rect 13320 19808 14657 19836
rect 13320 19796 13326 19808
rect 14645 19805 14657 19808
rect 14691 19805 14703 19839
rect 14645 19799 14703 19805
rect 16482 19796 16488 19848
rect 16540 19836 16546 19848
rect 16853 19839 16911 19845
rect 16853 19836 16865 19839
rect 16540 19808 16865 19836
rect 16540 19796 16546 19808
rect 16853 19805 16865 19808
rect 16899 19805 16911 19839
rect 16853 19799 16911 19805
rect 18782 19796 18788 19848
rect 18840 19836 18846 19848
rect 18877 19839 18935 19845
rect 18877 19836 18889 19839
rect 18840 19808 18889 19836
rect 18840 19796 18846 19808
rect 18877 19805 18889 19808
rect 18923 19805 18935 19839
rect 18877 19799 18935 19805
rect 20901 19839 20959 19845
rect 20901 19805 20913 19839
rect 20947 19836 20959 19839
rect 21836 19836 21864 19935
rect 22465 19907 22523 19913
rect 22465 19873 22477 19907
rect 22511 19904 22523 19907
rect 22646 19904 22652 19916
rect 22511 19876 22652 19904
rect 22511 19873 22523 19876
rect 22465 19867 22523 19873
rect 22646 19864 22652 19876
rect 22704 19864 22710 19916
rect 22741 19907 22799 19913
rect 22741 19873 22753 19907
rect 22787 19873 22799 19907
rect 25041 19907 25099 19913
rect 25041 19904 25053 19907
rect 22741 19867 22799 19873
rect 22940 19876 25053 19904
rect 20947 19808 21864 19836
rect 20947 19805 20959 19808
rect 20901 19799 20959 19805
rect 22094 19796 22100 19848
rect 22152 19836 22158 19848
rect 22281 19839 22339 19845
rect 22281 19836 22293 19839
rect 22152 19808 22293 19836
rect 22152 19796 22158 19808
rect 22281 19805 22293 19808
rect 22327 19836 22339 19839
rect 22756 19836 22784 19867
rect 22940 19836 22968 19876
rect 25041 19873 25053 19876
rect 25087 19873 25099 19907
rect 25041 19867 25099 19873
rect 22327 19808 22968 19836
rect 22327 19805 22339 19808
rect 22281 19799 22339 19805
rect 23014 19796 23020 19848
rect 23072 19836 23078 19848
rect 23385 19839 23443 19845
rect 23385 19836 23397 19839
rect 23072 19808 23397 19836
rect 23072 19796 23078 19808
rect 23385 19805 23397 19808
rect 23431 19805 23443 19839
rect 23385 19799 23443 19805
rect 23474 19796 23480 19848
rect 23532 19836 23538 19848
rect 23842 19836 23848 19848
rect 23532 19808 23848 19836
rect 23532 19796 23538 19808
rect 23842 19796 23848 19808
rect 23900 19836 23906 19848
rect 24397 19839 24455 19845
rect 24397 19836 24409 19839
rect 23900 19808 24409 19836
rect 23900 19796 23906 19808
rect 24397 19805 24409 19808
rect 24443 19805 24455 19839
rect 24397 19799 24455 19805
rect 24486 19796 24492 19848
rect 24544 19836 24550 19848
rect 24673 19839 24731 19845
rect 24673 19836 24685 19839
rect 24544 19808 24685 19836
rect 24544 19796 24550 19808
rect 24673 19805 24685 19808
rect 24719 19805 24731 19839
rect 24673 19799 24731 19805
rect 24762 19796 24768 19848
rect 24820 19836 24826 19848
rect 24949 19839 25007 19845
rect 24949 19836 24961 19839
rect 24820 19808 24961 19836
rect 24820 19796 24826 19808
rect 24949 19805 24961 19808
rect 24995 19805 25007 19839
rect 24949 19799 25007 19805
rect 25222 19796 25228 19848
rect 25280 19796 25286 19848
rect 4448 19740 5212 19768
rect 3605 19731 3663 19737
rect 3620 19700 3648 19731
rect 5184 19712 5212 19740
rect 5810 19728 5816 19780
rect 5868 19728 5874 19780
rect 6043 19771 6101 19777
rect 6043 19737 6055 19771
rect 6089 19768 6101 19771
rect 6454 19768 6460 19780
rect 6089 19740 6460 19768
rect 6089 19737 6101 19740
rect 6043 19731 6101 19737
rect 6454 19728 6460 19740
rect 6512 19728 6518 19780
rect 6549 19771 6607 19777
rect 6549 19737 6561 19771
rect 6595 19737 6607 19771
rect 6549 19731 6607 19737
rect 4798 19700 4804 19712
rect 3620 19672 4804 19700
rect 4798 19660 4804 19672
rect 4856 19660 4862 19712
rect 5166 19660 5172 19712
rect 5224 19660 5230 19712
rect 5537 19703 5595 19709
rect 5537 19669 5549 19703
rect 5583 19700 5595 19703
rect 6564 19700 6592 19731
rect 7006 19728 7012 19780
rect 7064 19728 7070 19780
rect 10980 19768 11008 19796
rect 11425 19771 11483 19777
rect 11425 19768 11437 19771
rect 10442 19740 11008 19768
rect 11072 19740 11437 19768
rect 5583 19672 6592 19700
rect 5583 19669 5595 19672
rect 5537 19663 5595 19669
rect 8570 19660 8576 19712
rect 8628 19660 8634 19712
rect 11072 19709 11100 19740
rect 11425 19737 11437 19740
rect 11471 19737 11483 19771
rect 13357 19771 13415 19777
rect 11425 19731 11483 19737
rect 12728 19740 13032 19768
rect 11057 19703 11115 19709
rect 11057 19669 11069 19703
rect 11103 19669 11115 19703
rect 11057 19663 11115 19669
rect 11146 19660 11152 19712
rect 11204 19700 11210 19712
rect 12728 19700 12756 19740
rect 11204 19672 12756 19700
rect 11204 19660 11210 19672
rect 12802 19660 12808 19712
rect 12860 19700 12866 19712
rect 13004 19709 13032 19740
rect 13357 19737 13369 19771
rect 13403 19768 13415 19771
rect 14093 19771 14151 19777
rect 14093 19768 14105 19771
rect 13403 19740 14105 19768
rect 13403 19737 13415 19740
rect 13357 19731 13415 19737
rect 14093 19737 14105 19740
rect 14139 19737 14151 19771
rect 14093 19731 14151 19737
rect 22189 19771 22247 19777
rect 22189 19737 22201 19771
rect 22235 19768 22247 19771
rect 24857 19771 24915 19777
rect 24857 19768 24869 19771
rect 22235 19740 24869 19768
rect 22235 19737 22247 19740
rect 22189 19731 22247 19737
rect 24857 19737 24869 19740
rect 24903 19737 24915 19771
rect 24857 19731 24915 19737
rect 12897 19703 12955 19709
rect 12897 19700 12909 19703
rect 12860 19672 12909 19700
rect 12860 19660 12866 19672
rect 12897 19669 12909 19672
rect 12943 19669 12955 19703
rect 12897 19663 12955 19669
rect 12989 19703 13047 19709
rect 12989 19669 13001 19703
rect 13035 19669 13047 19703
rect 12989 19663 13047 19669
rect 16298 19660 16304 19712
rect 16356 19660 16362 19712
rect 17310 19660 17316 19712
rect 17368 19660 17374 19712
rect 17678 19660 17684 19712
rect 17736 19660 17742 19712
rect 17773 19703 17831 19709
rect 17773 19669 17785 19703
rect 17819 19700 17831 19703
rect 18325 19703 18383 19709
rect 18325 19700 18337 19703
rect 17819 19672 18337 19700
rect 17819 19669 17831 19672
rect 17773 19663 17831 19669
rect 18325 19669 18337 19672
rect 18371 19669 18383 19703
rect 18325 19663 18383 19669
rect 20714 19660 20720 19712
rect 20772 19660 20778 19712
rect 23842 19660 23848 19712
rect 23900 19700 23906 19712
rect 24029 19703 24087 19709
rect 24029 19700 24041 19703
rect 23900 19672 24041 19700
rect 23900 19660 23906 19672
rect 24029 19669 24041 19672
rect 24075 19669 24087 19703
rect 24029 19663 24087 19669
rect 24118 19660 24124 19712
rect 24176 19700 24182 19712
rect 24489 19703 24547 19709
rect 24489 19700 24501 19703
rect 24176 19672 24501 19700
rect 24176 19660 24182 19672
rect 24489 19669 24501 19672
rect 24535 19669 24547 19703
rect 24489 19663 24547 19669
rect 25406 19660 25412 19712
rect 25464 19660 25470 19712
rect 1104 19610 26472 19632
rect 1104 19558 7252 19610
rect 7304 19558 7316 19610
rect 7368 19558 7380 19610
rect 7432 19558 7444 19610
rect 7496 19558 7508 19610
rect 7560 19558 13554 19610
rect 13606 19558 13618 19610
rect 13670 19558 13682 19610
rect 13734 19558 13746 19610
rect 13798 19558 13810 19610
rect 13862 19558 19856 19610
rect 19908 19558 19920 19610
rect 19972 19558 19984 19610
rect 20036 19558 20048 19610
rect 20100 19558 20112 19610
rect 20164 19558 26158 19610
rect 26210 19558 26222 19610
rect 26274 19558 26286 19610
rect 26338 19558 26350 19610
rect 26402 19558 26414 19610
rect 26466 19558 26472 19610
rect 1104 19536 26472 19558
rect 2682 19496 2688 19508
rect 1596 19468 2688 19496
rect 1596 19372 1624 19468
rect 2682 19456 2688 19468
rect 2740 19456 2746 19508
rect 2774 19456 2780 19508
rect 2832 19496 2838 19508
rect 3697 19499 3755 19505
rect 3697 19496 3709 19499
rect 2832 19468 3709 19496
rect 2832 19456 2838 19468
rect 3697 19465 3709 19468
rect 3743 19465 3755 19499
rect 4065 19499 4123 19505
rect 4065 19496 4077 19499
rect 3697 19459 3755 19465
rect 3896 19468 4077 19496
rect 1857 19431 1915 19437
rect 1857 19397 1869 19431
rect 1903 19428 1915 19431
rect 2130 19428 2136 19440
rect 1903 19400 2136 19428
rect 1903 19397 1915 19400
rect 1857 19391 1915 19397
rect 2130 19388 2136 19400
rect 2188 19388 2194 19440
rect 3326 19388 3332 19440
rect 3384 19428 3390 19440
rect 3605 19431 3663 19437
rect 3605 19428 3617 19431
rect 3384 19400 3617 19428
rect 3384 19388 3390 19400
rect 3605 19397 3617 19400
rect 3651 19428 3663 19431
rect 3896 19428 3924 19468
rect 4065 19465 4077 19468
rect 4111 19496 4123 19499
rect 4614 19496 4620 19508
rect 4111 19468 4620 19496
rect 4111 19465 4123 19468
rect 4065 19459 4123 19465
rect 4614 19456 4620 19468
rect 4672 19456 4678 19508
rect 5261 19499 5319 19505
rect 5261 19465 5273 19499
rect 5307 19496 5319 19499
rect 5350 19496 5356 19508
rect 5307 19468 5356 19496
rect 5307 19465 5319 19468
rect 5261 19459 5319 19465
rect 5350 19456 5356 19468
rect 5408 19456 5414 19508
rect 5721 19499 5779 19505
rect 5721 19465 5733 19499
rect 5767 19496 5779 19499
rect 5810 19496 5816 19508
rect 5767 19468 5816 19496
rect 5767 19465 5779 19468
rect 5721 19459 5779 19465
rect 5810 19456 5816 19468
rect 5868 19456 5874 19508
rect 6086 19496 6092 19508
rect 5920 19468 6092 19496
rect 3651 19400 3924 19428
rect 3651 19397 3663 19400
rect 3605 19391 3663 19397
rect 3970 19388 3976 19440
rect 4028 19428 4034 19440
rect 4028 19400 4292 19428
rect 4028 19388 4034 19400
rect 1578 19320 1584 19372
rect 1636 19320 1642 19372
rect 3142 19360 3148 19372
rect 2990 19332 3148 19360
rect 3142 19320 3148 19332
rect 3200 19320 3206 19372
rect 4264 19301 4292 19400
rect 5166 19320 5172 19372
rect 5224 19360 5230 19372
rect 5445 19363 5503 19369
rect 5445 19360 5457 19363
rect 5224 19332 5457 19360
rect 5224 19320 5230 19332
rect 5445 19329 5457 19332
rect 5491 19329 5503 19363
rect 5445 19323 5503 19329
rect 5626 19320 5632 19372
rect 5684 19320 5690 19372
rect 5920 19369 5948 19468
rect 6086 19456 6092 19468
rect 6144 19456 6150 19508
rect 6454 19456 6460 19508
rect 6512 19496 6518 19508
rect 7101 19499 7159 19505
rect 7101 19496 7113 19499
rect 6512 19468 7113 19496
rect 6512 19456 6518 19468
rect 7101 19465 7113 19468
rect 7147 19465 7159 19499
rect 12434 19496 12440 19508
rect 7101 19459 7159 19465
rect 11532 19468 12440 19496
rect 6196 19400 6500 19428
rect 6196 19372 6224 19400
rect 5905 19363 5963 19369
rect 5905 19329 5917 19363
rect 5951 19329 5963 19363
rect 5905 19323 5963 19329
rect 6089 19363 6147 19369
rect 6089 19329 6101 19363
rect 6135 19329 6147 19363
rect 6089 19323 6147 19329
rect 4157 19295 4215 19301
rect 4157 19261 4169 19295
rect 4203 19261 4215 19295
rect 4157 19255 4215 19261
rect 4249 19295 4307 19301
rect 4249 19261 4261 19295
rect 4295 19261 4307 19295
rect 4249 19255 4307 19261
rect 4172 19224 4200 19255
rect 6104 19224 6132 19323
rect 6178 19320 6184 19372
rect 6236 19320 6242 19372
rect 6362 19320 6368 19372
rect 6420 19320 6426 19372
rect 6472 19369 6500 19400
rect 8570 19388 8576 19440
rect 8628 19428 8634 19440
rect 8665 19431 8723 19437
rect 8665 19428 8677 19431
rect 8628 19400 8677 19428
rect 8628 19388 8634 19400
rect 8665 19397 8677 19400
rect 8711 19397 8723 19431
rect 8665 19391 8723 19397
rect 9674 19388 9680 19440
rect 9732 19388 9738 19440
rect 6457 19363 6515 19369
rect 6457 19329 6469 19363
rect 6503 19329 6515 19363
rect 6457 19323 6515 19329
rect 7745 19363 7803 19369
rect 7745 19329 7757 19363
rect 7791 19360 7803 19363
rect 8018 19360 8024 19372
rect 7791 19332 8024 19360
rect 7791 19329 7803 19332
rect 7745 19323 7803 19329
rect 8018 19320 8024 19332
rect 8076 19320 8082 19372
rect 8294 19320 8300 19372
rect 8352 19360 8358 19372
rect 8389 19363 8447 19369
rect 8389 19360 8401 19363
rect 8352 19332 8401 19360
rect 8352 19320 8358 19332
rect 8389 19329 8401 19332
rect 8435 19329 8447 19363
rect 8389 19323 8447 19329
rect 11146 19320 11152 19372
rect 11204 19320 11210 19372
rect 11532 19369 11560 19468
rect 12434 19456 12440 19468
rect 12492 19496 12498 19508
rect 12492 19468 14780 19496
rect 12492 19456 12498 19468
rect 14752 19372 14780 19468
rect 16482 19456 16488 19508
rect 16540 19456 16546 19508
rect 16574 19456 16580 19508
rect 16632 19456 16638 19508
rect 17310 19456 17316 19508
rect 17368 19456 17374 19508
rect 17770 19456 17776 19508
rect 17828 19496 17834 19508
rect 18414 19496 18420 19508
rect 17828 19468 18420 19496
rect 17828 19456 17834 19468
rect 18414 19456 18420 19468
rect 18472 19456 18478 19508
rect 21637 19499 21695 19505
rect 21637 19465 21649 19499
rect 21683 19496 21695 19499
rect 22094 19496 22100 19508
rect 21683 19468 22100 19496
rect 21683 19465 21695 19468
rect 21637 19459 21695 19465
rect 22094 19456 22100 19468
rect 22152 19456 22158 19508
rect 24026 19456 24032 19508
rect 24084 19496 24090 19508
rect 24397 19499 24455 19505
rect 24397 19496 24409 19499
rect 24084 19468 24409 19496
rect 24084 19456 24090 19468
rect 24397 19465 24409 19468
rect 24443 19465 24455 19499
rect 24397 19459 24455 19465
rect 15470 19388 15476 19440
rect 15528 19388 15534 19440
rect 11517 19363 11575 19369
rect 11517 19329 11529 19363
rect 11563 19329 11575 19363
rect 11517 19323 11575 19329
rect 12894 19320 12900 19372
rect 12952 19320 12958 19372
rect 14734 19320 14740 19372
rect 14792 19320 14798 19372
rect 9398 19252 9404 19304
rect 9456 19292 9462 19304
rect 10137 19295 10195 19301
rect 9456 19264 10088 19292
rect 9456 19252 9462 19264
rect 4172 19196 6132 19224
rect 10060 19224 10088 19264
rect 10137 19261 10149 19295
rect 10183 19292 10195 19295
rect 10318 19292 10324 19304
rect 10183 19264 10324 19292
rect 10183 19261 10195 19264
rect 10137 19255 10195 19261
rect 10318 19252 10324 19264
rect 10376 19292 10382 19304
rect 10781 19295 10839 19301
rect 10781 19292 10793 19295
rect 10376 19264 10793 19292
rect 10376 19252 10382 19264
rect 10781 19261 10793 19264
rect 10827 19261 10839 19295
rect 11793 19295 11851 19301
rect 11793 19292 11805 19295
rect 10781 19255 10839 19261
rect 11348 19264 11805 19292
rect 11348 19233 11376 19264
rect 11793 19261 11805 19264
rect 11839 19261 11851 19295
rect 11793 19255 11851 19261
rect 12158 19252 12164 19304
rect 12216 19292 12222 19304
rect 14642 19292 14648 19304
rect 12216 19264 14648 19292
rect 12216 19252 12222 19264
rect 14642 19252 14648 19264
rect 14700 19252 14706 19304
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19292 15071 19295
rect 15102 19292 15108 19304
rect 15059 19264 15108 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 15102 19252 15108 19264
rect 15160 19252 15166 19304
rect 16592 19292 16620 19456
rect 17328 19428 17356 19456
rect 16868 19400 17356 19428
rect 17788 19428 17816 19456
rect 17788 19400 17894 19428
rect 16868 19369 16896 19400
rect 22830 19388 22836 19440
rect 22888 19388 22894 19440
rect 16853 19363 16911 19369
rect 16853 19329 16865 19363
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 21266 19320 21272 19372
rect 21324 19360 21330 19372
rect 21910 19360 21916 19372
rect 21324 19332 21916 19360
rect 21324 19320 21330 19332
rect 21910 19320 21916 19332
rect 21968 19320 21974 19372
rect 22738 19320 22744 19372
rect 22796 19360 22802 19372
rect 23014 19360 23020 19372
rect 22796 19332 23020 19360
rect 22796 19320 22802 19332
rect 23014 19320 23020 19332
rect 23072 19320 23078 19372
rect 23658 19320 23664 19372
rect 23716 19360 23722 19372
rect 24213 19363 24271 19369
rect 24213 19360 24225 19363
rect 23716 19332 24225 19360
rect 23716 19320 23722 19332
rect 24213 19329 24225 19332
rect 24259 19329 24271 19363
rect 24213 19323 24271 19329
rect 25041 19363 25099 19369
rect 25041 19329 25053 19363
rect 25087 19360 25099 19363
rect 25222 19360 25228 19372
rect 25087 19332 25228 19360
rect 25087 19329 25099 19332
rect 25041 19323 25099 19329
rect 25222 19320 25228 19332
rect 25280 19320 25286 19372
rect 17126 19292 17132 19304
rect 16592 19264 17132 19292
rect 17126 19252 17132 19264
rect 17184 19252 17190 19304
rect 17405 19295 17463 19301
rect 17405 19292 17417 19295
rect 17236 19264 17417 19292
rect 11333 19227 11391 19233
rect 10060 19196 11284 19224
rect 6012 19168 6040 19196
rect 5994 19116 6000 19168
rect 6052 19116 6058 19168
rect 10226 19116 10232 19168
rect 10284 19116 10290 19168
rect 11256 19156 11284 19196
rect 11333 19193 11345 19227
rect 11379 19193 11391 19227
rect 11333 19187 11391 19193
rect 13262 19184 13268 19236
rect 13320 19184 13326 19236
rect 17037 19227 17095 19233
rect 17037 19193 17049 19227
rect 17083 19224 17095 19227
rect 17236 19224 17264 19264
rect 17405 19261 17417 19264
rect 17451 19261 17463 19295
rect 17405 19255 17463 19261
rect 18874 19252 18880 19304
rect 18932 19292 18938 19304
rect 19153 19295 19211 19301
rect 19153 19292 19165 19295
rect 18932 19264 19165 19292
rect 18932 19252 18938 19264
rect 19153 19261 19165 19264
rect 19199 19261 19211 19295
rect 19153 19255 19211 19261
rect 19889 19295 19947 19301
rect 19889 19261 19901 19295
rect 19935 19261 19947 19295
rect 19889 19255 19947 19261
rect 20165 19295 20223 19301
rect 20165 19261 20177 19295
rect 20211 19292 20223 19295
rect 20714 19292 20720 19304
rect 20211 19264 20720 19292
rect 20211 19261 20223 19264
rect 20165 19255 20223 19261
rect 17083 19196 17264 19224
rect 17083 19193 17095 19196
rect 17037 19187 17095 19193
rect 12158 19156 12164 19168
rect 11256 19128 12164 19156
rect 12158 19116 12164 19128
rect 12216 19116 12222 19168
rect 12250 19116 12256 19168
rect 12308 19156 12314 19168
rect 16942 19156 16948 19168
rect 12308 19128 16948 19156
rect 12308 19116 12314 19128
rect 16942 19116 16948 19128
rect 17000 19116 17006 19168
rect 18138 19116 18144 19168
rect 18196 19156 18202 19168
rect 18782 19156 18788 19168
rect 18196 19128 18788 19156
rect 18196 19116 18202 19128
rect 18782 19116 18788 19128
rect 18840 19156 18846 19168
rect 18877 19159 18935 19165
rect 18877 19156 18889 19159
rect 18840 19128 18889 19156
rect 18840 19116 18846 19128
rect 18877 19125 18889 19128
rect 18923 19125 18935 19159
rect 18877 19119 18935 19125
rect 19610 19116 19616 19168
rect 19668 19156 19674 19168
rect 19797 19159 19855 19165
rect 19797 19156 19809 19159
rect 19668 19128 19809 19156
rect 19668 19116 19674 19128
rect 19797 19125 19809 19128
rect 19843 19125 19855 19159
rect 19904 19156 19932 19255
rect 20714 19252 20720 19264
rect 20772 19252 20778 19304
rect 22002 19252 22008 19304
rect 22060 19292 22066 19304
rect 22097 19295 22155 19301
rect 22097 19292 22109 19295
rect 22060 19264 22109 19292
rect 22060 19252 22066 19264
rect 22097 19261 22109 19264
rect 22143 19261 22155 19295
rect 22097 19255 22155 19261
rect 23474 19252 23480 19304
rect 23532 19292 23538 19304
rect 24486 19292 24492 19304
rect 23532 19264 24492 19292
rect 23532 19252 23538 19264
rect 24486 19252 24492 19264
rect 24544 19252 24550 19304
rect 20714 19156 20720 19168
rect 19904 19128 20720 19156
rect 19797 19119 19855 19125
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 22925 19159 22983 19165
rect 22925 19156 22937 19159
rect 22152 19128 22937 19156
rect 22152 19116 22158 19128
rect 22925 19125 22937 19128
rect 22971 19125 22983 19159
rect 22925 19119 22983 19125
rect 23658 19116 23664 19168
rect 23716 19116 23722 19168
rect 1104 19066 26312 19088
rect 1104 19014 4101 19066
rect 4153 19014 4165 19066
rect 4217 19014 4229 19066
rect 4281 19014 4293 19066
rect 4345 19014 4357 19066
rect 4409 19014 10403 19066
rect 10455 19014 10467 19066
rect 10519 19014 10531 19066
rect 10583 19014 10595 19066
rect 10647 19014 10659 19066
rect 10711 19014 16705 19066
rect 16757 19014 16769 19066
rect 16821 19014 16833 19066
rect 16885 19014 16897 19066
rect 16949 19014 16961 19066
rect 17013 19014 23007 19066
rect 23059 19014 23071 19066
rect 23123 19014 23135 19066
rect 23187 19014 23199 19066
rect 23251 19014 23263 19066
rect 23315 19014 26312 19066
rect 1104 18992 26312 19014
rect 5166 18912 5172 18964
rect 5224 18912 5230 18964
rect 5626 18912 5632 18964
rect 5684 18952 5690 18964
rect 5721 18955 5779 18961
rect 5721 18952 5733 18955
rect 5684 18924 5733 18952
rect 5684 18912 5690 18924
rect 5721 18921 5733 18924
rect 5767 18921 5779 18955
rect 5721 18915 5779 18921
rect 8754 18912 8760 18964
rect 8812 18952 8818 18964
rect 9309 18955 9367 18961
rect 9309 18952 9321 18955
rect 8812 18924 9321 18952
rect 8812 18912 8818 18924
rect 9309 18921 9321 18924
rect 9355 18921 9367 18955
rect 9309 18915 9367 18921
rect 10778 18912 10784 18964
rect 10836 18912 10842 18964
rect 10870 18912 10876 18964
rect 10928 18952 10934 18964
rect 14921 18955 14979 18961
rect 10928 18924 12664 18952
rect 10928 18912 10934 18924
rect 1578 18776 1584 18828
rect 1636 18776 1642 18828
rect 5994 18816 6000 18828
rect 5368 18788 6000 18816
rect 3605 18751 3663 18757
rect 3605 18717 3617 18751
rect 3651 18748 3663 18751
rect 4154 18748 4160 18760
rect 3651 18720 4160 18748
rect 3651 18717 3663 18720
rect 3605 18711 3663 18717
rect 4154 18708 4160 18720
rect 4212 18748 4218 18760
rect 4982 18748 4988 18760
rect 4212 18720 4988 18748
rect 4212 18708 4218 18720
rect 4982 18708 4988 18720
rect 5040 18748 5046 18760
rect 5368 18757 5396 18788
rect 5994 18776 6000 18788
rect 6052 18776 6058 18828
rect 9398 18776 9404 18828
rect 9456 18816 9462 18828
rect 9861 18819 9919 18825
rect 9861 18816 9873 18819
rect 9456 18788 9873 18816
rect 9456 18776 9462 18788
rect 9861 18785 9873 18788
rect 9907 18785 9919 18819
rect 10796 18816 10824 18912
rect 9861 18779 9919 18785
rect 10704 18788 10824 18816
rect 5353 18751 5411 18757
rect 5353 18748 5365 18751
rect 5040 18720 5365 18748
rect 5040 18708 5046 18720
rect 5353 18717 5365 18720
rect 5399 18717 5411 18751
rect 5353 18711 5411 18717
rect 5537 18751 5595 18757
rect 5537 18717 5549 18751
rect 5583 18717 5595 18751
rect 5537 18711 5595 18717
rect 1854 18640 1860 18692
rect 1912 18640 1918 18692
rect 3234 18680 3240 18692
rect 3082 18652 3240 18680
rect 3234 18640 3240 18652
rect 3292 18640 3298 18692
rect 5552 18680 5580 18711
rect 5626 18708 5632 18760
rect 5684 18708 5690 18760
rect 5721 18751 5779 18757
rect 5721 18717 5733 18751
rect 5767 18717 5779 18751
rect 5721 18711 5779 18717
rect 5736 18680 5764 18711
rect 5810 18708 5816 18760
rect 5868 18708 5874 18760
rect 9677 18751 9735 18757
rect 9677 18717 9689 18751
rect 9723 18748 9735 18751
rect 10226 18748 10232 18760
rect 9723 18720 10232 18748
rect 9723 18717 9735 18720
rect 9677 18711 9735 18717
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 10318 18708 10324 18760
rect 10376 18748 10382 18760
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 10376 18720 10425 18748
rect 10376 18708 10382 18720
rect 10413 18717 10425 18720
rect 10459 18717 10471 18751
rect 10597 18751 10655 18757
rect 10597 18748 10609 18751
rect 10413 18711 10471 18717
rect 10520 18720 10609 18748
rect 5552 18652 5764 18680
rect 5736 18612 5764 18652
rect 9769 18683 9827 18689
rect 9769 18649 9781 18683
rect 9815 18680 9827 18683
rect 9950 18680 9956 18692
rect 9815 18652 9956 18680
rect 9815 18649 9827 18652
rect 9769 18643 9827 18649
rect 9950 18640 9956 18652
rect 10008 18640 10014 18692
rect 6178 18612 6184 18624
rect 5736 18584 6184 18612
rect 6178 18572 6184 18584
rect 6236 18572 6242 18624
rect 10226 18572 10232 18624
rect 10284 18612 10290 18624
rect 10520 18612 10548 18720
rect 10597 18717 10609 18720
rect 10643 18717 10655 18751
rect 10597 18711 10655 18717
rect 10704 18689 10732 18788
rect 10778 18708 10784 18760
rect 10836 18748 10842 18760
rect 10888 18748 10916 18912
rect 10965 18887 11023 18893
rect 10965 18853 10977 18887
rect 11011 18853 11023 18887
rect 10965 18847 11023 18853
rect 10836 18720 10916 18748
rect 10980 18748 11008 18847
rect 12526 18844 12532 18896
rect 12584 18844 12590 18896
rect 12636 18884 12664 18924
rect 14921 18921 14933 18955
rect 14967 18952 14979 18955
rect 15102 18952 15108 18964
rect 14967 18924 15108 18952
rect 14967 18921 14979 18924
rect 14921 18915 14979 18921
rect 15102 18912 15108 18924
rect 15160 18912 15166 18964
rect 16206 18952 16212 18964
rect 16132 18924 16212 18952
rect 15378 18884 15384 18896
rect 12636 18856 15384 18884
rect 15378 18844 15384 18856
rect 15436 18844 15442 18896
rect 15562 18844 15568 18896
rect 15620 18844 15626 18896
rect 15657 18887 15715 18893
rect 15657 18853 15669 18887
rect 15703 18853 15715 18887
rect 15657 18847 15715 18853
rect 13262 18816 13268 18828
rect 12268 18788 13268 18816
rect 11885 18751 11943 18757
rect 11885 18748 11897 18751
rect 10980 18720 11897 18748
rect 10836 18708 10842 18720
rect 11885 18717 11897 18720
rect 11931 18717 11943 18751
rect 11885 18711 11943 18717
rect 12033 18751 12091 18757
rect 12033 18717 12045 18751
rect 12079 18748 12091 18751
rect 12268 18748 12296 18788
rect 13262 18776 13268 18788
rect 13320 18776 13326 18828
rect 15672 18816 15700 18847
rect 16132 18816 16160 18924
rect 16206 18912 16212 18924
rect 16264 18952 16270 18964
rect 19334 18952 19340 18964
rect 16264 18924 19340 18952
rect 16264 18912 16270 18924
rect 14752 18788 15700 18816
rect 15764 18788 16160 18816
rect 12079 18720 12296 18748
rect 12391 18751 12449 18757
rect 12079 18717 12091 18720
rect 12033 18711 12091 18717
rect 12391 18717 12403 18751
rect 12437 18748 12449 18751
rect 12710 18748 12716 18760
rect 12437 18720 12716 18748
rect 12437 18717 12449 18720
rect 12391 18711 12449 18717
rect 12710 18708 12716 18720
rect 12768 18708 12774 18760
rect 14752 18757 14780 18788
rect 14737 18751 14795 18757
rect 14737 18717 14749 18751
rect 14783 18717 14795 18751
rect 14737 18711 14795 18717
rect 15010 18708 15016 18760
rect 15068 18708 15074 18760
rect 15378 18708 15384 18760
rect 15436 18748 15442 18760
rect 15764 18748 15792 18788
rect 16206 18776 16212 18828
rect 16264 18776 16270 18828
rect 15436 18720 15792 18748
rect 16025 18751 16083 18757
rect 15436 18708 15442 18720
rect 16025 18717 16037 18751
rect 16071 18748 16083 18751
rect 16298 18748 16304 18760
rect 16071 18720 16304 18748
rect 16071 18717 16083 18720
rect 16025 18711 16083 18717
rect 16298 18708 16304 18720
rect 16356 18708 16362 18760
rect 16482 18708 16488 18760
rect 16540 18708 16546 18760
rect 16853 18751 16911 18757
rect 16853 18717 16865 18751
rect 16899 18748 16911 18751
rect 16960 18748 16988 18924
rect 19334 18912 19340 18924
rect 19392 18912 19398 18964
rect 22189 18955 22247 18961
rect 22189 18921 22201 18955
rect 22235 18952 22247 18955
rect 23474 18952 23480 18964
rect 22235 18924 23480 18952
rect 22235 18921 22247 18924
rect 22189 18915 22247 18921
rect 23474 18912 23480 18924
rect 23532 18912 23538 18964
rect 18506 18844 18512 18896
rect 18564 18884 18570 18896
rect 18564 18856 19840 18884
rect 18564 18844 18570 18856
rect 17126 18776 17132 18828
rect 17184 18776 17190 18828
rect 17770 18776 17776 18828
rect 17828 18816 17834 18828
rect 19812 18825 19840 18856
rect 19705 18819 19763 18825
rect 19705 18816 19717 18819
rect 17828 18788 19717 18816
rect 17828 18776 17834 18788
rect 19705 18785 19717 18788
rect 19751 18785 19763 18819
rect 19705 18779 19763 18785
rect 19797 18819 19855 18825
rect 19797 18785 19809 18819
rect 19843 18785 19855 18819
rect 19797 18779 19855 18785
rect 20441 18819 20499 18825
rect 20441 18785 20453 18819
rect 20487 18816 20499 18819
rect 20714 18816 20720 18828
rect 20487 18788 20720 18816
rect 20487 18785 20499 18788
rect 20441 18779 20499 18785
rect 20714 18776 20720 18788
rect 20772 18816 20778 18828
rect 22002 18816 22008 18828
rect 20772 18788 22008 18816
rect 20772 18776 20778 18788
rect 22002 18776 22008 18788
rect 22060 18816 22066 18828
rect 22373 18819 22431 18825
rect 22373 18816 22385 18819
rect 22060 18788 22385 18816
rect 22060 18776 22066 18788
rect 22373 18785 22385 18788
rect 22419 18785 22431 18819
rect 22373 18779 22431 18785
rect 22741 18819 22799 18825
rect 22741 18785 22753 18819
rect 22787 18816 22799 18819
rect 23658 18816 23664 18828
rect 22787 18788 23664 18816
rect 22787 18785 22799 18788
rect 22741 18779 22799 18785
rect 23658 18776 23664 18788
rect 23716 18776 23722 18828
rect 16899 18720 16988 18748
rect 16899 18717 16911 18720
rect 16853 18711 16911 18717
rect 19610 18708 19616 18760
rect 19668 18708 19674 18760
rect 24167 18751 24225 18757
rect 24167 18717 24179 18751
rect 24213 18748 24225 18751
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 24213 18720 24593 18748
rect 24213 18717 24225 18720
rect 24167 18711 24225 18717
rect 24581 18717 24593 18720
rect 24627 18748 24639 18751
rect 25222 18748 25228 18760
rect 24627 18720 25228 18748
rect 24627 18717 24639 18720
rect 24581 18711 24639 18717
rect 25222 18708 25228 18720
rect 25280 18708 25286 18760
rect 10689 18683 10747 18689
rect 10689 18649 10701 18683
rect 10735 18649 10747 18683
rect 10689 18643 10747 18649
rect 12158 18640 12164 18692
rect 12216 18640 12222 18692
rect 12253 18683 12311 18689
rect 12253 18649 12265 18683
rect 12299 18680 12311 18683
rect 12802 18680 12808 18692
rect 12299 18652 12808 18680
rect 12299 18649 12311 18652
rect 12253 18643 12311 18649
rect 12802 18640 12808 18652
rect 12860 18640 12866 18692
rect 15197 18683 15255 18689
rect 15197 18649 15209 18683
rect 15243 18649 15255 18683
rect 15197 18643 15255 18649
rect 10594 18612 10600 18624
rect 10284 18584 10600 18612
rect 10284 18572 10290 18584
rect 10594 18572 10600 18584
rect 10652 18612 10658 18624
rect 15212 18612 15240 18643
rect 15286 18640 15292 18692
rect 15344 18640 15350 18692
rect 15562 18640 15568 18692
rect 15620 18680 15626 18692
rect 16574 18680 16580 18692
rect 15620 18652 16580 18680
rect 15620 18640 15626 18652
rect 16574 18640 16580 18652
rect 16632 18640 16638 18692
rect 16666 18640 16672 18692
rect 16724 18640 16730 18692
rect 16761 18683 16819 18689
rect 16761 18649 16773 18683
rect 16807 18680 16819 18683
rect 16807 18652 17356 18680
rect 16807 18649 16819 18652
rect 16761 18643 16819 18649
rect 15930 18612 15936 18624
rect 10652 18584 15936 18612
rect 10652 18572 10658 18584
rect 15930 18572 15936 18584
rect 15988 18572 15994 18624
rect 16114 18572 16120 18624
rect 16172 18572 16178 18624
rect 17034 18572 17040 18624
rect 17092 18572 17098 18624
rect 17328 18612 17356 18652
rect 17402 18640 17408 18692
rect 17460 18640 17466 18692
rect 18414 18640 18420 18692
rect 18472 18640 18478 18692
rect 20717 18683 20775 18689
rect 20717 18649 20729 18683
rect 20763 18680 20775 18683
rect 20990 18680 20996 18692
rect 20763 18652 20996 18680
rect 20763 18649 20775 18652
rect 20717 18643 20775 18649
rect 20990 18640 20996 18652
rect 21048 18640 21054 18692
rect 21942 18652 22048 18680
rect 22020 18624 22048 18652
rect 22112 18652 22324 18680
rect 18138 18612 18144 18624
rect 17328 18584 18144 18612
rect 18138 18572 18144 18584
rect 18196 18572 18202 18624
rect 18874 18572 18880 18624
rect 18932 18572 18938 18624
rect 19242 18572 19248 18624
rect 19300 18572 19306 18624
rect 22002 18572 22008 18624
rect 22060 18612 22066 18624
rect 22112 18612 22140 18652
rect 22060 18584 22140 18612
rect 22296 18612 22324 18652
rect 23032 18652 23138 18680
rect 23032 18612 23060 18652
rect 22296 18584 23060 18612
rect 22060 18572 22066 18584
rect 24486 18572 24492 18624
rect 24544 18572 24550 18624
rect 1104 18522 26472 18544
rect 1104 18470 7252 18522
rect 7304 18470 7316 18522
rect 7368 18470 7380 18522
rect 7432 18470 7444 18522
rect 7496 18470 7508 18522
rect 7560 18470 13554 18522
rect 13606 18470 13618 18522
rect 13670 18470 13682 18522
rect 13734 18470 13746 18522
rect 13798 18470 13810 18522
rect 13862 18470 19856 18522
rect 19908 18470 19920 18522
rect 19972 18470 19984 18522
rect 20036 18470 20048 18522
rect 20100 18470 20112 18522
rect 20164 18470 26158 18522
rect 26210 18470 26222 18522
rect 26274 18470 26286 18522
rect 26338 18470 26350 18522
rect 26402 18470 26414 18522
rect 26466 18470 26472 18522
rect 1104 18448 26472 18470
rect 1854 18368 1860 18420
rect 1912 18408 1918 18420
rect 2225 18411 2283 18417
rect 2225 18408 2237 18411
rect 1912 18380 2237 18408
rect 1912 18368 1918 18380
rect 2225 18377 2237 18380
rect 2271 18377 2283 18411
rect 2225 18371 2283 18377
rect 2685 18411 2743 18417
rect 2685 18377 2697 18411
rect 2731 18377 2743 18411
rect 2685 18371 2743 18377
rect 2409 18275 2467 18281
rect 2409 18241 2421 18275
rect 2455 18272 2467 18275
rect 2700 18272 2728 18371
rect 3510 18368 3516 18420
rect 3568 18368 3574 18420
rect 4154 18368 4160 18420
rect 4212 18368 4218 18420
rect 6914 18368 6920 18420
rect 6972 18368 6978 18420
rect 8202 18368 8208 18420
rect 8260 18368 8266 18420
rect 9493 18411 9551 18417
rect 9493 18377 9505 18411
rect 9539 18408 9551 18411
rect 16114 18408 16120 18420
rect 9539 18380 16120 18408
rect 9539 18377 9551 18380
rect 9493 18371 9551 18377
rect 3053 18343 3111 18349
rect 3053 18309 3065 18343
rect 3099 18340 3111 18343
rect 4172 18340 4200 18368
rect 8220 18340 8248 18368
rect 9674 18340 9680 18352
rect 3099 18312 4200 18340
rect 7760 18312 8248 18340
rect 9246 18312 9680 18340
rect 3099 18309 3111 18312
rect 3053 18303 3111 18309
rect 2455 18244 2728 18272
rect 3145 18275 3203 18281
rect 2455 18241 2467 18244
rect 2409 18235 2467 18241
rect 3145 18241 3157 18275
rect 3191 18272 3203 18275
rect 3510 18272 3516 18284
rect 3191 18244 3516 18272
rect 3191 18241 3203 18244
rect 3145 18235 3203 18241
rect 3510 18232 3516 18244
rect 3568 18232 3574 18284
rect 4614 18232 4620 18284
rect 4672 18272 4678 18284
rect 5353 18275 5411 18281
rect 5353 18272 5365 18275
rect 4672 18244 5365 18272
rect 4672 18232 4678 18244
rect 5353 18241 5365 18244
rect 5399 18241 5411 18275
rect 5353 18235 5411 18241
rect 5537 18275 5595 18281
rect 5537 18241 5549 18275
rect 5583 18272 5595 18275
rect 5902 18272 5908 18284
rect 5583 18244 5908 18272
rect 5583 18241 5595 18244
rect 5537 18235 5595 18241
rect 5902 18232 5908 18244
rect 5960 18232 5966 18284
rect 6362 18232 6368 18284
rect 6420 18272 6426 18284
rect 6549 18275 6607 18281
rect 6549 18272 6561 18275
rect 6420 18244 6561 18272
rect 6420 18232 6426 18244
rect 6549 18241 6561 18244
rect 6595 18241 6607 18275
rect 6549 18235 6607 18241
rect 6641 18275 6699 18281
rect 6641 18241 6653 18275
rect 6687 18272 6699 18275
rect 6822 18272 6828 18284
rect 6687 18244 6828 18272
rect 6687 18241 6699 18244
rect 6641 18235 6699 18241
rect 6822 18232 6828 18244
rect 6880 18232 6886 18284
rect 7760 18281 7788 18312
rect 9508 18284 9536 18312
rect 9674 18300 9680 18312
rect 9732 18300 9738 18352
rect 7745 18275 7803 18281
rect 7745 18241 7757 18275
rect 7791 18241 7803 18275
rect 7745 18235 7803 18241
rect 9490 18232 9496 18284
rect 9548 18232 9554 18284
rect 10152 18272 10180 18380
rect 16114 18368 16120 18380
rect 16172 18368 16178 18420
rect 17402 18368 17408 18420
rect 17460 18368 17466 18420
rect 19242 18408 19248 18420
rect 18156 18380 19248 18408
rect 10594 18300 10600 18352
rect 10652 18300 10658 18352
rect 10689 18343 10747 18349
rect 10689 18309 10701 18343
rect 10735 18340 10747 18343
rect 10735 18312 10916 18340
rect 10735 18309 10747 18312
rect 10689 18303 10747 18309
rect 10888 18284 10916 18312
rect 12158 18300 12164 18352
rect 12216 18340 12222 18352
rect 15470 18340 15476 18352
rect 12216 18312 12572 18340
rect 14858 18312 15476 18340
rect 12216 18300 12222 18312
rect 10229 18275 10287 18281
rect 10229 18272 10241 18275
rect 10152 18244 10241 18272
rect 10229 18241 10241 18244
rect 10275 18241 10287 18275
rect 10229 18235 10287 18241
rect 10413 18275 10471 18281
rect 10413 18241 10425 18275
rect 10459 18241 10471 18275
rect 10413 18235 10471 18241
rect 3326 18164 3332 18216
rect 3384 18204 3390 18216
rect 3970 18204 3976 18216
rect 3384 18176 3976 18204
rect 3384 18164 3390 18176
rect 3970 18164 3976 18176
rect 4028 18164 4034 18216
rect 4157 18207 4215 18213
rect 4157 18173 4169 18207
rect 4203 18204 4215 18207
rect 4430 18204 4436 18216
rect 4203 18176 4436 18204
rect 4203 18173 4215 18176
rect 4157 18167 4215 18173
rect 4430 18164 4436 18176
rect 4488 18164 4494 18216
rect 6178 18164 6184 18216
rect 6236 18164 6242 18216
rect 6454 18164 6460 18216
rect 6512 18164 6518 18216
rect 6733 18207 6791 18213
rect 6733 18173 6745 18207
rect 6779 18173 6791 18207
rect 6733 18167 6791 18173
rect 1946 18096 1952 18148
rect 2004 18136 2010 18148
rect 6196 18136 6224 18164
rect 6748 18136 6776 18167
rect 8018 18164 8024 18216
rect 8076 18164 8082 18216
rect 10134 18164 10140 18216
rect 10192 18204 10198 18216
rect 10428 18204 10456 18235
rect 10778 18232 10784 18284
rect 10836 18232 10842 18284
rect 10870 18232 10876 18284
rect 10928 18232 10934 18284
rect 12544 18281 12572 18312
rect 15470 18300 15476 18312
rect 15528 18300 15534 18352
rect 15930 18300 15936 18352
rect 15988 18340 15994 18352
rect 16666 18340 16672 18352
rect 15988 18312 16672 18340
rect 15988 18300 15994 18312
rect 16666 18300 16672 18312
rect 16724 18340 16730 18352
rect 17770 18340 17776 18352
rect 16724 18312 17776 18340
rect 16724 18300 16730 18312
rect 17770 18300 17776 18312
rect 17828 18300 17834 18352
rect 12253 18275 12311 18281
rect 12253 18272 12265 18275
rect 10980 18244 12265 18272
rect 10192 18176 10456 18204
rect 10192 18164 10198 18176
rect 10980 18145 11008 18244
rect 12253 18241 12265 18244
rect 12299 18241 12311 18275
rect 12253 18235 12311 18241
rect 12391 18275 12449 18281
rect 12391 18241 12403 18275
rect 12437 18241 12449 18275
rect 12391 18235 12449 18241
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18241 12587 18275
rect 12529 18235 12587 18241
rect 2004 18108 5671 18136
rect 6196 18108 6776 18136
rect 10965 18139 11023 18145
rect 2004 18096 2010 18108
rect 5534 18028 5540 18080
rect 5592 18028 5598 18080
rect 5643 18068 5671 18108
rect 10965 18105 10977 18139
rect 11011 18105 11023 18139
rect 10965 18099 11023 18105
rect 12406 18080 12434 18235
rect 12544 18204 12572 18235
rect 12618 18232 12624 18284
rect 12676 18232 12682 18284
rect 12710 18232 12716 18284
rect 12768 18281 12774 18284
rect 12768 18272 12776 18281
rect 12768 18244 12813 18272
rect 12768 18235 12776 18244
rect 12768 18232 12774 18235
rect 15286 18232 15292 18284
rect 15344 18272 15350 18284
rect 15838 18272 15844 18284
rect 15344 18244 15844 18272
rect 15344 18232 15350 18244
rect 15838 18232 15844 18244
rect 15896 18232 15902 18284
rect 17589 18275 17647 18281
rect 17589 18241 17601 18275
rect 17635 18272 17647 18275
rect 18156 18272 18184 18380
rect 19242 18368 19248 18380
rect 19300 18368 19306 18420
rect 20990 18368 20996 18420
rect 21048 18368 21054 18420
rect 24486 18408 24492 18420
rect 21192 18380 24492 18408
rect 17635 18244 18184 18272
rect 17635 18241 17647 18244
rect 17589 18235 17647 18241
rect 18414 18232 18420 18284
rect 18472 18232 18478 18284
rect 21192 18281 21220 18380
rect 24486 18368 24492 18380
rect 24544 18368 24550 18420
rect 21545 18343 21603 18349
rect 21545 18309 21557 18343
rect 21591 18340 21603 18343
rect 22094 18340 22100 18352
rect 21591 18312 22100 18340
rect 21591 18309 21603 18312
rect 21545 18303 21603 18309
rect 22094 18300 22100 18312
rect 22152 18300 22158 18352
rect 23385 18343 23443 18349
rect 23385 18309 23397 18343
rect 23431 18340 23443 18343
rect 23750 18340 23756 18352
rect 23431 18312 23756 18340
rect 23431 18309 23443 18312
rect 23385 18303 23443 18309
rect 23750 18300 23756 18312
rect 23808 18300 23814 18352
rect 19797 18275 19855 18281
rect 19797 18241 19809 18275
rect 19843 18272 19855 18275
rect 21177 18275 21235 18281
rect 19843 18244 20760 18272
rect 19843 18241 19855 18244
rect 19797 18235 19855 18241
rect 12544 18176 13032 18204
rect 8478 18068 8484 18080
rect 5643 18040 8484 18068
rect 8478 18028 8484 18040
rect 8536 18028 8542 18080
rect 9674 18028 9680 18080
rect 9732 18028 9738 18080
rect 12406 18040 12440 18080
rect 12434 18028 12440 18040
rect 12492 18028 12498 18080
rect 12802 18028 12808 18080
rect 12860 18068 12866 18080
rect 12897 18071 12955 18077
rect 12897 18068 12909 18071
rect 12860 18040 12909 18068
rect 12860 18028 12866 18040
rect 12897 18037 12909 18040
rect 12943 18037 12955 18071
rect 13004 18068 13032 18176
rect 13354 18164 13360 18216
rect 13412 18164 13418 18216
rect 13630 18164 13636 18216
rect 13688 18164 13694 18216
rect 15010 18164 15016 18216
rect 15068 18204 15074 18216
rect 15105 18207 15163 18213
rect 15105 18204 15117 18207
rect 15068 18176 15117 18204
rect 15068 18164 15074 18176
rect 15105 18173 15117 18176
rect 15151 18204 15163 18207
rect 17221 18207 17279 18213
rect 17221 18204 17233 18207
rect 15151 18176 17233 18204
rect 15151 18173 15163 18176
rect 15105 18167 15163 18173
rect 17221 18173 17233 18176
rect 17267 18173 17279 18207
rect 17221 18167 17279 18173
rect 17678 18164 17684 18216
rect 17736 18204 17742 18216
rect 18138 18204 18144 18216
rect 17736 18176 18144 18204
rect 17736 18164 17742 18176
rect 18138 18164 18144 18176
rect 18196 18164 18202 18216
rect 18432 18204 18460 18232
rect 20732 18216 20760 18244
rect 21177 18241 21189 18275
rect 21223 18241 21235 18275
rect 21177 18235 21235 18241
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18272 21327 18275
rect 21358 18272 21364 18284
rect 21315 18244 21364 18272
rect 21315 18241 21327 18244
rect 21269 18235 21327 18241
rect 21358 18232 21364 18244
rect 21416 18232 21422 18284
rect 21910 18232 21916 18284
rect 21968 18272 21974 18284
rect 21968 18244 22310 18272
rect 21968 18232 21974 18244
rect 18248 18176 18460 18204
rect 14826 18096 14832 18148
rect 14884 18096 14890 18148
rect 15470 18096 15476 18148
rect 15528 18136 15534 18148
rect 18248 18136 18276 18176
rect 19518 18164 19524 18216
rect 19576 18164 19582 18216
rect 20441 18207 20499 18213
rect 20441 18173 20453 18207
rect 20487 18173 20499 18207
rect 20441 18167 20499 18173
rect 20456 18136 20484 18167
rect 20714 18164 20720 18216
rect 20772 18164 20778 18216
rect 21637 18207 21695 18213
rect 21637 18173 21649 18207
rect 21683 18204 21695 18207
rect 22646 18204 22652 18216
rect 21683 18176 22652 18204
rect 21683 18173 21695 18176
rect 21637 18167 21695 18173
rect 22646 18164 22652 18176
rect 22704 18204 22710 18216
rect 22830 18204 22836 18216
rect 22704 18176 22836 18204
rect 22704 18164 22710 18176
rect 22830 18164 22836 18176
rect 22888 18164 22894 18216
rect 23661 18207 23719 18213
rect 23661 18173 23673 18207
rect 23707 18204 23719 18207
rect 24854 18204 24860 18216
rect 23707 18176 24860 18204
rect 23707 18173 23719 18176
rect 23661 18167 23719 18173
rect 24854 18164 24860 18176
rect 24912 18164 24918 18216
rect 15528 18108 18276 18136
rect 19720 18108 20484 18136
rect 15528 18096 15534 18108
rect 13446 18068 13452 18080
rect 13004 18040 13452 18068
rect 12897 18031 12955 18037
rect 13446 18028 13452 18040
rect 13504 18068 13510 18080
rect 14844 18068 14872 18096
rect 13504 18040 14872 18068
rect 13504 18028 13510 18040
rect 15286 18028 15292 18080
rect 15344 18028 15350 18080
rect 16574 18028 16580 18080
rect 16632 18068 16638 18080
rect 16669 18071 16727 18077
rect 16669 18068 16681 18071
rect 16632 18040 16681 18068
rect 16632 18028 16638 18040
rect 16669 18037 16681 18040
rect 16715 18037 16727 18071
rect 16669 18031 16727 18037
rect 18046 18028 18052 18080
rect 18104 18068 18110 18080
rect 19720 18068 19748 18108
rect 18104 18040 19748 18068
rect 18104 18028 18110 18040
rect 19886 18028 19892 18080
rect 19944 18028 19950 18080
rect 21913 18071 21971 18077
rect 21913 18037 21925 18071
rect 21959 18068 21971 18071
rect 22094 18068 22100 18080
rect 21959 18040 22100 18068
rect 21959 18037 21971 18040
rect 21913 18031 21971 18037
rect 22094 18028 22100 18040
rect 22152 18028 22158 18080
rect 1104 17978 26312 18000
rect 1104 17926 4101 17978
rect 4153 17926 4165 17978
rect 4217 17926 4229 17978
rect 4281 17926 4293 17978
rect 4345 17926 4357 17978
rect 4409 17926 10403 17978
rect 10455 17926 10467 17978
rect 10519 17926 10531 17978
rect 10583 17926 10595 17978
rect 10647 17926 10659 17978
rect 10711 17926 16705 17978
rect 16757 17926 16769 17978
rect 16821 17926 16833 17978
rect 16885 17926 16897 17978
rect 16949 17926 16961 17978
rect 17013 17926 23007 17978
rect 23059 17926 23071 17978
rect 23123 17926 23135 17978
rect 23187 17926 23199 17978
rect 23251 17926 23263 17978
rect 23315 17926 26312 17978
rect 1104 17904 26312 17926
rect 5721 17867 5779 17873
rect 5721 17833 5733 17867
rect 5767 17864 5779 17867
rect 6086 17864 6092 17876
rect 5767 17836 6092 17864
rect 5767 17833 5779 17836
rect 5721 17827 5779 17833
rect 6086 17824 6092 17836
rect 6144 17824 6150 17876
rect 6181 17867 6239 17873
rect 6181 17833 6193 17867
rect 6227 17864 6239 17867
rect 6454 17864 6460 17876
rect 6227 17836 6460 17864
rect 6227 17833 6239 17836
rect 6181 17827 6239 17833
rect 6454 17824 6460 17836
rect 6512 17824 6518 17876
rect 7653 17867 7711 17873
rect 7653 17833 7665 17867
rect 7699 17864 7711 17867
rect 8018 17864 8024 17876
rect 7699 17836 8024 17864
rect 7699 17833 7711 17836
rect 7653 17827 7711 17833
rect 8018 17824 8024 17836
rect 8076 17824 8082 17876
rect 9766 17824 9772 17876
rect 9824 17864 9830 17876
rect 9824 17836 12572 17864
rect 9824 17824 9830 17836
rect 6362 17756 6368 17808
rect 6420 17756 6426 17808
rect 6546 17756 6552 17808
rect 6604 17796 6610 17808
rect 6730 17796 6736 17808
rect 6604 17768 6736 17796
rect 6604 17756 6610 17768
rect 6730 17756 6736 17768
rect 6788 17796 6794 17808
rect 11333 17799 11391 17805
rect 6788 17768 8064 17796
rect 6788 17756 6794 17768
rect 5169 17731 5227 17737
rect 5169 17728 5181 17731
rect 3528 17700 5181 17728
rect 3528 17672 3556 17700
rect 5169 17697 5181 17700
rect 5215 17728 5227 17731
rect 5626 17728 5632 17740
rect 5215 17700 5632 17728
rect 5215 17697 5227 17700
rect 5169 17691 5227 17697
rect 5626 17688 5632 17700
rect 5684 17688 5690 17740
rect 6380 17728 6408 17756
rect 6825 17731 6883 17737
rect 5736 17700 6776 17728
rect 5736 17672 5764 17700
rect 3510 17620 3516 17672
rect 3568 17620 3574 17672
rect 4522 17620 4528 17672
rect 4580 17660 4586 17672
rect 4982 17660 4988 17672
rect 4580 17632 4988 17660
rect 4580 17620 4586 17632
rect 4982 17620 4988 17632
rect 5040 17620 5046 17672
rect 5258 17620 5264 17672
rect 5316 17620 5322 17672
rect 5350 17620 5356 17672
rect 5408 17620 5414 17672
rect 5445 17663 5503 17669
rect 5445 17629 5457 17663
rect 5491 17660 5503 17663
rect 5718 17660 5724 17672
rect 5491 17632 5724 17660
rect 5491 17629 5503 17632
rect 5445 17623 5503 17629
rect 5718 17620 5724 17632
rect 5776 17620 5782 17672
rect 5813 17663 5871 17669
rect 5813 17629 5825 17663
rect 5859 17629 5871 17663
rect 5813 17623 5871 17629
rect 5828 17592 5856 17623
rect 5994 17620 6000 17672
rect 6052 17660 6058 17672
rect 6270 17660 6276 17672
rect 6052 17632 6276 17660
rect 6052 17620 6058 17632
rect 6270 17620 6276 17632
rect 6328 17620 6334 17672
rect 6362 17620 6368 17672
rect 6420 17620 6426 17672
rect 6457 17663 6515 17669
rect 6457 17629 6469 17663
rect 6503 17629 6515 17663
rect 6457 17623 6515 17629
rect 6472 17592 6500 17623
rect 6546 17620 6552 17672
rect 6604 17620 6610 17672
rect 6641 17663 6699 17669
rect 6641 17629 6653 17663
rect 6687 17629 6699 17663
rect 6748 17660 6776 17700
rect 6825 17697 6837 17731
rect 6871 17728 6883 17731
rect 6871 17700 7972 17728
rect 6871 17697 6883 17700
rect 6825 17691 6883 17697
rect 7098 17660 7104 17672
rect 6748 17632 7104 17660
rect 6641 17623 6699 17629
rect 5184 17564 6500 17592
rect 5184 17536 5212 17564
rect 6656 17536 6684 17623
rect 7098 17620 7104 17632
rect 7156 17660 7162 17672
rect 7944 17669 7972 17700
rect 7193 17663 7251 17669
rect 7193 17660 7205 17663
rect 7156 17632 7205 17660
rect 7156 17620 7162 17632
rect 7193 17629 7205 17632
rect 7239 17629 7251 17663
rect 7193 17623 7251 17629
rect 7561 17663 7619 17669
rect 7561 17629 7573 17663
rect 7607 17660 7619 17663
rect 7837 17663 7895 17669
rect 7837 17660 7849 17663
rect 7607 17632 7849 17660
rect 7607 17629 7619 17632
rect 7561 17623 7619 17629
rect 7837 17629 7849 17632
rect 7883 17629 7895 17663
rect 7837 17623 7895 17629
rect 7929 17663 7987 17669
rect 7929 17629 7941 17663
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 8036 17601 8064 17768
rect 11333 17765 11345 17799
rect 11379 17796 11391 17799
rect 11790 17796 11796 17808
rect 11379 17768 11796 17796
rect 11379 17765 11391 17768
rect 11333 17759 11391 17765
rect 11790 17756 11796 17768
rect 11848 17756 11854 17808
rect 8110 17688 8116 17740
rect 8168 17728 8174 17740
rect 8297 17731 8355 17737
rect 8297 17728 8309 17731
rect 8168 17700 8309 17728
rect 8168 17688 8174 17700
rect 8297 17697 8309 17700
rect 8343 17697 8355 17731
rect 8297 17691 8355 17697
rect 12069 17731 12127 17737
rect 12069 17697 12081 17731
rect 12115 17728 12127 17731
rect 12250 17728 12256 17740
rect 12115 17700 12256 17728
rect 12115 17697 12127 17700
rect 12069 17691 12127 17697
rect 12250 17688 12256 17700
rect 12308 17688 12314 17740
rect 9674 17620 9680 17672
rect 9732 17620 9738 17672
rect 10870 17620 10876 17672
rect 10928 17620 10934 17672
rect 11149 17663 11207 17669
rect 11149 17629 11161 17663
rect 11195 17660 11207 17663
rect 12544 17660 12572 17836
rect 13630 17824 13636 17876
rect 13688 17824 13694 17876
rect 13740 17836 15424 17864
rect 13740 17796 13768 17836
rect 13280 17768 13768 17796
rect 15396 17796 15424 17836
rect 15838 17824 15844 17876
rect 15896 17824 15902 17876
rect 18322 17864 18328 17876
rect 16960 17836 18328 17864
rect 15933 17799 15991 17805
rect 15933 17796 15945 17799
rect 15396 17768 15945 17796
rect 12618 17688 12624 17740
rect 12676 17728 12682 17740
rect 13170 17728 13176 17740
rect 12676 17700 13176 17728
rect 12676 17688 12682 17700
rect 13170 17688 13176 17700
rect 13228 17688 13234 17740
rect 13280 17660 13308 17768
rect 15933 17765 15945 17768
rect 15979 17765 15991 17799
rect 15933 17759 15991 17765
rect 13354 17688 13360 17740
rect 13412 17728 13418 17740
rect 14093 17731 14151 17737
rect 14093 17728 14105 17731
rect 13412 17700 14105 17728
rect 13412 17688 13418 17700
rect 14093 17697 14105 17700
rect 14139 17728 14151 17731
rect 14734 17728 14740 17740
rect 14139 17700 14740 17728
rect 14139 17697 14151 17700
rect 14093 17691 14151 17697
rect 14734 17688 14740 17700
rect 14792 17728 14798 17740
rect 15010 17728 15016 17740
rect 14792 17700 15016 17728
rect 14792 17688 14798 17700
rect 15010 17688 15016 17700
rect 15068 17688 15074 17740
rect 16206 17688 16212 17740
rect 16264 17728 16270 17740
rect 16485 17731 16543 17737
rect 16485 17728 16497 17731
rect 16264 17700 16497 17728
rect 16264 17688 16270 17700
rect 16485 17697 16497 17700
rect 16531 17697 16543 17731
rect 16485 17691 16543 17697
rect 13449 17663 13507 17669
rect 13449 17660 13461 17663
rect 11195 17632 11468 17660
rect 12544 17632 12756 17660
rect 13280 17632 13461 17660
rect 11195 17629 11207 17632
rect 11149 17623 11207 17629
rect 7377 17595 7435 17601
rect 7377 17561 7389 17595
rect 7423 17592 7435 17595
rect 8021 17595 8079 17601
rect 7423 17564 7972 17592
rect 7423 17561 7435 17564
rect 7377 17555 7435 17561
rect 7944 17536 7972 17564
rect 8021 17561 8033 17595
rect 8067 17561 8079 17595
rect 8021 17555 8079 17561
rect 8159 17595 8217 17601
rect 8159 17561 8171 17595
rect 8205 17592 8217 17595
rect 9692 17592 9720 17620
rect 8205 17564 9720 17592
rect 8205 17561 8217 17564
rect 8159 17555 8217 17561
rect 5166 17484 5172 17536
rect 5224 17484 5230 17536
rect 6638 17484 6644 17536
rect 6696 17484 6702 17536
rect 7926 17484 7932 17536
rect 7984 17484 7990 17536
rect 10226 17484 10232 17536
rect 10284 17484 10290 17536
rect 11440 17533 11468 17632
rect 11793 17595 11851 17601
rect 11793 17561 11805 17595
rect 11839 17592 11851 17595
rect 12621 17595 12679 17601
rect 12621 17592 12633 17595
rect 11839 17564 12633 17592
rect 11839 17561 11851 17564
rect 11793 17555 11851 17561
rect 12621 17561 12633 17564
rect 12667 17561 12679 17595
rect 12621 17555 12679 17561
rect 11425 17527 11483 17533
rect 11425 17493 11437 17527
rect 11471 17493 11483 17527
rect 11425 17487 11483 17493
rect 11514 17484 11520 17536
rect 11572 17524 11578 17536
rect 11885 17527 11943 17533
rect 11885 17524 11897 17527
rect 11572 17496 11897 17524
rect 11572 17484 11578 17496
rect 11885 17493 11897 17496
rect 11931 17493 11943 17527
rect 12728 17524 12756 17632
rect 13449 17629 13461 17632
rect 13495 17629 13507 17663
rect 13449 17623 13507 17629
rect 13725 17663 13783 17669
rect 13725 17629 13737 17663
rect 13771 17660 13783 17663
rect 13998 17660 14004 17672
rect 13771 17632 14004 17660
rect 13771 17629 13783 17632
rect 13725 17623 13783 17629
rect 13998 17620 14004 17632
rect 14056 17620 14062 17672
rect 15470 17620 15476 17672
rect 15528 17620 15534 17672
rect 16301 17663 16359 17669
rect 16301 17629 16313 17663
rect 16347 17660 16359 17663
rect 16574 17660 16580 17672
rect 16347 17632 16580 17660
rect 16347 17629 16359 17632
rect 16301 17623 16359 17629
rect 16574 17620 16580 17632
rect 16632 17620 16638 17672
rect 14369 17595 14427 17601
rect 14369 17592 14381 17595
rect 13924 17564 14381 17592
rect 13446 17524 13452 17536
rect 12728 17496 13452 17524
rect 11885 17487 11943 17493
rect 13446 17484 13452 17496
rect 13504 17484 13510 17536
rect 13924 17533 13952 17564
rect 14369 17561 14381 17564
rect 14415 17561 14427 17595
rect 16960 17592 16988 17836
rect 18322 17824 18328 17836
rect 18380 17824 18386 17876
rect 18785 17867 18843 17873
rect 18785 17833 18797 17867
rect 18831 17864 18843 17867
rect 19518 17864 19524 17876
rect 18831 17836 19524 17864
rect 18831 17833 18843 17836
rect 18785 17827 18843 17833
rect 19518 17824 19524 17836
rect 19576 17824 19582 17876
rect 22097 17867 22155 17873
rect 22097 17833 22109 17867
rect 22143 17833 22155 17867
rect 22097 17827 22155 17833
rect 18874 17796 18880 17808
rect 17328 17768 18880 17796
rect 17034 17620 17040 17672
rect 17092 17620 17098 17672
rect 17185 17663 17243 17669
rect 17185 17629 17197 17663
rect 17231 17660 17243 17663
rect 17328 17660 17356 17768
rect 18874 17756 18880 17768
rect 18932 17756 18938 17808
rect 22112 17796 22140 17827
rect 22186 17824 22192 17876
rect 22244 17864 22250 17876
rect 22370 17864 22376 17876
rect 22244 17836 22376 17864
rect 22244 17824 22250 17836
rect 22370 17824 22376 17836
rect 22428 17824 22434 17876
rect 22646 17824 22652 17876
rect 22704 17864 22710 17876
rect 22704 17836 23152 17864
rect 22704 17824 22710 17836
rect 23017 17799 23075 17805
rect 22112 17768 22692 17796
rect 17402 17688 17408 17740
rect 17460 17728 17466 17740
rect 17865 17731 17923 17737
rect 17865 17728 17877 17731
rect 17460 17700 17877 17728
rect 17460 17688 17466 17700
rect 17865 17697 17877 17700
rect 17911 17697 17923 17731
rect 17865 17691 17923 17697
rect 18156 17700 19932 17728
rect 17231 17632 17356 17660
rect 17231 17629 17243 17632
rect 17185 17623 17243 17629
rect 17494 17620 17500 17672
rect 17552 17669 17558 17672
rect 17552 17660 17560 17669
rect 17552 17632 17597 17660
rect 17552 17623 17560 17632
rect 17552 17620 17558 17623
rect 18046 17620 18052 17672
rect 18104 17620 18110 17672
rect 18156 17669 18184 17700
rect 19904 17672 19932 17700
rect 20806 17688 20812 17740
rect 20864 17728 20870 17740
rect 22664 17728 22692 17768
rect 23017 17765 23029 17799
rect 23063 17765 23075 17799
rect 23124 17796 23152 17836
rect 23750 17824 23756 17876
rect 23808 17824 23814 17876
rect 23937 17867 23995 17873
rect 23937 17833 23949 17867
rect 23983 17864 23995 17867
rect 24118 17864 24124 17876
rect 23983 17836 24124 17864
rect 23983 17833 23995 17836
rect 23937 17827 23995 17833
rect 23952 17796 23980 17827
rect 24118 17824 24124 17836
rect 24176 17824 24182 17876
rect 23124 17768 23980 17796
rect 23017 17759 23075 17765
rect 23032 17728 23060 17759
rect 23109 17731 23167 17737
rect 23109 17728 23121 17731
rect 20864 17700 22416 17728
rect 22664 17700 22968 17728
rect 23032 17700 23121 17728
rect 20864 17688 20870 17700
rect 18141 17663 18199 17669
rect 18141 17629 18153 17663
rect 18187 17629 18199 17663
rect 18601 17663 18659 17669
rect 18601 17660 18613 17663
rect 18141 17623 18199 17629
rect 18524 17632 18613 17660
rect 17313 17595 17371 17601
rect 17313 17592 17325 17595
rect 16960 17564 17325 17592
rect 14369 17555 14427 17561
rect 17313 17561 17325 17564
rect 17359 17561 17371 17595
rect 17313 17555 17371 17561
rect 17405 17595 17463 17601
rect 17405 17561 17417 17595
rect 17451 17592 17463 17595
rect 18064 17592 18092 17620
rect 17451 17564 18092 17592
rect 17451 17561 17463 17564
rect 17405 17555 17463 17561
rect 13909 17527 13967 17533
rect 13909 17493 13921 17527
rect 13955 17493 13967 17527
rect 13909 17487 13967 17493
rect 16390 17484 16396 17536
rect 16448 17484 16454 17536
rect 17681 17527 17739 17533
rect 17681 17493 17693 17527
rect 17727 17524 17739 17527
rect 17954 17524 17960 17536
rect 17727 17496 17960 17524
rect 17727 17493 17739 17496
rect 17681 17487 17739 17493
rect 17954 17484 17960 17496
rect 18012 17484 18018 17536
rect 18049 17527 18107 17533
rect 18049 17493 18061 17527
rect 18095 17524 18107 17527
rect 18138 17524 18144 17536
rect 18095 17496 18144 17524
rect 18095 17493 18107 17496
rect 18049 17487 18107 17493
rect 18138 17484 18144 17496
rect 18196 17484 18202 17536
rect 18524 17533 18552 17632
rect 18601 17629 18613 17632
rect 18647 17629 18659 17663
rect 18601 17623 18659 17629
rect 19886 17620 19892 17672
rect 19944 17620 19950 17672
rect 21637 17663 21695 17669
rect 21637 17660 21649 17663
rect 20916 17632 21649 17660
rect 20916 17604 20944 17632
rect 21637 17629 21649 17632
rect 21683 17629 21695 17663
rect 21637 17623 21695 17629
rect 21726 17620 21732 17672
rect 21784 17660 21790 17672
rect 22005 17663 22063 17669
rect 22005 17660 22017 17663
rect 21784 17632 22017 17660
rect 21784 17620 21790 17632
rect 22005 17629 22017 17632
rect 22051 17629 22063 17663
rect 22005 17623 22063 17629
rect 22094 17620 22100 17672
rect 22152 17660 22158 17672
rect 22388 17669 22416 17700
rect 22281 17663 22339 17669
rect 22281 17660 22293 17663
rect 22152 17632 22293 17660
rect 22152 17620 22158 17632
rect 22281 17629 22293 17632
rect 22327 17629 22339 17663
rect 22281 17623 22339 17629
rect 22373 17663 22431 17669
rect 22373 17629 22385 17663
rect 22419 17629 22431 17663
rect 22373 17623 22431 17629
rect 20898 17552 20904 17604
rect 20956 17552 20962 17604
rect 22296 17592 22324 17623
rect 22462 17620 22468 17672
rect 22520 17620 22526 17672
rect 22646 17620 22652 17672
rect 22704 17620 22710 17672
rect 22830 17620 22836 17672
rect 22888 17620 22894 17672
rect 22940 17660 22968 17700
rect 23109 17697 23121 17700
rect 23155 17697 23167 17731
rect 25406 17728 25412 17740
rect 23109 17691 23167 17697
rect 23216 17700 25412 17728
rect 23216 17660 23244 17700
rect 25406 17688 25412 17700
rect 25464 17688 25470 17740
rect 22940 17632 23244 17660
rect 23382 17620 23388 17672
rect 23440 17620 23446 17672
rect 23845 17663 23903 17669
rect 23845 17660 23857 17663
rect 23676 17632 23857 17660
rect 22741 17595 22799 17601
rect 22741 17592 22753 17595
rect 22296 17564 22753 17592
rect 22741 17561 22753 17564
rect 22787 17592 22799 17595
rect 23400 17592 23428 17620
rect 22787 17564 23428 17592
rect 22787 17561 22799 17564
rect 22741 17555 22799 17561
rect 23676 17536 23704 17632
rect 23845 17629 23857 17632
rect 23891 17660 23903 17663
rect 23934 17660 23940 17672
rect 23891 17632 23940 17660
rect 23891 17629 23903 17632
rect 23845 17623 23903 17629
rect 23934 17620 23940 17632
rect 23992 17620 23998 17672
rect 18509 17527 18567 17533
rect 18509 17493 18521 17527
rect 18555 17493 18567 17527
rect 18509 17487 18567 17493
rect 21821 17527 21879 17533
rect 21821 17493 21833 17527
rect 21867 17524 21879 17527
rect 22186 17524 22192 17536
rect 21867 17496 22192 17524
rect 21867 17493 21879 17496
rect 21821 17487 21879 17493
rect 22186 17484 22192 17496
rect 22244 17484 22250 17536
rect 23658 17484 23664 17536
rect 23716 17484 23722 17536
rect 1104 17434 26472 17456
rect 1104 17382 7252 17434
rect 7304 17382 7316 17434
rect 7368 17382 7380 17434
rect 7432 17382 7444 17434
rect 7496 17382 7508 17434
rect 7560 17382 13554 17434
rect 13606 17382 13618 17434
rect 13670 17382 13682 17434
rect 13734 17382 13746 17434
rect 13798 17382 13810 17434
rect 13862 17382 19856 17434
rect 19908 17382 19920 17434
rect 19972 17382 19984 17434
rect 20036 17382 20048 17434
rect 20100 17382 20112 17434
rect 20164 17382 26158 17434
rect 26210 17382 26222 17434
rect 26274 17382 26286 17434
rect 26338 17382 26350 17434
rect 26402 17382 26414 17434
rect 26466 17382 26472 17434
rect 1104 17360 26472 17382
rect 4617 17323 4675 17329
rect 4617 17289 4629 17323
rect 4663 17320 4675 17323
rect 5350 17320 5356 17332
rect 4663 17292 5356 17320
rect 4663 17289 4675 17292
rect 4617 17283 4675 17289
rect 5350 17280 5356 17292
rect 5408 17280 5414 17332
rect 6362 17280 6368 17332
rect 6420 17320 6426 17332
rect 7101 17323 7159 17329
rect 7101 17320 7113 17323
rect 6420 17292 7113 17320
rect 6420 17280 6426 17292
rect 7101 17289 7113 17292
rect 7147 17289 7159 17323
rect 7101 17283 7159 17289
rect 9769 17323 9827 17329
rect 9769 17289 9781 17323
rect 9815 17320 9827 17323
rect 10226 17320 10232 17332
rect 9815 17292 10232 17320
rect 9815 17289 9827 17292
rect 9769 17283 9827 17289
rect 10226 17280 10232 17292
rect 10284 17280 10290 17332
rect 11057 17323 11115 17329
rect 11057 17289 11069 17323
rect 11103 17320 11115 17323
rect 11514 17320 11520 17332
rect 11103 17292 11520 17320
rect 11103 17289 11115 17292
rect 11057 17283 11115 17289
rect 3605 17255 3663 17261
rect 3605 17221 3617 17255
rect 3651 17252 3663 17255
rect 3651 17224 5212 17252
rect 3651 17221 3663 17224
rect 3605 17215 3663 17221
rect 3234 17184 3240 17196
rect 2990 17156 3240 17184
rect 3234 17144 3240 17156
rect 3292 17144 3298 17196
rect 4157 17187 4215 17193
rect 4157 17153 4169 17187
rect 4203 17184 4215 17187
rect 4449 17187 4507 17193
rect 4203 17156 4384 17184
rect 4203 17153 4215 17156
rect 4157 17147 4215 17153
rect 1578 17076 1584 17128
rect 1636 17076 1642 17128
rect 1854 17076 1860 17128
rect 1912 17076 1918 17128
rect 4249 17119 4307 17125
rect 4249 17085 4261 17119
rect 4295 17085 4307 17119
rect 4356 17116 4384 17156
rect 4449 17153 4461 17187
rect 4495 17184 4507 17187
rect 4540 17184 4568 17224
rect 5184 17196 5212 17224
rect 5368 17224 6408 17252
rect 5368 17196 5396 17224
rect 6380 17196 6408 17224
rect 6546 17212 6552 17264
rect 6604 17252 6610 17264
rect 6604 17224 7052 17252
rect 6604 17212 6610 17224
rect 7024 17196 7052 17224
rect 9582 17212 9588 17264
rect 9640 17252 9646 17264
rect 9677 17255 9735 17261
rect 9677 17252 9689 17255
rect 9640 17224 9689 17252
rect 9640 17212 9646 17224
rect 9677 17221 9689 17224
rect 9723 17252 9735 17255
rect 11072 17252 11100 17283
rect 11514 17280 11520 17292
rect 11572 17280 11578 17332
rect 12710 17280 12716 17332
rect 12768 17320 12774 17332
rect 12768 17292 12940 17320
rect 12768 17280 12774 17292
rect 11882 17252 11888 17264
rect 9723 17224 11100 17252
rect 11256 17224 11888 17252
rect 9723 17221 9735 17224
rect 9677 17215 9735 17221
rect 4495 17156 4568 17184
rect 4495 17153 4507 17156
rect 4449 17147 4507 17153
rect 4982 17144 4988 17196
rect 5040 17144 5046 17196
rect 5166 17144 5172 17196
rect 5224 17144 5230 17196
rect 5350 17144 5356 17196
rect 5408 17144 5414 17196
rect 5442 17144 5448 17196
rect 5500 17144 5506 17196
rect 5534 17144 5540 17196
rect 5592 17144 5598 17196
rect 6181 17187 6239 17193
rect 6181 17153 6193 17187
rect 6227 17184 6239 17187
rect 6270 17184 6276 17196
rect 6227 17156 6276 17184
rect 6227 17153 6239 17156
rect 6181 17147 6239 17153
rect 6270 17144 6276 17156
rect 6328 17144 6334 17196
rect 6362 17144 6368 17196
rect 6420 17144 6426 17196
rect 6825 17187 6883 17193
rect 6825 17153 6837 17187
rect 6871 17153 6883 17187
rect 6825 17147 6883 17153
rect 4706 17116 4712 17128
rect 4356 17088 4712 17116
rect 4249 17079 4307 17085
rect 4264 17048 4292 17079
rect 4706 17076 4712 17088
rect 4764 17116 4770 17128
rect 5460 17116 5488 17144
rect 4764 17088 5488 17116
rect 4764 17076 4770 17088
rect 5810 17076 5816 17128
rect 5868 17076 5874 17128
rect 6638 17116 6644 17128
rect 6104 17088 6644 17116
rect 4798 17048 4804 17060
rect 4264 17020 4804 17048
rect 4798 17008 4804 17020
rect 4856 17048 4862 17060
rect 5828 17048 5856 17076
rect 4856 17020 5856 17048
rect 4856 17008 4862 17020
rect 6104 16992 6132 17088
rect 6638 17076 6644 17088
rect 6696 17116 6702 17128
rect 6840 17116 6868 17147
rect 7006 17144 7012 17196
rect 7064 17144 7070 17196
rect 9030 17144 9036 17196
rect 9088 17144 9094 17196
rect 10321 17187 10379 17193
rect 10321 17153 10333 17187
rect 10367 17184 10379 17187
rect 10965 17187 11023 17193
rect 10367 17156 10640 17184
rect 10367 17153 10379 17156
rect 10321 17147 10379 17153
rect 6696 17088 6868 17116
rect 6696 17076 6702 17088
rect 7098 17076 7104 17128
rect 7156 17108 7162 17128
rect 7156 17080 7193 17108
rect 7156 17076 7162 17080
rect 9766 17076 9772 17128
rect 9824 17116 9830 17128
rect 9861 17119 9919 17125
rect 9861 17116 9873 17119
rect 9824 17088 9873 17116
rect 9824 17076 9830 17088
rect 9861 17085 9873 17088
rect 9907 17085 9919 17119
rect 9861 17079 9919 17085
rect 7101 17071 7159 17076
rect 6270 17008 6276 17060
rect 6328 17048 6334 17060
rect 6822 17048 6828 17060
rect 6328 17020 6828 17048
rect 6328 17008 6334 17020
rect 6822 17008 6828 17020
rect 6880 17048 6886 17060
rect 6917 17051 6975 17057
rect 6917 17048 6929 17051
rect 6880 17020 6929 17048
rect 6880 17008 6886 17020
rect 6917 17017 6929 17020
rect 6963 17017 6975 17051
rect 6917 17011 6975 17017
rect 8754 17008 8760 17060
rect 8812 17048 8818 17060
rect 10612 17057 10640 17156
rect 10965 17153 10977 17187
rect 11011 17184 11023 17187
rect 11146 17184 11152 17196
rect 11011 17156 11152 17184
rect 11011 17153 11023 17156
rect 10965 17147 11023 17153
rect 11146 17144 11152 17156
rect 11204 17144 11210 17196
rect 11256 17125 11284 17224
rect 11882 17212 11888 17224
rect 11940 17212 11946 17264
rect 12912 17196 12940 17292
rect 13170 17280 13176 17332
rect 13228 17320 13234 17332
rect 13265 17323 13323 17329
rect 13265 17320 13277 17323
rect 13228 17292 13277 17320
rect 13228 17280 13234 17292
rect 13265 17289 13277 17292
rect 13311 17289 13323 17323
rect 13265 17283 13323 17289
rect 13998 17280 14004 17332
rect 14056 17320 14062 17332
rect 14277 17323 14335 17329
rect 14277 17320 14289 17323
rect 14056 17292 14289 17320
rect 14056 17280 14062 17292
rect 14277 17289 14289 17292
rect 14323 17289 14335 17323
rect 14277 17283 14335 17289
rect 14737 17323 14795 17329
rect 14737 17289 14749 17323
rect 14783 17320 14795 17323
rect 15286 17320 15292 17332
rect 14783 17292 15292 17320
rect 14783 17289 14795 17292
rect 14737 17283 14795 17289
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 18417 17323 18475 17329
rect 18417 17289 18429 17323
rect 18463 17320 18475 17323
rect 18506 17320 18512 17332
rect 18463 17292 18512 17320
rect 18463 17289 18475 17292
rect 18417 17283 18475 17289
rect 14645 17255 14703 17261
rect 14645 17252 14657 17255
rect 14016 17224 14657 17252
rect 14016 17196 14044 17224
rect 14645 17221 14657 17224
rect 14691 17252 14703 17255
rect 15657 17255 15715 17261
rect 15657 17252 15669 17255
rect 14691 17224 15669 17252
rect 14691 17221 14703 17224
rect 14645 17215 14703 17221
rect 15657 17221 15669 17224
rect 15703 17252 15715 17255
rect 16390 17252 16396 17264
rect 15703 17224 16396 17252
rect 15703 17221 15715 17224
rect 15657 17215 15715 17221
rect 16390 17212 16396 17224
rect 16448 17212 16454 17264
rect 12894 17144 12900 17196
rect 12952 17144 12958 17196
rect 13998 17144 14004 17196
rect 14056 17144 14062 17196
rect 15565 17187 15623 17193
rect 15565 17153 15577 17187
rect 15611 17184 15623 17187
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 15611 17156 16681 17184
rect 15611 17153 15623 17156
rect 15565 17147 15623 17153
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 18432 17184 18460 17283
rect 18506 17280 18512 17292
rect 18564 17280 18570 17332
rect 18800 17292 20208 17320
rect 18800 17264 18828 17292
rect 18782 17212 18788 17264
rect 18840 17212 18846 17264
rect 20180 17261 20208 17292
rect 22462 17280 22468 17332
rect 22520 17320 22526 17332
rect 23293 17323 23351 17329
rect 23293 17320 23305 17323
rect 22520 17292 23305 17320
rect 22520 17280 22526 17292
rect 23293 17289 23305 17292
rect 23339 17289 23351 17323
rect 23293 17283 23351 17289
rect 19949 17255 20007 17261
rect 19949 17252 19961 17255
rect 19444 17224 19961 17252
rect 19444 17196 19472 17224
rect 19949 17221 19961 17224
rect 19995 17221 20007 17255
rect 19949 17215 20007 17221
rect 20165 17255 20223 17261
rect 20165 17221 20177 17255
rect 20211 17221 20223 17255
rect 20165 17215 20223 17221
rect 16669 17147 16727 17153
rect 16776 17156 18460 17184
rect 11241 17119 11299 17125
rect 11241 17085 11253 17119
rect 11287 17085 11299 17119
rect 11517 17119 11575 17125
rect 11517 17116 11529 17119
rect 11241 17079 11299 17085
rect 11440 17088 11529 17116
rect 9309 17051 9367 17057
rect 9309 17048 9321 17051
rect 8812 17020 9321 17048
rect 8812 17008 8818 17020
rect 9309 17017 9321 17020
rect 9355 17017 9367 17051
rect 9309 17011 9367 17017
rect 10597 17051 10655 17057
rect 10597 17017 10609 17051
rect 10643 17017 10655 17051
rect 11440 17048 11468 17088
rect 11517 17085 11529 17088
rect 11563 17085 11575 17119
rect 11517 17079 11575 17085
rect 11790 17076 11796 17128
rect 11848 17076 11854 17128
rect 11882 17076 11888 17128
rect 11940 17116 11946 17128
rect 13354 17116 13360 17128
rect 11940 17088 12940 17116
rect 11940 17076 11946 17088
rect 12912 17060 12940 17088
rect 13188 17088 13360 17116
rect 10597 17011 10655 17017
rect 10796 17020 11468 17048
rect 10796 16992 10824 17020
rect 4433 16983 4491 16989
rect 4433 16949 4445 16983
rect 4479 16980 4491 16983
rect 4982 16980 4988 16992
rect 4479 16952 4988 16980
rect 4479 16949 4491 16952
rect 4433 16943 4491 16949
rect 4982 16940 4988 16952
rect 5040 16940 5046 16992
rect 6086 16940 6092 16992
rect 6144 16940 6150 16992
rect 6178 16940 6184 16992
rect 6236 16940 6242 16992
rect 6454 16940 6460 16992
rect 6512 16980 6518 16992
rect 6733 16983 6791 16989
rect 6733 16980 6745 16983
rect 6512 16952 6745 16980
rect 6512 16940 6518 16952
rect 6733 16949 6745 16952
rect 6779 16949 6791 16983
rect 6733 16943 6791 16949
rect 8846 16940 8852 16992
rect 8904 16940 8910 16992
rect 10318 16940 10324 16992
rect 10376 16980 10382 16992
rect 10505 16983 10563 16989
rect 10505 16980 10517 16983
rect 10376 16952 10517 16980
rect 10376 16940 10382 16952
rect 10505 16949 10517 16952
rect 10551 16949 10563 16983
rect 10505 16943 10563 16949
rect 10778 16940 10784 16992
rect 10836 16940 10842 16992
rect 11440 16980 11468 17020
rect 12894 17008 12900 17060
rect 12952 17008 12958 17060
rect 13188 16980 13216 17088
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 13446 17076 13452 17128
rect 13504 17116 13510 17128
rect 14921 17119 14979 17125
rect 14921 17116 14933 17119
rect 13504 17088 14933 17116
rect 13504 17076 13510 17088
rect 14921 17085 14933 17088
rect 14967 17116 14979 17119
rect 14967 17088 15240 17116
rect 14967 17085 14979 17088
rect 14921 17079 14979 17085
rect 15102 17008 15108 17060
rect 15160 17008 15166 17060
rect 15212 17048 15240 17088
rect 15286 17076 15292 17128
rect 15344 17116 15350 17128
rect 15841 17119 15899 17125
rect 15841 17116 15853 17119
rect 15344 17088 15853 17116
rect 15344 17076 15350 17088
rect 15841 17085 15853 17088
rect 15887 17116 15899 17119
rect 16776 17116 16804 17156
rect 18506 17144 18512 17196
rect 18564 17144 18570 17196
rect 19058 17144 19064 17196
rect 19116 17144 19122 17196
rect 19426 17144 19432 17196
rect 19484 17144 19490 17196
rect 21358 17144 21364 17196
rect 21416 17144 21422 17196
rect 21542 17144 21548 17196
rect 21600 17144 21606 17196
rect 23934 17144 23940 17196
rect 23992 17184 23998 17196
rect 24762 17184 24768 17196
rect 23992 17156 24768 17184
rect 23992 17144 23998 17156
rect 24762 17144 24768 17156
rect 24820 17144 24826 17196
rect 25961 17187 26019 17193
rect 25961 17153 25973 17187
rect 26007 17153 26019 17187
rect 25961 17147 26019 17153
rect 15887 17088 16804 17116
rect 15887 17085 15899 17088
rect 15841 17079 15899 17085
rect 17034 17076 17040 17128
rect 17092 17116 17098 17128
rect 17221 17119 17279 17125
rect 17221 17116 17233 17119
rect 17092 17088 17233 17116
rect 17092 17076 17098 17088
rect 17221 17085 17233 17088
rect 17267 17085 17279 17119
rect 17862 17116 17868 17128
rect 17221 17079 17279 17085
rect 17328 17088 17868 17116
rect 17328 17048 17356 17088
rect 17862 17076 17868 17088
rect 17920 17076 17926 17128
rect 25976 17116 26004 17147
rect 26326 17116 26332 17128
rect 25976 17088 26332 17116
rect 26326 17076 26332 17088
rect 26384 17076 26390 17128
rect 15212 17020 17356 17048
rect 17402 17008 17408 17060
rect 17460 17048 17466 17060
rect 18785 17051 18843 17057
rect 18785 17048 18797 17051
rect 17460 17020 18797 17048
rect 17460 17008 17466 17020
rect 18785 17017 18797 17020
rect 18831 17017 18843 17051
rect 18785 17011 18843 17017
rect 11440 16952 13216 16980
rect 13262 16940 13268 16992
rect 13320 16980 13326 16992
rect 15120 16980 15148 17008
rect 13320 16952 15148 16980
rect 13320 16940 13326 16952
rect 15194 16940 15200 16992
rect 15252 16940 15258 16992
rect 19702 16940 19708 16992
rect 19760 16980 19766 16992
rect 19797 16983 19855 16989
rect 19797 16980 19809 16983
rect 19760 16952 19809 16980
rect 19760 16940 19766 16952
rect 19797 16949 19809 16952
rect 19843 16949 19855 16983
rect 19797 16943 19855 16949
rect 19978 16940 19984 16992
rect 20036 16940 20042 16992
rect 21545 16983 21603 16989
rect 21545 16949 21557 16983
rect 21591 16980 21603 16983
rect 22094 16980 22100 16992
rect 21591 16952 22100 16980
rect 21591 16949 21603 16952
rect 21545 16943 21603 16949
rect 22094 16940 22100 16952
rect 22152 16940 22158 16992
rect 25590 16940 25596 16992
rect 25648 16980 25654 16992
rect 25777 16983 25835 16989
rect 25777 16980 25789 16983
rect 25648 16952 25789 16980
rect 25648 16940 25654 16952
rect 25777 16949 25789 16952
rect 25823 16949 25835 16983
rect 25777 16943 25835 16949
rect 1104 16890 26312 16912
rect 1104 16838 4101 16890
rect 4153 16838 4165 16890
rect 4217 16838 4229 16890
rect 4281 16838 4293 16890
rect 4345 16838 4357 16890
rect 4409 16838 10403 16890
rect 10455 16838 10467 16890
rect 10519 16838 10531 16890
rect 10583 16838 10595 16890
rect 10647 16838 10659 16890
rect 10711 16838 16705 16890
rect 16757 16838 16769 16890
rect 16821 16838 16833 16890
rect 16885 16838 16897 16890
rect 16949 16838 16961 16890
rect 17013 16838 23007 16890
rect 23059 16838 23071 16890
rect 23123 16838 23135 16890
rect 23187 16838 23199 16890
rect 23251 16838 23263 16890
rect 23315 16838 26312 16890
rect 1104 16816 26312 16838
rect 1854 16736 1860 16788
rect 1912 16776 1918 16788
rect 2133 16779 2191 16785
rect 2133 16776 2145 16779
rect 1912 16748 2145 16776
rect 1912 16736 1918 16748
rect 2133 16745 2145 16748
rect 2179 16745 2191 16779
rect 2133 16739 2191 16745
rect 4801 16779 4859 16785
rect 4801 16745 4813 16779
rect 4847 16776 4859 16779
rect 5258 16776 5264 16788
rect 4847 16748 5264 16776
rect 4847 16745 4859 16748
rect 4801 16739 4859 16745
rect 5258 16736 5264 16748
rect 5316 16736 5322 16788
rect 6086 16736 6092 16788
rect 6144 16736 6150 16788
rect 10318 16736 10324 16788
rect 10376 16736 10382 16788
rect 10689 16779 10747 16785
rect 10689 16745 10701 16779
rect 10735 16776 10747 16779
rect 10870 16776 10876 16788
rect 10735 16748 10876 16776
rect 10735 16745 10747 16748
rect 10689 16739 10747 16745
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 11146 16736 11152 16788
rect 11204 16776 11210 16788
rect 11204 16748 12296 16776
rect 11204 16736 11210 16748
rect 4706 16668 4712 16720
rect 4764 16708 4770 16720
rect 5902 16708 5908 16720
rect 4764 16680 5908 16708
rect 4764 16668 4770 16680
rect 5902 16668 5908 16680
rect 5960 16668 5966 16720
rect 10336 16708 10364 16736
rect 10336 16680 10916 16708
rect 1486 16600 1492 16652
rect 1544 16600 1550 16652
rect 3326 16600 3332 16652
rect 3384 16600 3390 16652
rect 3973 16643 4031 16649
rect 3973 16609 3985 16643
rect 4019 16640 4031 16643
rect 4341 16643 4399 16649
rect 4019 16612 4292 16640
rect 4019 16609 4031 16612
rect 3973 16603 4031 16609
rect 2317 16575 2375 16581
rect 2317 16541 2329 16575
rect 2363 16541 2375 16575
rect 2317 16535 2375 16541
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16541 4215 16575
rect 4264 16572 4292 16612
rect 4341 16609 4353 16643
rect 4387 16640 4399 16643
rect 5350 16640 5356 16652
rect 4387 16612 5356 16640
rect 4387 16609 4399 16612
rect 4341 16603 4399 16609
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 5445 16643 5503 16649
rect 5445 16609 5457 16643
rect 5491 16640 5503 16643
rect 6454 16640 6460 16652
rect 5491 16612 6460 16640
rect 5491 16609 5503 16612
rect 5445 16603 5503 16609
rect 6454 16600 6460 16612
rect 6512 16600 6518 16652
rect 7009 16643 7067 16649
rect 7009 16609 7021 16643
rect 7055 16640 7067 16643
rect 7650 16640 7656 16652
rect 7055 16612 7656 16640
rect 7055 16609 7067 16612
rect 7009 16603 7067 16609
rect 7650 16600 7656 16612
rect 7708 16640 7714 16652
rect 8110 16640 8116 16652
rect 7708 16612 8116 16640
rect 7708 16600 7714 16612
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 10778 16600 10784 16652
rect 10836 16600 10842 16652
rect 10888 16640 10916 16680
rect 11057 16643 11115 16649
rect 11057 16640 11069 16643
rect 10888 16612 11069 16640
rect 11057 16609 11069 16612
rect 11103 16609 11115 16643
rect 11057 16603 11115 16609
rect 4264 16544 4660 16572
rect 4157 16535 4215 16541
rect 1765 16507 1823 16513
rect 1765 16473 1777 16507
rect 1811 16504 1823 16507
rect 2222 16504 2228 16516
rect 1811 16476 2228 16504
rect 1811 16473 1823 16476
rect 1765 16467 1823 16473
rect 2222 16464 2228 16476
rect 2280 16464 2286 16516
rect 2332 16436 2360 16535
rect 4172 16504 4200 16535
rect 4632 16516 4660 16544
rect 5166 16532 5172 16584
rect 5224 16532 5230 16584
rect 5534 16532 5540 16584
rect 5592 16572 5598 16584
rect 6089 16575 6147 16581
rect 6089 16572 6101 16575
rect 5592 16544 6101 16572
rect 5592 16532 5598 16544
rect 6089 16541 6101 16544
rect 6135 16541 6147 16575
rect 6089 16535 6147 16541
rect 6273 16575 6331 16581
rect 6273 16541 6285 16575
rect 6319 16572 6331 16575
rect 6362 16572 6368 16584
rect 6319 16544 6368 16572
rect 6319 16541 6331 16544
rect 6273 16535 6331 16541
rect 6362 16532 6368 16544
rect 6420 16532 6426 16584
rect 6546 16532 6552 16584
rect 6604 16532 6610 16584
rect 6730 16532 6736 16584
rect 6788 16532 6794 16584
rect 8573 16575 8631 16581
rect 8573 16541 8585 16575
rect 8619 16572 8631 16575
rect 8754 16572 8760 16584
rect 8619 16544 8760 16572
rect 8619 16541 8631 16544
rect 8573 16535 8631 16541
rect 8754 16532 8760 16544
rect 8812 16532 8818 16584
rect 8938 16532 8944 16584
rect 8996 16532 9002 16584
rect 12268 16572 12296 16748
rect 12434 16736 12440 16788
rect 12492 16776 12498 16788
rect 12529 16779 12587 16785
rect 12529 16776 12541 16779
rect 12492 16748 12541 16776
rect 12492 16736 12498 16748
rect 12529 16745 12541 16748
rect 12575 16745 12587 16779
rect 12529 16739 12587 16745
rect 12544 16640 12572 16739
rect 12894 16736 12900 16788
rect 12952 16776 12958 16788
rect 13262 16776 13268 16788
rect 12952 16748 13268 16776
rect 12952 16736 12958 16748
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 14645 16779 14703 16785
rect 14645 16745 14657 16779
rect 14691 16776 14703 16779
rect 15270 16779 15328 16785
rect 15270 16776 15282 16779
rect 14691 16748 15282 16776
rect 14691 16745 14703 16748
rect 14645 16739 14703 16745
rect 15270 16745 15282 16748
rect 15316 16745 15328 16779
rect 15270 16739 15328 16745
rect 16390 16736 16396 16788
rect 16448 16776 16454 16788
rect 18417 16779 18475 16785
rect 16448 16748 17356 16776
rect 16448 16736 16454 16748
rect 13173 16643 13231 16649
rect 13173 16640 13185 16643
rect 12544 16612 13185 16640
rect 13173 16609 13185 16612
rect 13219 16609 13231 16643
rect 13173 16603 13231 16609
rect 15010 16600 15016 16652
rect 15068 16600 15074 16652
rect 17328 16649 17356 16748
rect 18417 16745 18429 16779
rect 18463 16776 18475 16779
rect 18506 16776 18512 16788
rect 18463 16748 18512 16776
rect 18463 16745 18475 16748
rect 18417 16739 18475 16745
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 18601 16779 18659 16785
rect 18601 16745 18613 16779
rect 18647 16745 18659 16779
rect 18601 16739 18659 16745
rect 18616 16708 18644 16739
rect 19334 16736 19340 16788
rect 19392 16736 19398 16788
rect 23569 16779 23627 16785
rect 23569 16745 23581 16779
rect 23615 16776 23627 16779
rect 23934 16776 23940 16788
rect 23615 16748 23940 16776
rect 23615 16745 23627 16748
rect 23569 16739 23627 16745
rect 23934 16736 23940 16748
rect 23992 16736 23998 16788
rect 18432 16680 18644 16708
rect 18432 16652 18460 16680
rect 16761 16643 16819 16649
rect 16761 16609 16773 16643
rect 16807 16609 16819 16643
rect 16761 16603 16819 16609
rect 17313 16643 17371 16649
rect 17313 16609 17325 16643
rect 17359 16609 17371 16643
rect 17313 16603 17371 16609
rect 12621 16575 12679 16581
rect 12621 16572 12633 16575
rect 12268 16544 12633 16572
rect 12621 16541 12633 16544
rect 12667 16541 12679 16575
rect 12621 16535 12679 16541
rect 14461 16575 14519 16581
rect 14461 16541 14473 16575
rect 14507 16572 14519 16575
rect 14507 16544 14872 16572
rect 14507 16541 14519 16544
rect 14461 16535 14519 16541
rect 4433 16507 4491 16513
rect 4433 16504 4445 16507
rect 4172 16476 4445 16504
rect 4433 16473 4445 16476
rect 4479 16473 4491 16507
rect 4433 16467 4491 16473
rect 2685 16439 2743 16445
rect 2685 16436 2697 16439
rect 2332 16408 2697 16436
rect 2685 16405 2697 16408
rect 2731 16405 2743 16439
rect 2685 16399 2743 16405
rect 3050 16396 3056 16448
rect 3108 16396 3114 16448
rect 3145 16439 3203 16445
rect 3145 16405 3157 16439
rect 3191 16436 3203 16439
rect 3602 16436 3608 16448
rect 3191 16408 3608 16436
rect 3191 16405 3203 16408
rect 3145 16399 3203 16405
rect 3602 16396 3608 16408
rect 3660 16396 3666 16448
rect 4448 16436 4476 16467
rect 4614 16464 4620 16516
rect 4672 16464 4678 16516
rect 4706 16464 4712 16516
rect 4764 16464 4770 16516
rect 6914 16513 6920 16516
rect 6641 16507 6699 16513
rect 6641 16504 6653 16507
rect 5644 16476 6653 16504
rect 4724 16436 4752 16464
rect 5644 16448 5672 16476
rect 6641 16473 6653 16476
rect 6687 16473 6699 16507
rect 6641 16467 6699 16473
rect 6871 16507 6920 16513
rect 6871 16473 6883 16507
rect 6917 16473 6920 16507
rect 6871 16467 6920 16473
rect 6914 16464 6920 16467
rect 6972 16464 6978 16516
rect 9217 16507 9275 16513
rect 9217 16504 9229 16507
rect 8772 16476 9229 16504
rect 4448 16408 4752 16436
rect 5626 16396 5632 16448
rect 5684 16396 5690 16448
rect 5997 16439 6055 16445
rect 5997 16405 6009 16439
rect 6043 16436 6055 16439
rect 6270 16436 6276 16448
rect 6043 16408 6276 16436
rect 6043 16405 6055 16408
rect 5997 16399 6055 16405
rect 6270 16396 6276 16408
rect 6328 16396 6334 16448
rect 6362 16396 6368 16448
rect 6420 16396 6426 16448
rect 8772 16445 8800 16476
rect 9217 16473 9229 16476
rect 9263 16473 9275 16507
rect 9217 16467 9275 16473
rect 9490 16464 9496 16516
rect 9548 16504 9554 16516
rect 12710 16504 12716 16516
rect 9548 16476 9706 16504
rect 10520 16476 11546 16504
rect 12406 16476 12716 16504
rect 9548 16464 9554 16476
rect 8757 16439 8815 16445
rect 8757 16405 8769 16439
rect 8803 16405 8815 16439
rect 9600 16436 9628 16476
rect 10520 16436 10548 16476
rect 9600 16408 10548 16436
rect 11440 16436 11468 16476
rect 12066 16436 12072 16448
rect 11440 16408 12072 16436
rect 8757 16399 8815 16405
rect 12066 16396 12072 16408
rect 12124 16436 12130 16448
rect 12406 16436 12434 16476
rect 12710 16464 12716 16476
rect 12768 16464 12774 16516
rect 12124 16408 12434 16436
rect 12124 16396 12130 16408
rect 14734 16396 14740 16448
rect 14792 16396 14798 16448
rect 14844 16436 14872 16544
rect 14918 16532 14924 16584
rect 14976 16532 14982 16584
rect 16776 16572 16804 16603
rect 17402 16600 17408 16652
rect 17460 16600 17466 16652
rect 17770 16600 17776 16652
rect 17828 16640 17834 16652
rect 17828 16612 18368 16640
rect 17828 16600 17834 16612
rect 17034 16572 17040 16584
rect 16776 16544 17040 16572
rect 17034 16532 17040 16544
rect 17092 16572 17098 16584
rect 18233 16575 18291 16581
rect 18233 16572 18245 16575
rect 17092 16544 18245 16572
rect 17092 16532 17098 16544
rect 18233 16541 18245 16544
rect 18279 16541 18291 16575
rect 18340 16572 18368 16612
rect 18414 16600 18420 16652
rect 18472 16600 18478 16652
rect 18506 16600 18512 16652
rect 18564 16640 18570 16652
rect 19981 16643 20039 16649
rect 19981 16640 19993 16643
rect 18564 16612 19993 16640
rect 18564 16600 18570 16612
rect 19981 16609 19993 16612
rect 20027 16609 20039 16643
rect 19981 16603 20039 16609
rect 20898 16600 20904 16652
rect 20956 16640 20962 16652
rect 21177 16643 21235 16649
rect 21177 16640 21189 16643
rect 20956 16612 21189 16640
rect 20956 16600 20962 16612
rect 21177 16609 21189 16612
rect 21223 16609 21235 16643
rect 21177 16603 21235 16609
rect 22097 16643 22155 16649
rect 22097 16609 22109 16643
rect 22143 16640 22155 16643
rect 23474 16640 23480 16652
rect 22143 16612 23480 16640
rect 22143 16609 22155 16612
rect 22097 16603 22155 16609
rect 23474 16600 23480 16612
rect 23532 16600 23538 16652
rect 18524 16572 18552 16600
rect 18340 16544 18552 16572
rect 18233 16535 18291 16541
rect 18782 16532 18788 16584
rect 18840 16572 18846 16584
rect 18969 16575 19027 16581
rect 18969 16572 18981 16575
rect 18840 16544 18981 16572
rect 18840 16532 18846 16544
rect 18969 16541 18981 16544
rect 19015 16541 19027 16575
rect 18969 16535 19027 16541
rect 19334 16532 19340 16584
rect 19392 16572 19398 16584
rect 19797 16575 19855 16581
rect 19797 16572 19809 16575
rect 19392 16544 19809 16572
rect 19392 16532 19398 16544
rect 19797 16541 19809 16544
rect 19843 16541 19855 16575
rect 19797 16535 19855 16541
rect 20717 16575 20775 16581
rect 20717 16541 20729 16575
rect 20763 16541 20775 16575
rect 20717 16535 20775 16541
rect 15562 16464 15568 16516
rect 15620 16504 15626 16516
rect 17221 16507 17279 16513
rect 15620 16476 15778 16504
rect 15620 16464 15626 16476
rect 17221 16473 17233 16507
rect 17267 16504 17279 16507
rect 17681 16507 17739 16513
rect 17681 16504 17693 16507
rect 17267 16476 17693 16504
rect 17267 16473 17279 16476
rect 17221 16467 17279 16473
rect 17681 16473 17693 16476
rect 17727 16473 17739 16507
rect 17681 16467 17739 16473
rect 18601 16507 18659 16513
rect 18601 16473 18613 16507
rect 18647 16473 18659 16507
rect 18601 16467 18659 16473
rect 19613 16507 19671 16513
rect 19613 16473 19625 16507
rect 19659 16504 19671 16507
rect 19702 16504 19708 16516
rect 19659 16476 19708 16504
rect 19659 16473 19671 16476
rect 19613 16467 19671 16473
rect 16853 16439 16911 16445
rect 16853 16436 16865 16439
rect 14844 16408 16865 16436
rect 16853 16405 16865 16408
rect 16899 16405 16911 16439
rect 18616 16436 18644 16467
rect 19702 16464 19708 16476
rect 19760 16464 19766 16516
rect 19978 16464 19984 16516
rect 20036 16464 20042 16516
rect 20732 16504 20760 16535
rect 20806 16532 20812 16584
rect 20864 16572 20870 16584
rect 21085 16575 21143 16581
rect 21085 16572 21097 16575
rect 20864 16544 21097 16572
rect 20864 16532 20870 16544
rect 21085 16541 21097 16544
rect 21131 16541 21143 16575
rect 21085 16535 21143 16541
rect 20990 16504 20996 16516
rect 20732 16476 20996 16504
rect 20990 16464 20996 16476
rect 21048 16464 21054 16516
rect 18874 16436 18880 16448
rect 18616 16408 18880 16436
rect 16853 16399 16911 16405
rect 18874 16396 18880 16408
rect 18932 16436 18938 16448
rect 19996 16436 20024 16464
rect 18932 16408 20024 16436
rect 21100 16436 21128 16535
rect 21818 16532 21824 16584
rect 21876 16532 21882 16584
rect 23566 16504 23572 16516
rect 23322 16476 23572 16504
rect 23566 16464 23572 16476
rect 23624 16464 23630 16516
rect 23382 16436 23388 16448
rect 21100 16408 23388 16436
rect 18932 16396 18938 16408
rect 23382 16396 23388 16408
rect 23440 16396 23446 16448
rect 1104 16346 26472 16368
rect 1104 16294 7252 16346
rect 7304 16294 7316 16346
rect 7368 16294 7380 16346
rect 7432 16294 7444 16346
rect 7496 16294 7508 16346
rect 7560 16294 13554 16346
rect 13606 16294 13618 16346
rect 13670 16294 13682 16346
rect 13734 16294 13746 16346
rect 13798 16294 13810 16346
rect 13862 16294 19856 16346
rect 19908 16294 19920 16346
rect 19972 16294 19984 16346
rect 20036 16294 20048 16346
rect 20100 16294 20112 16346
rect 20164 16294 26158 16346
rect 26210 16294 26222 16346
rect 26274 16294 26286 16346
rect 26338 16294 26350 16346
rect 26402 16294 26414 16346
rect 26466 16294 26472 16346
rect 1104 16272 26472 16294
rect 5626 16192 5632 16244
rect 5684 16192 5690 16244
rect 6546 16192 6552 16244
rect 6604 16192 6610 16244
rect 6914 16192 6920 16244
rect 6972 16192 6978 16244
rect 7653 16235 7711 16241
rect 7653 16201 7665 16235
rect 7699 16201 7711 16235
rect 7653 16195 7711 16201
rect 2961 16167 3019 16173
rect 2961 16133 2973 16167
rect 3007 16164 3019 16167
rect 3510 16164 3516 16176
rect 3007 16136 3516 16164
rect 3007 16133 3019 16136
rect 2961 16127 3019 16133
rect 3510 16124 3516 16136
rect 3568 16124 3574 16176
rect 4982 16124 4988 16176
rect 5040 16164 5046 16176
rect 6564 16164 6592 16192
rect 7668 16164 7696 16195
rect 9490 16192 9496 16244
rect 9548 16232 9554 16244
rect 9548 16204 9812 16232
rect 9548 16192 9554 16204
rect 8938 16164 8944 16176
rect 5040 16136 5488 16164
rect 6564 16136 7696 16164
rect 8404 16136 8944 16164
rect 5040 16124 5046 16136
rect 2225 16099 2283 16105
rect 2225 16065 2237 16099
rect 2271 16065 2283 16099
rect 2225 16059 2283 16065
rect 2240 16028 2268 16059
rect 2498 16056 2504 16108
rect 2556 16056 2562 16108
rect 3050 16056 3056 16108
rect 3108 16096 3114 16108
rect 5166 16096 5172 16108
rect 3108 16068 5172 16096
rect 3108 16056 3114 16068
rect 3237 16031 3295 16037
rect 2240 16000 2636 16028
rect 2608 15969 2636 16000
rect 3237 15997 3249 16031
rect 3283 16028 3295 16031
rect 3326 16028 3332 16040
rect 3283 16000 3332 16028
rect 3283 15997 3295 16000
rect 3237 15991 3295 15997
rect 3326 15988 3332 16000
rect 3384 15988 3390 16040
rect 5092 16037 5120 16068
rect 5166 16056 5172 16068
rect 5224 16056 5230 16108
rect 5258 16056 5264 16108
rect 5316 16096 5322 16108
rect 5353 16099 5411 16105
rect 5353 16096 5365 16099
rect 5316 16068 5365 16096
rect 5316 16056 5322 16068
rect 5353 16065 5365 16068
rect 5399 16065 5411 16099
rect 5353 16059 5411 16065
rect 5460 16037 5488 16136
rect 5537 16099 5595 16105
rect 5537 16065 5549 16099
rect 5583 16096 5595 16099
rect 5718 16096 5724 16108
rect 5583 16068 5724 16096
rect 5583 16065 5595 16068
rect 5537 16059 5595 16065
rect 5718 16056 5724 16068
rect 5776 16056 5782 16108
rect 6270 16056 6276 16108
rect 6328 16096 6334 16108
rect 6730 16096 6736 16108
rect 6328 16068 6736 16096
rect 6328 16056 6334 16068
rect 6730 16056 6736 16068
rect 6788 16056 6794 16108
rect 6914 16056 6920 16108
rect 6972 16096 6978 16108
rect 8404 16105 8432 16136
rect 8938 16124 8944 16136
rect 8996 16124 9002 16176
rect 7561 16099 7619 16105
rect 7561 16096 7573 16099
rect 6972 16068 7573 16096
rect 6972 16056 6978 16068
rect 7561 16065 7573 16068
rect 7607 16096 7619 16099
rect 8389 16099 8447 16105
rect 7607 16068 8340 16096
rect 7607 16065 7619 16068
rect 7561 16059 7619 16065
rect 5077 16031 5135 16037
rect 5077 15997 5089 16031
rect 5123 15997 5135 16031
rect 5077 15991 5135 15997
rect 5445 16031 5503 16037
rect 5445 15997 5457 16031
rect 5491 16028 5503 16031
rect 7006 16028 7012 16040
rect 5491 16000 7012 16028
rect 5491 15997 5503 16000
rect 5445 15991 5503 15997
rect 2593 15963 2651 15969
rect 2593 15929 2605 15963
rect 2639 15929 2651 15963
rect 2593 15923 2651 15929
rect 2038 15852 2044 15904
rect 2096 15852 2102 15904
rect 2314 15852 2320 15904
rect 2372 15852 2378 15904
rect 5092 15892 5120 15991
rect 7006 15988 7012 16000
rect 7064 15988 7070 16040
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 7837 16031 7895 16037
rect 7837 16028 7849 16031
rect 7156 16000 7849 16028
rect 7156 15988 7162 16000
rect 7837 15997 7849 16000
rect 7883 15997 7895 16031
rect 7837 15991 7895 15997
rect 7929 16031 7987 16037
rect 7929 15997 7941 16031
rect 7975 15997 7987 16031
rect 7929 15991 7987 15997
rect 5169 15963 5227 15969
rect 5169 15929 5181 15963
rect 5215 15960 5227 15963
rect 5350 15960 5356 15972
rect 5215 15932 5356 15960
rect 5215 15929 5227 15932
rect 5169 15923 5227 15929
rect 5350 15920 5356 15932
rect 5408 15920 5414 15972
rect 6822 15920 6828 15972
rect 6880 15920 6886 15972
rect 6840 15892 6868 15920
rect 5092 15864 6868 15892
rect 7834 15852 7840 15904
rect 7892 15892 7898 15904
rect 7944 15892 7972 15991
rect 8018 15988 8024 16040
rect 8076 15988 8082 16040
rect 8113 16031 8171 16037
rect 8113 15997 8125 16031
rect 8159 15997 8171 16031
rect 8312 16028 8340 16068
rect 8389 16065 8401 16099
rect 8435 16065 8447 16099
rect 9784 16082 9812 16204
rect 10134 16192 10140 16244
rect 10192 16192 10198 16244
rect 14734 16192 14740 16244
rect 14792 16192 14798 16244
rect 16301 16235 16359 16241
rect 16301 16201 16313 16235
rect 16347 16232 16359 16235
rect 16942 16232 16948 16244
rect 16347 16204 16948 16232
rect 16347 16201 16359 16204
rect 16301 16195 16359 16201
rect 16942 16192 16948 16204
rect 17000 16192 17006 16244
rect 17034 16192 17040 16244
rect 17092 16192 17098 16244
rect 17218 16192 17224 16244
rect 17276 16232 17282 16244
rect 20809 16235 20867 16241
rect 17276 16204 19472 16232
rect 17276 16192 17282 16204
rect 10152 16096 10180 16192
rect 14752 16164 14780 16192
rect 14829 16167 14887 16173
rect 14829 16164 14841 16167
rect 14752 16136 14841 16164
rect 14829 16133 14841 16136
rect 14875 16133 14887 16167
rect 14829 16127 14887 16133
rect 15470 16124 15476 16176
rect 15528 16124 15534 16176
rect 16960 16164 16988 16192
rect 16868 16136 16988 16164
rect 10781 16099 10839 16105
rect 10781 16096 10793 16099
rect 10152 16068 10793 16096
rect 8389 16059 8447 16065
rect 10781 16065 10793 16068
rect 10827 16065 10839 16099
rect 10781 16059 10839 16065
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 16868 16105 16896 16136
rect 17052 16105 17080 16192
rect 19444 16176 19472 16204
rect 20809 16201 20821 16235
rect 20855 16232 20867 16235
rect 21358 16232 21364 16244
rect 20855 16204 21364 16232
rect 20855 16201 20867 16204
rect 20809 16195 20867 16201
rect 21358 16192 21364 16204
rect 21416 16192 21422 16244
rect 21818 16192 21824 16244
rect 21876 16232 21882 16244
rect 24854 16232 24860 16244
rect 21876 16204 24860 16232
rect 21876 16192 21882 16204
rect 24854 16192 24860 16204
rect 24912 16232 24918 16244
rect 24912 16204 25820 16232
rect 24912 16192 24918 16204
rect 17862 16124 17868 16176
rect 17920 16124 17926 16176
rect 19153 16131 19211 16137
rect 19153 16108 19165 16131
rect 19199 16108 19211 16131
rect 19426 16124 19432 16176
rect 19484 16164 19490 16176
rect 19613 16167 19671 16173
rect 19613 16164 19625 16167
rect 19484 16136 19625 16164
rect 19484 16124 19490 16136
rect 19613 16133 19625 16136
rect 19659 16164 19671 16167
rect 19659 16136 20668 16164
rect 19659 16133 19671 16136
rect 19613 16127 19671 16133
rect 20640 16108 20668 16136
rect 20714 16124 20720 16176
rect 20772 16164 20778 16176
rect 21836 16164 21864 16192
rect 20772 16136 21864 16164
rect 20772 16124 20778 16136
rect 16669 16099 16727 16105
rect 16669 16096 16681 16099
rect 16632 16068 16681 16096
rect 16632 16056 16638 16068
rect 16669 16065 16681 16068
rect 16715 16065 16727 16099
rect 16669 16059 16727 16065
rect 16817 16099 16896 16105
rect 16817 16065 16829 16099
rect 16863 16068 16896 16099
rect 16945 16099 17003 16105
rect 16863 16065 16875 16068
rect 16817 16059 16875 16065
rect 16945 16065 16957 16099
rect 16991 16065 17003 16099
rect 16945 16059 17003 16065
rect 17037 16099 17095 16105
rect 17037 16065 17049 16099
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 17175 16099 17233 16105
rect 17175 16065 17187 16099
rect 17221 16096 17233 16099
rect 17494 16096 17500 16108
rect 17221 16068 17500 16096
rect 17221 16065 17233 16068
rect 17175 16059 17233 16065
rect 13998 16028 14004 16040
rect 8312 16000 14004 16028
rect 8113 15991 8171 15997
rect 8128 15960 8156 15991
rect 13998 15988 14004 16000
rect 14056 15988 14062 16040
rect 14090 15988 14096 16040
rect 14148 16028 14154 16040
rect 14553 16031 14611 16037
rect 14553 16028 14565 16031
rect 14148 16000 14565 16028
rect 14148 15988 14154 16000
rect 14553 15997 14565 16000
rect 14599 15997 14611 16031
rect 14553 15991 14611 15997
rect 14826 15988 14832 16040
rect 14884 16028 14890 16040
rect 16960 16028 16988 16059
rect 17494 16056 17500 16068
rect 17552 16056 17558 16108
rect 18233 16099 18291 16105
rect 18233 16065 18245 16099
rect 18279 16065 18291 16099
rect 18233 16059 18291 16065
rect 14884 16000 16988 16028
rect 18248 16028 18276 16059
rect 18414 16056 18420 16108
rect 18472 16056 18478 16108
rect 18874 16056 18880 16108
rect 18932 16056 18938 16108
rect 19150 16056 19156 16108
rect 19208 16056 19214 16108
rect 19705 16099 19763 16105
rect 19705 16096 19717 16099
rect 19260 16068 19717 16096
rect 18782 16028 18788 16040
rect 18248 16000 18788 16028
rect 14884 15988 14890 16000
rect 8036 15932 8156 15960
rect 8036 15904 8064 15932
rect 18340 15904 18368 16000
rect 18782 15988 18788 16000
rect 18840 16028 18846 16040
rect 19260 16028 19288 16068
rect 19705 16065 19717 16068
rect 19751 16065 19763 16099
rect 19705 16059 19763 16065
rect 19889 16099 19947 16105
rect 19889 16065 19901 16099
rect 19935 16096 19947 16099
rect 19981 16099 20039 16105
rect 19981 16096 19993 16099
rect 19935 16068 19993 16096
rect 19935 16065 19947 16068
rect 19889 16059 19947 16065
rect 19981 16065 19993 16068
rect 20027 16065 20039 16099
rect 19981 16059 20039 16065
rect 20622 16056 20628 16108
rect 20680 16056 20686 16108
rect 20165 16031 20223 16037
rect 20165 16028 20177 16031
rect 18840 16000 19288 16028
rect 20088 16000 20177 16028
rect 18840 15988 18846 16000
rect 19153 15963 19211 15969
rect 19153 15929 19165 15963
rect 19199 15960 19211 15963
rect 19978 15960 19984 15972
rect 19199 15932 19984 15960
rect 19199 15929 19211 15932
rect 19153 15923 19211 15929
rect 19978 15920 19984 15932
rect 20036 15920 20042 15972
rect 7892 15864 7972 15892
rect 7892 15852 7898 15864
rect 8018 15852 8024 15904
rect 8076 15852 8082 15904
rect 8652 15895 8710 15901
rect 8652 15861 8664 15895
rect 8698 15892 8710 15895
rect 8846 15892 8852 15904
rect 8698 15864 8852 15892
rect 8698 15861 8710 15864
rect 8652 15855 8710 15861
rect 8846 15852 8852 15864
rect 8904 15852 8910 15904
rect 10226 15852 10232 15904
rect 10284 15852 10290 15904
rect 17310 15852 17316 15904
rect 17368 15852 17374 15904
rect 18322 15852 18328 15904
rect 18380 15852 18386 15904
rect 18690 15852 18696 15904
rect 18748 15892 18754 15904
rect 20088 15892 20116 16000
rect 20165 15997 20177 16000
rect 20211 15997 20223 16031
rect 20165 15991 20223 15997
rect 20438 15988 20444 16040
rect 20496 16028 20502 16040
rect 20824 16028 20852 16136
rect 21836 16105 21864 16136
rect 22094 16124 22100 16176
rect 22152 16124 22158 16176
rect 23382 16124 23388 16176
rect 23440 16164 23446 16176
rect 23845 16167 23903 16173
rect 23845 16164 23857 16167
rect 23440 16136 23857 16164
rect 23440 16124 23446 16136
rect 23845 16133 23857 16136
rect 23891 16133 23903 16167
rect 23845 16127 23903 16133
rect 25498 16124 25504 16176
rect 25556 16124 25562 16176
rect 20901 16099 20959 16105
rect 20901 16065 20913 16099
rect 20947 16065 20959 16099
rect 20901 16059 20959 16065
rect 21821 16099 21879 16105
rect 21821 16065 21833 16099
rect 21867 16065 21879 16099
rect 23566 16096 23572 16108
rect 23230 16082 23572 16096
rect 21821 16059 21879 16065
rect 23216 16068 23572 16082
rect 20496 16000 20852 16028
rect 20496 15988 20502 16000
rect 20916 15960 20944 16059
rect 21637 16031 21695 16037
rect 21637 15997 21649 16031
rect 21683 16028 21695 16031
rect 21726 16028 21732 16040
rect 21683 16000 21732 16028
rect 21683 15997 21695 16000
rect 21637 15991 21695 15997
rect 21726 15988 21732 16000
rect 21784 15988 21790 16040
rect 23216 16028 23244 16068
rect 23566 16056 23572 16068
rect 23624 16096 23630 16108
rect 24486 16096 24492 16108
rect 23624 16068 24492 16096
rect 23624 16056 23630 16068
rect 24486 16056 24492 16068
rect 24544 16056 24550 16108
rect 25792 16040 25820 16204
rect 21836 16000 23244 16028
rect 21836 15972 21864 16000
rect 25774 15988 25780 16040
rect 25832 15988 25838 16040
rect 20916 15932 21036 15960
rect 21008 15901 21036 15932
rect 21818 15920 21824 15972
rect 21876 15920 21882 15972
rect 18748 15864 20116 15892
rect 20993 15895 21051 15901
rect 18748 15852 18754 15864
rect 20993 15861 21005 15895
rect 21039 15892 21051 15895
rect 21358 15892 21364 15904
rect 21039 15864 21364 15892
rect 21039 15861 21051 15864
rect 20993 15855 21051 15861
rect 21358 15852 21364 15864
rect 21416 15852 21422 15904
rect 24026 15852 24032 15904
rect 24084 15852 24090 15904
rect 1104 15802 26312 15824
rect 1104 15750 4101 15802
rect 4153 15750 4165 15802
rect 4217 15750 4229 15802
rect 4281 15750 4293 15802
rect 4345 15750 4357 15802
rect 4409 15750 10403 15802
rect 10455 15750 10467 15802
rect 10519 15750 10531 15802
rect 10583 15750 10595 15802
rect 10647 15750 10659 15802
rect 10711 15750 16705 15802
rect 16757 15750 16769 15802
rect 16821 15750 16833 15802
rect 16885 15750 16897 15802
rect 16949 15750 16961 15802
rect 17013 15750 23007 15802
rect 23059 15750 23071 15802
rect 23123 15750 23135 15802
rect 23187 15750 23199 15802
rect 23251 15750 23263 15802
rect 23315 15750 26312 15802
rect 1104 15728 26312 15750
rect 1844 15691 1902 15697
rect 1844 15657 1856 15691
rect 1890 15688 1902 15691
rect 2314 15688 2320 15700
rect 1890 15660 2320 15688
rect 1890 15657 1902 15660
rect 1844 15651 1902 15657
rect 2314 15648 2320 15660
rect 2372 15648 2378 15700
rect 2498 15648 2504 15700
rect 2556 15688 2562 15700
rect 3789 15691 3847 15697
rect 3789 15688 3801 15691
rect 2556 15660 3801 15688
rect 2556 15648 2562 15660
rect 3789 15657 3801 15660
rect 3835 15657 3847 15691
rect 3789 15651 3847 15657
rect 4154 15648 4160 15700
rect 4212 15688 4218 15700
rect 4706 15688 4712 15700
rect 4212 15660 4712 15688
rect 4212 15648 4218 15660
rect 4706 15648 4712 15660
rect 4764 15688 4770 15700
rect 4764 15660 6500 15688
rect 4764 15648 4770 15660
rect 6472 15620 6500 15660
rect 6914 15648 6920 15700
rect 6972 15648 6978 15700
rect 7006 15648 7012 15700
rect 7064 15688 7070 15700
rect 8018 15688 8024 15700
rect 7064 15660 8024 15688
rect 7064 15648 7070 15660
rect 8018 15648 8024 15660
rect 8076 15648 8082 15700
rect 9030 15648 9036 15700
rect 9088 15688 9094 15700
rect 9217 15691 9275 15697
rect 9217 15688 9229 15691
rect 9088 15660 9229 15688
rect 9088 15648 9094 15660
rect 9217 15657 9229 15660
rect 9263 15657 9275 15691
rect 9217 15651 9275 15657
rect 10226 15648 10232 15700
rect 10284 15648 10290 15700
rect 10318 15648 10324 15700
rect 10376 15688 10382 15700
rect 11698 15688 11704 15700
rect 10376 15660 11704 15688
rect 10376 15648 10382 15660
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 17037 15691 17095 15697
rect 17037 15657 17049 15691
rect 17083 15688 17095 15691
rect 18138 15688 18144 15700
rect 17083 15660 18144 15688
rect 17083 15657 17095 15660
rect 17037 15651 17095 15657
rect 18138 15648 18144 15660
rect 18196 15648 18202 15700
rect 19058 15648 19064 15700
rect 19116 15688 19122 15700
rect 19245 15691 19303 15697
rect 19245 15688 19257 15691
rect 19116 15660 19257 15688
rect 19116 15648 19122 15660
rect 19245 15657 19257 15660
rect 19291 15657 19303 15691
rect 19245 15651 19303 15657
rect 19334 15648 19340 15700
rect 19392 15648 19398 15700
rect 21726 15648 21732 15700
rect 21784 15688 21790 15700
rect 21784 15660 22094 15688
rect 21784 15648 21790 15660
rect 4264 15592 4752 15620
rect 6472 15592 7144 15620
rect 1578 15512 1584 15564
rect 1636 15552 1642 15564
rect 2590 15552 2596 15564
rect 1636 15524 2596 15552
rect 1636 15512 1642 15524
rect 2590 15512 2596 15524
rect 2648 15552 2654 15564
rect 4264 15552 4292 15592
rect 4724 15564 4752 15592
rect 2648 15524 4292 15552
rect 4341 15555 4399 15561
rect 2648 15512 2654 15524
rect 4341 15521 4353 15555
rect 4387 15521 4399 15555
rect 4341 15515 4399 15521
rect 3234 15484 3240 15496
rect 2990 15456 3240 15484
rect 3234 15444 3240 15456
rect 3292 15444 3298 15496
rect 3326 15444 3332 15496
rect 3384 15484 3390 15496
rect 4062 15484 4068 15496
rect 3384 15456 4068 15484
rect 3384 15444 3390 15456
rect 4062 15444 4068 15456
rect 4120 15484 4126 15496
rect 4356 15484 4384 15515
rect 4706 15512 4712 15564
rect 4764 15552 4770 15564
rect 5169 15555 5227 15561
rect 5169 15552 5181 15555
rect 4764 15524 5181 15552
rect 4764 15512 4770 15524
rect 5169 15521 5181 15524
rect 5215 15552 5227 15555
rect 7116 15552 7144 15592
rect 7834 15552 7840 15564
rect 5215 15524 7052 15552
rect 7116 15524 7840 15552
rect 5215 15521 5227 15524
rect 5169 15515 5227 15521
rect 4120 15456 4384 15484
rect 4120 15444 4126 15456
rect 4982 15444 4988 15496
rect 5040 15444 5046 15496
rect 7024 15493 7052 15524
rect 7834 15512 7840 15524
rect 7892 15512 7898 15564
rect 9398 15512 9404 15564
rect 9456 15552 9462 15564
rect 9769 15555 9827 15561
rect 9769 15552 9781 15555
rect 9456 15524 9781 15552
rect 9456 15512 9462 15524
rect 9769 15521 9781 15524
rect 9815 15521 9827 15555
rect 9769 15515 9827 15521
rect 7009 15487 7067 15493
rect 7009 15453 7021 15487
rect 7055 15453 7067 15487
rect 9490 15484 9496 15496
rect 8418 15456 9496 15484
rect 7009 15447 7067 15453
rect 3602 15376 3608 15428
rect 3660 15416 3666 15428
rect 5000 15416 5028 15444
rect 3660 15388 5028 15416
rect 5445 15419 5503 15425
rect 3660 15376 3666 15388
rect 4172 15357 4200 15388
rect 5445 15385 5457 15419
rect 5491 15385 5503 15419
rect 5445 15379 5503 15385
rect 4157 15351 4215 15357
rect 4157 15317 4169 15351
rect 4203 15317 4215 15351
rect 4157 15311 4215 15317
rect 4249 15351 4307 15357
rect 4249 15317 4261 15351
rect 4295 15348 4307 15351
rect 4338 15348 4344 15360
rect 4295 15320 4344 15348
rect 4295 15317 4307 15320
rect 4249 15311 4307 15317
rect 4338 15308 4344 15320
rect 4396 15348 4402 15360
rect 4614 15348 4620 15360
rect 4396 15320 4620 15348
rect 4396 15308 4402 15320
rect 4614 15308 4620 15320
rect 4672 15308 4678 15360
rect 5460 15348 5488 15379
rect 5902 15376 5908 15428
rect 5960 15376 5966 15428
rect 6362 15348 6368 15360
rect 5460 15320 6368 15348
rect 6362 15308 6368 15320
rect 6420 15308 6426 15360
rect 7024 15348 7052 15447
rect 9490 15444 9496 15456
rect 9548 15444 9554 15496
rect 9585 15487 9643 15493
rect 9585 15453 9597 15487
rect 9631 15484 9643 15487
rect 10244 15484 10272 15648
rect 17221 15623 17279 15629
rect 17221 15589 17233 15623
rect 17267 15620 17279 15623
rect 19352 15620 19380 15648
rect 17267 15592 19380 15620
rect 17267 15589 17279 15592
rect 17221 15583 17279 15589
rect 19978 15580 19984 15632
rect 20036 15620 20042 15632
rect 20036 15592 20392 15620
rect 20036 15580 20042 15592
rect 12342 15512 12348 15564
rect 12400 15552 12406 15564
rect 12529 15555 12587 15561
rect 12529 15552 12541 15555
rect 12400 15524 12541 15552
rect 12400 15512 12406 15524
rect 12529 15521 12541 15524
rect 12575 15521 12587 15555
rect 12529 15515 12587 15521
rect 17770 15512 17776 15564
rect 17828 15552 17834 15564
rect 18414 15552 18420 15564
rect 17828 15524 18420 15552
rect 17828 15512 17834 15524
rect 18414 15512 18420 15524
rect 18472 15552 18478 15564
rect 19521 15555 19579 15561
rect 19521 15552 19533 15555
rect 18472 15524 19533 15552
rect 18472 15512 18478 15524
rect 19521 15521 19533 15524
rect 19567 15521 19579 15555
rect 19521 15515 19579 15521
rect 20364 15496 20392 15592
rect 9631 15456 10272 15484
rect 9631 15453 9643 15456
rect 9585 15447 9643 15453
rect 11422 15444 11428 15496
rect 11480 15484 11486 15496
rect 11517 15487 11575 15493
rect 11517 15484 11529 15487
rect 11480 15456 11529 15484
rect 11480 15444 11486 15456
rect 11517 15453 11529 15456
rect 11563 15453 11575 15487
rect 11517 15447 11575 15453
rect 11885 15487 11943 15493
rect 11885 15453 11897 15487
rect 11931 15484 11943 15487
rect 14093 15487 14151 15493
rect 11931 15456 12020 15484
rect 11931 15453 11943 15456
rect 11885 15447 11943 15453
rect 7190 15376 7196 15428
rect 7248 15416 7254 15428
rect 7285 15419 7343 15425
rect 7285 15416 7297 15419
rect 7248 15388 7297 15416
rect 7248 15376 7254 15388
rect 7285 15385 7297 15388
rect 7331 15385 7343 15419
rect 7285 15379 7343 15385
rect 8018 15348 8024 15360
rect 7024 15320 8024 15348
rect 8018 15308 8024 15320
rect 8076 15308 8082 15360
rect 8757 15351 8815 15357
rect 8757 15317 8769 15351
rect 8803 15348 8815 15351
rect 8846 15348 8852 15360
rect 8803 15320 8852 15348
rect 8803 15317 8815 15320
rect 8757 15311 8815 15317
rect 8846 15308 8852 15320
rect 8904 15348 8910 15360
rect 9582 15348 9588 15360
rect 8904 15320 9588 15348
rect 8904 15308 8910 15320
rect 9582 15308 9588 15320
rect 9640 15348 9646 15360
rect 9677 15351 9735 15357
rect 9677 15348 9689 15351
rect 9640 15320 9689 15348
rect 9640 15308 9646 15320
rect 9677 15317 9689 15320
rect 9723 15317 9735 15351
rect 9677 15311 9735 15317
rect 11330 15308 11336 15360
rect 11388 15308 11394 15360
rect 11698 15308 11704 15360
rect 11756 15308 11762 15360
rect 11992 15357 12020 15456
rect 14093 15453 14105 15487
rect 14139 15484 14151 15487
rect 14182 15484 14188 15496
rect 14139 15456 14188 15484
rect 14139 15453 14151 15456
rect 14093 15447 14151 15453
rect 14182 15444 14188 15456
rect 14240 15444 14246 15496
rect 16206 15444 16212 15496
rect 16264 15484 16270 15496
rect 17313 15487 17371 15493
rect 17313 15484 17325 15487
rect 16264 15456 17325 15484
rect 16264 15444 16270 15456
rect 17313 15453 17325 15456
rect 17359 15453 17371 15487
rect 17313 15447 17371 15453
rect 18506 15444 18512 15496
rect 18564 15444 18570 15496
rect 18601 15487 18659 15493
rect 18601 15453 18613 15487
rect 18647 15484 18659 15487
rect 18690 15484 18696 15496
rect 18647 15456 18696 15484
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 18690 15444 18696 15456
rect 18748 15444 18754 15496
rect 18874 15444 18880 15496
rect 18932 15484 18938 15496
rect 19061 15487 19119 15493
rect 18932 15456 18977 15484
rect 18932 15444 18938 15456
rect 19061 15453 19073 15487
rect 19107 15484 19119 15487
rect 19334 15484 19340 15496
rect 19107 15456 19340 15484
rect 19107 15453 19119 15456
rect 19061 15447 19119 15453
rect 19334 15444 19340 15456
rect 19392 15444 19398 15496
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 20165 15487 20223 15493
rect 20165 15484 20177 15487
rect 19484 15456 20177 15484
rect 19484 15444 19490 15456
rect 20165 15453 20177 15456
rect 20211 15453 20223 15487
rect 20165 15447 20223 15453
rect 20346 15444 20352 15496
rect 20404 15444 20410 15496
rect 20438 15444 20444 15496
rect 20496 15444 20502 15496
rect 21818 15444 21824 15496
rect 21876 15444 21882 15496
rect 12437 15419 12495 15425
rect 12437 15385 12449 15419
rect 12483 15416 12495 15419
rect 12526 15416 12532 15428
rect 12483 15388 12532 15416
rect 12483 15385 12495 15388
rect 12437 15379 12495 15385
rect 12526 15376 12532 15388
rect 12584 15376 12590 15428
rect 16853 15419 16911 15425
rect 16853 15385 16865 15419
rect 16899 15416 16911 15419
rect 16899 15388 17632 15416
rect 16899 15385 16911 15388
rect 16853 15379 16911 15385
rect 11977 15351 12035 15357
rect 11977 15317 11989 15351
rect 12023 15317 12035 15351
rect 11977 15311 12035 15317
rect 12345 15351 12403 15357
rect 12345 15317 12357 15351
rect 12391 15348 12403 15351
rect 13446 15348 13452 15360
rect 12391 15320 13452 15348
rect 12391 15317 12403 15320
rect 12345 15311 12403 15317
rect 13446 15308 13452 15320
rect 13504 15308 13510 15360
rect 14277 15351 14335 15357
rect 14277 15317 14289 15351
rect 14323 15348 14335 15351
rect 14366 15348 14372 15360
rect 14323 15320 14372 15348
rect 14323 15317 14335 15320
rect 14277 15311 14335 15317
rect 14366 15308 14372 15320
rect 14424 15308 14430 15360
rect 17063 15351 17121 15357
rect 17063 15317 17075 15351
rect 17109 15348 17121 15351
rect 17218 15348 17224 15360
rect 17109 15320 17224 15348
rect 17109 15317 17121 15320
rect 17063 15311 17121 15317
rect 17218 15308 17224 15320
rect 17276 15308 17282 15360
rect 17604 15348 17632 15388
rect 17678 15376 17684 15428
rect 17736 15376 17742 15428
rect 17862 15376 17868 15428
rect 17920 15376 17926 15428
rect 19150 15416 19156 15428
rect 18248 15388 19156 15416
rect 18248 15360 18276 15388
rect 19150 15376 19156 15388
rect 19208 15416 19214 15428
rect 19981 15419 20039 15425
rect 19981 15416 19993 15419
rect 19208 15388 19993 15416
rect 19208 15376 19214 15388
rect 19981 15385 19993 15388
rect 20027 15385 20039 15419
rect 19981 15379 20039 15385
rect 20714 15376 20720 15428
rect 20772 15376 20778 15428
rect 22066 15416 22094 15660
rect 22554 15648 22560 15700
rect 22612 15688 22618 15700
rect 23201 15691 23259 15697
rect 23201 15688 23213 15691
rect 22612 15660 23213 15688
rect 22612 15648 22618 15660
rect 23201 15657 23213 15660
rect 23247 15657 23259 15691
rect 23201 15651 23259 15657
rect 23474 15648 23480 15700
rect 23532 15648 23538 15700
rect 24026 15648 24032 15700
rect 24084 15648 24090 15700
rect 22278 15512 22284 15564
rect 22336 15512 22342 15564
rect 24044 15552 24072 15648
rect 24397 15555 24455 15561
rect 24397 15552 24409 15555
rect 24044 15524 24409 15552
rect 24397 15521 24409 15524
rect 24443 15521 24455 15555
rect 24397 15515 24455 15521
rect 23661 15487 23719 15493
rect 23661 15484 23673 15487
rect 23400 15456 23673 15484
rect 23017 15419 23075 15425
rect 23017 15416 23029 15419
rect 22066 15388 23029 15416
rect 18230 15348 18236 15360
rect 17604 15320 18236 15348
rect 18230 15308 18236 15320
rect 18288 15308 18294 15360
rect 18322 15308 18328 15360
rect 18380 15348 18386 15360
rect 19426 15348 19432 15360
rect 18380 15320 19432 15348
rect 18380 15308 18386 15320
rect 19426 15308 19432 15320
rect 19484 15308 19490 15360
rect 19610 15308 19616 15360
rect 19668 15348 19674 15360
rect 22204 15357 22232 15388
rect 23017 15385 23029 15388
rect 23063 15385 23075 15419
rect 23017 15379 23075 15385
rect 20257 15351 20315 15357
rect 20257 15348 20269 15351
rect 19668 15320 20269 15348
rect 19668 15308 19674 15320
rect 20257 15317 20269 15320
rect 20303 15317 20315 15351
rect 20257 15311 20315 15317
rect 22189 15351 22247 15357
rect 22189 15317 22201 15351
rect 22235 15317 22247 15351
rect 22189 15311 22247 15317
rect 22922 15308 22928 15360
rect 22980 15308 22986 15360
rect 23106 15308 23112 15360
rect 23164 15348 23170 15360
rect 23400 15357 23428 15456
rect 23661 15453 23673 15456
rect 23707 15453 23719 15487
rect 23661 15447 23719 15453
rect 23217 15351 23275 15357
rect 23217 15348 23229 15351
rect 23164 15320 23229 15348
rect 23164 15308 23170 15320
rect 23217 15317 23229 15320
rect 23263 15317 23275 15351
rect 23217 15311 23275 15317
rect 23385 15351 23443 15357
rect 23385 15317 23397 15351
rect 23431 15317 23443 15351
rect 23385 15311 23443 15317
rect 25041 15351 25099 15357
rect 25041 15317 25053 15351
rect 25087 15348 25099 15351
rect 25222 15348 25228 15360
rect 25087 15320 25228 15348
rect 25087 15317 25099 15320
rect 25041 15311 25099 15317
rect 25222 15308 25228 15320
rect 25280 15308 25286 15360
rect 1104 15258 26472 15280
rect 1104 15206 7252 15258
rect 7304 15206 7316 15258
rect 7368 15206 7380 15258
rect 7432 15206 7444 15258
rect 7496 15206 7508 15258
rect 7560 15206 13554 15258
rect 13606 15206 13618 15258
rect 13670 15206 13682 15258
rect 13734 15206 13746 15258
rect 13798 15206 13810 15258
rect 13862 15206 19856 15258
rect 19908 15206 19920 15258
rect 19972 15206 19984 15258
rect 20036 15206 20048 15258
rect 20100 15206 20112 15258
rect 20164 15206 26158 15258
rect 26210 15206 26222 15258
rect 26274 15206 26286 15258
rect 26338 15206 26350 15258
rect 26402 15206 26414 15258
rect 26466 15206 26472 15258
rect 1104 15184 26472 15206
rect 2038 15104 2044 15156
rect 2096 15104 2102 15156
rect 4062 15104 4068 15156
rect 4120 15104 4126 15156
rect 4154 15104 4160 15156
rect 4212 15104 4218 15156
rect 5718 15104 5724 15156
rect 5776 15144 5782 15156
rect 6454 15144 6460 15156
rect 5776 15116 6460 15144
rect 5776 15104 5782 15116
rect 6454 15104 6460 15116
rect 6512 15104 6518 15156
rect 6917 15147 6975 15153
rect 6917 15113 6929 15147
rect 6963 15144 6975 15147
rect 7098 15144 7104 15156
rect 6963 15116 7104 15144
rect 6963 15113 6975 15116
rect 6917 15107 6975 15113
rect 7098 15104 7104 15116
rect 7156 15104 7162 15156
rect 10965 15147 11023 15153
rect 10965 15113 10977 15147
rect 11011 15144 11023 15147
rect 11333 15147 11391 15153
rect 11011 15116 11284 15144
rect 11011 15113 11023 15116
rect 10965 15107 11023 15113
rect 1857 15079 1915 15085
rect 1857 15045 1869 15079
rect 1903 15076 1915 15079
rect 2056 15076 2084 15104
rect 3234 15076 3240 15088
rect 1903 15048 2084 15076
rect 3082 15048 3240 15076
rect 1903 15045 1915 15048
rect 1857 15039 1915 15045
rect 3234 15036 3240 15048
rect 3292 15036 3298 15088
rect 4080 15076 4108 15104
rect 4080 15048 4292 15076
rect 1578 14968 1584 15020
rect 1636 14968 1642 15020
rect 3510 14968 3516 15020
rect 3568 15008 3574 15020
rect 3605 15011 3663 15017
rect 3605 15008 3617 15011
rect 3568 14980 3617 15008
rect 3568 14968 3574 14980
rect 3605 14977 3617 14980
rect 3651 15008 3663 15011
rect 3970 15008 3976 15020
rect 3651 14980 3976 15008
rect 3651 14977 3663 14980
rect 3605 14971 3663 14977
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 4065 15011 4123 15017
rect 4065 14977 4077 15011
rect 4111 14977 4123 15011
rect 4065 14971 4123 14977
rect 4080 14872 4108 14971
rect 4264 14949 4292 15048
rect 7374 15036 7380 15088
rect 7432 15076 7438 15088
rect 7469 15079 7527 15085
rect 7469 15076 7481 15079
rect 7432 15048 7481 15076
rect 7432 15036 7438 15048
rect 7469 15045 7481 15048
rect 7515 15076 7527 15079
rect 7650 15076 7656 15088
rect 7515 15048 7656 15076
rect 7515 15045 7527 15048
rect 7469 15039 7527 15045
rect 7650 15036 7656 15048
rect 7708 15036 7714 15088
rect 6178 14968 6184 15020
rect 6236 15008 6242 15020
rect 6365 15011 6423 15017
rect 6365 15008 6377 15011
rect 6236 14980 6377 15008
rect 6236 14968 6242 14980
rect 6365 14977 6377 14980
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 4249 14943 4307 14949
rect 4249 14909 4261 14943
rect 4295 14909 4307 14943
rect 6380 14940 6408 14971
rect 6546 14968 6552 15020
rect 6604 15008 6610 15020
rect 6641 15011 6699 15017
rect 6641 15008 6653 15011
rect 6604 14980 6653 15008
rect 6604 14968 6610 14980
rect 6641 14977 6653 14980
rect 6687 14977 6699 15011
rect 6641 14971 6699 14977
rect 7190 14968 7196 15020
rect 7248 14968 7254 15020
rect 8846 14968 8852 15020
rect 8904 14968 8910 15020
rect 11256 15008 11284 15116
rect 11333 15113 11345 15147
rect 11379 15144 11391 15147
rect 11422 15144 11428 15156
rect 11379 15116 11428 15144
rect 11379 15113 11391 15116
rect 11333 15107 11391 15113
rect 11422 15104 11428 15116
rect 11480 15104 11486 15156
rect 27062 15144 27068 15156
rect 11532 15116 14136 15144
rect 11422 15008 11428 15020
rect 10796 14980 11100 15008
rect 11256 14980 11428 15008
rect 6730 14940 6736 14952
rect 6380 14912 6736 14940
rect 4249 14903 4307 14909
rect 6730 14900 6736 14912
rect 6788 14900 6794 14952
rect 10796 14949 10824 14980
rect 11072 14952 11100 14980
rect 11422 14968 11428 14980
rect 11480 14968 11486 15020
rect 11532 15017 11560 15116
rect 14108 15088 14136 15116
rect 15304 15116 27068 15144
rect 11698 15036 11704 15088
rect 11756 15076 11762 15088
rect 11793 15079 11851 15085
rect 11793 15076 11805 15079
rect 11756 15048 11805 15076
rect 11756 15036 11762 15048
rect 11793 15045 11805 15048
rect 11839 15045 11851 15079
rect 11793 15039 11851 15045
rect 12066 15036 12072 15088
rect 12124 15076 12130 15088
rect 12250 15076 12256 15088
rect 12124 15048 12256 15076
rect 12124 15036 12130 15048
rect 12250 15036 12256 15048
rect 12308 15036 12314 15088
rect 14090 15036 14096 15088
rect 14148 15036 14154 15088
rect 15304 15085 15332 15116
rect 27062 15104 27068 15116
rect 27120 15104 27126 15156
rect 15289 15079 15347 15085
rect 15289 15045 15301 15079
rect 15335 15045 15347 15079
rect 15289 15039 15347 15045
rect 16758 15036 16764 15088
rect 16816 15076 16822 15088
rect 17770 15076 17776 15088
rect 16816 15048 17776 15076
rect 16816 15036 16822 15048
rect 17770 15036 17776 15048
rect 17828 15076 17834 15088
rect 17925 15079 17983 15085
rect 17925 15076 17937 15079
rect 17828 15048 17937 15076
rect 17828 15036 17834 15048
rect 17925 15045 17937 15048
rect 17971 15045 17983 15079
rect 17925 15039 17983 15045
rect 18141 15079 18199 15085
rect 18141 15045 18153 15079
rect 18187 15076 18199 15079
rect 18230 15076 18236 15088
rect 18187 15048 18236 15076
rect 18187 15045 18199 15048
rect 18141 15039 18199 15045
rect 18230 15036 18236 15048
rect 18288 15036 18294 15088
rect 19150 15036 19156 15088
rect 19208 15036 19214 15088
rect 21192 15048 21588 15076
rect 11517 15011 11575 15017
rect 11517 14977 11529 15011
rect 11563 14977 11575 15011
rect 11517 14971 11575 14977
rect 7101 14943 7159 14949
rect 7101 14909 7113 14943
rect 7147 14909 7159 14943
rect 7101 14903 7159 14909
rect 7561 14943 7619 14949
rect 7561 14909 7573 14943
rect 7607 14940 7619 14943
rect 8205 14943 8263 14949
rect 8205 14940 8217 14943
rect 7607 14912 8217 14940
rect 7607 14909 7619 14912
rect 7561 14903 7619 14909
rect 8205 14909 8217 14912
rect 8251 14909 8263 14943
rect 8205 14903 8263 14909
rect 10781 14943 10839 14949
rect 10781 14909 10793 14943
rect 10827 14909 10839 14943
rect 10781 14903 10839 14909
rect 10873 14943 10931 14949
rect 10873 14909 10885 14943
rect 10919 14909 10931 14943
rect 10873 14903 10931 14909
rect 4338 14872 4344 14884
rect 4080 14844 4344 14872
rect 4338 14832 4344 14844
rect 4396 14872 4402 14884
rect 4798 14872 4804 14884
rect 4396 14844 4804 14872
rect 4396 14832 4402 14844
rect 4798 14832 4804 14844
rect 4856 14832 4862 14884
rect 6641 14875 6699 14881
rect 6641 14841 6653 14875
rect 6687 14872 6699 14875
rect 7116 14872 7144 14903
rect 6687 14844 7144 14872
rect 10888 14872 10916 14903
rect 11054 14900 11060 14952
rect 11112 14900 11118 14952
rect 11238 14900 11244 14952
rect 11296 14940 11302 14952
rect 11532 14940 11560 14971
rect 12802 14940 12808 14952
rect 11296 14912 11560 14940
rect 11624 14912 12808 14940
rect 11296 14900 11302 14912
rect 11624 14872 11652 14912
rect 12802 14900 12808 14912
rect 12860 14900 12866 14952
rect 18138 14900 18144 14952
rect 18196 14900 18202 14952
rect 18248 14949 18276 15036
rect 19981 15011 20039 15017
rect 19981 14977 19993 15011
rect 20027 15008 20039 15011
rect 20438 15008 20444 15020
rect 20027 14980 20444 15008
rect 20027 14977 20039 14980
rect 19981 14971 20039 14977
rect 20438 14968 20444 14980
rect 20496 14968 20502 15020
rect 20990 14968 20996 15020
rect 21048 14968 21054 15020
rect 21192 15017 21220 15048
rect 21560 15020 21588 15048
rect 24486 15036 24492 15088
rect 24544 15036 24550 15088
rect 25222 15036 25228 15088
rect 25280 15076 25286 15088
rect 25501 15079 25559 15085
rect 25501 15076 25513 15079
rect 25280 15048 25513 15076
rect 25280 15036 25286 15048
rect 25501 15045 25513 15048
rect 25547 15045 25559 15079
rect 25501 15039 25559 15045
rect 21177 15011 21235 15017
rect 21177 14977 21189 15011
rect 21223 14977 21235 15011
rect 21177 14971 21235 14977
rect 21358 14968 21364 15020
rect 21416 14968 21422 15020
rect 21542 14968 21548 15020
rect 21600 15008 21606 15020
rect 23106 15008 23112 15020
rect 21600 14980 23112 15008
rect 21600 14968 21606 14980
rect 23106 14968 23112 14980
rect 23164 14968 23170 15020
rect 25774 14968 25780 15020
rect 25832 14968 25838 15020
rect 18233 14943 18291 14949
rect 18233 14909 18245 14943
rect 18279 14909 18291 14943
rect 18233 14903 18291 14909
rect 19702 14900 19708 14952
rect 19760 14900 19766 14952
rect 21008 14940 21036 14968
rect 21008 14912 21220 14940
rect 10888 14844 11652 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 17678 14832 17684 14884
rect 17736 14832 17742 14884
rect 3694 14764 3700 14816
rect 3752 14764 3758 14816
rect 4890 14764 4896 14816
rect 4948 14804 4954 14816
rect 9582 14804 9588 14816
rect 4948 14776 9588 14804
rect 4948 14764 4954 14776
rect 9582 14764 9588 14776
rect 9640 14804 9646 14816
rect 10134 14804 10140 14816
rect 9640 14776 10140 14804
rect 9640 14764 9646 14776
rect 10134 14764 10140 14776
rect 10192 14764 10198 14816
rect 13265 14807 13323 14813
rect 13265 14773 13277 14807
rect 13311 14804 13323 14807
rect 13446 14804 13452 14816
rect 13311 14776 13452 14804
rect 13311 14773 13323 14776
rect 13265 14767 13323 14773
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 13998 14764 14004 14816
rect 14056 14804 14062 14816
rect 17586 14804 17592 14816
rect 14056 14776 17592 14804
rect 14056 14764 14062 14776
rect 17586 14764 17592 14776
rect 17644 14764 17650 14816
rect 17696 14804 17724 14832
rect 17773 14807 17831 14813
rect 17773 14804 17785 14807
rect 17696 14776 17785 14804
rect 17773 14773 17785 14776
rect 17819 14773 17831 14807
rect 17773 14767 17831 14773
rect 17957 14807 18015 14813
rect 17957 14773 17969 14807
rect 18003 14804 18015 14807
rect 18156 14804 18184 14900
rect 20714 14832 20720 14884
rect 20772 14872 20778 14884
rect 20993 14875 21051 14881
rect 20993 14872 21005 14875
rect 20772 14844 21005 14872
rect 20772 14832 20778 14844
rect 20993 14841 21005 14844
rect 21039 14841 21051 14875
rect 21192 14872 21220 14912
rect 21266 14900 21272 14952
rect 21324 14900 21330 14952
rect 21453 14943 21511 14949
rect 21453 14909 21465 14943
rect 21499 14909 21511 14943
rect 21453 14903 21511 14909
rect 21468 14872 21496 14903
rect 21192 14844 21496 14872
rect 20993 14835 21051 14841
rect 18003 14776 18184 14804
rect 18003 14773 18015 14776
rect 17957 14767 18015 14773
rect 23382 14764 23388 14816
rect 23440 14804 23446 14816
rect 24029 14807 24087 14813
rect 24029 14804 24041 14807
rect 23440 14776 24041 14804
rect 23440 14764 23446 14776
rect 24029 14773 24041 14776
rect 24075 14804 24087 14807
rect 25038 14804 25044 14816
rect 24075 14776 25044 14804
rect 24075 14773 24087 14776
rect 24029 14767 24087 14773
rect 25038 14764 25044 14776
rect 25096 14764 25102 14816
rect 1104 14714 26312 14736
rect 1104 14662 4101 14714
rect 4153 14662 4165 14714
rect 4217 14662 4229 14714
rect 4281 14662 4293 14714
rect 4345 14662 4357 14714
rect 4409 14662 10403 14714
rect 10455 14662 10467 14714
rect 10519 14662 10531 14714
rect 10583 14662 10595 14714
rect 10647 14662 10659 14714
rect 10711 14662 16705 14714
rect 16757 14662 16769 14714
rect 16821 14662 16833 14714
rect 16885 14662 16897 14714
rect 16949 14662 16961 14714
rect 17013 14662 23007 14714
rect 23059 14662 23071 14714
rect 23123 14662 23135 14714
rect 23187 14662 23199 14714
rect 23251 14662 23263 14714
rect 23315 14662 26312 14714
rect 1104 14640 26312 14662
rect 3694 14560 3700 14612
rect 3752 14560 3758 14612
rect 6454 14560 6460 14612
rect 6512 14560 6518 14612
rect 6917 14603 6975 14609
rect 6917 14569 6929 14603
rect 6963 14600 6975 14603
rect 7190 14600 7196 14612
rect 6963 14572 7196 14600
rect 6963 14569 6975 14572
rect 6917 14563 6975 14569
rect 7190 14560 7196 14572
rect 7248 14560 7254 14612
rect 11054 14600 11060 14612
rect 10796 14572 11060 14600
rect 3142 14356 3148 14408
rect 3200 14356 3206 14408
rect 3513 14399 3571 14405
rect 3513 14365 3525 14399
rect 3559 14396 3571 14399
rect 3712 14396 3740 14560
rect 6472 14532 6500 14560
rect 6472 14504 6684 14532
rect 3970 14424 3976 14476
rect 4028 14464 4034 14476
rect 6546 14464 6552 14476
rect 4028 14436 6552 14464
rect 4028 14424 4034 14436
rect 5920 14408 5948 14436
rect 6546 14424 6552 14436
rect 6604 14424 6610 14476
rect 6656 14473 6684 14504
rect 7742 14492 7748 14544
rect 7800 14532 7806 14544
rect 8110 14532 8116 14544
rect 7800 14504 8116 14532
rect 7800 14492 7806 14504
rect 8110 14492 8116 14504
rect 8168 14532 8174 14544
rect 10686 14532 10692 14544
rect 8168 14504 10692 14532
rect 8168 14492 8174 14504
rect 10686 14492 10692 14504
rect 10744 14492 10750 14544
rect 6641 14467 6699 14473
rect 6641 14433 6653 14467
rect 6687 14433 6699 14467
rect 6641 14427 6699 14433
rect 6730 14424 6736 14476
rect 6788 14424 6794 14476
rect 10594 14464 10600 14476
rect 9692 14436 10600 14464
rect 3559 14368 3740 14396
rect 3559 14365 3571 14368
rect 3513 14359 3571 14365
rect 5902 14356 5908 14408
rect 5960 14356 5966 14408
rect 6457 14399 6515 14405
rect 6457 14365 6469 14399
rect 6503 14396 6515 14399
rect 6914 14396 6920 14408
rect 6503 14368 6920 14396
rect 6503 14365 6515 14368
rect 6457 14359 6515 14365
rect 6914 14356 6920 14368
rect 6972 14396 6978 14408
rect 9692 14405 9720 14436
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 10796 14473 10824 14572
rect 11054 14560 11060 14572
rect 11112 14600 11118 14612
rect 11112 14572 12388 14600
rect 11112 14560 11118 14572
rect 12360 14544 12388 14572
rect 18138 14560 18144 14612
rect 18196 14600 18202 14612
rect 19610 14600 19616 14612
rect 18196 14572 19616 14600
rect 18196 14560 18202 14572
rect 12342 14492 12348 14544
rect 12400 14492 12406 14544
rect 18693 14535 18751 14541
rect 18693 14501 18705 14535
rect 18739 14501 18751 14535
rect 18693 14495 18751 14501
rect 18785 14535 18843 14541
rect 18785 14501 18797 14535
rect 18831 14532 18843 14535
rect 18874 14532 18880 14544
rect 18831 14504 18880 14532
rect 18831 14501 18843 14504
rect 18785 14495 18843 14501
rect 10781 14467 10839 14473
rect 10781 14433 10793 14467
rect 10827 14433 10839 14467
rect 10781 14427 10839 14433
rect 11241 14467 11299 14473
rect 11241 14433 11253 14467
rect 11287 14464 11299 14467
rect 11330 14464 11336 14476
rect 11287 14436 11336 14464
rect 11287 14433 11299 14436
rect 11241 14427 11299 14433
rect 11330 14424 11336 14436
rect 11388 14424 11394 14476
rect 11606 14424 11612 14476
rect 11664 14464 11670 14476
rect 11974 14464 11980 14476
rect 11664 14436 11980 14464
rect 11664 14424 11670 14436
rect 11974 14424 11980 14436
rect 12032 14464 12038 14476
rect 12713 14467 12771 14473
rect 12713 14464 12725 14467
rect 12032 14436 12725 14464
rect 12032 14424 12038 14436
rect 12713 14433 12725 14436
rect 12759 14433 12771 14467
rect 12713 14427 12771 14433
rect 14366 14424 14372 14476
rect 14424 14424 14430 14476
rect 18230 14424 18236 14476
rect 18288 14464 18294 14476
rect 18325 14467 18383 14473
rect 18325 14464 18337 14467
rect 18288 14436 18337 14464
rect 18288 14424 18294 14436
rect 18325 14433 18337 14436
rect 18371 14433 18383 14467
rect 18708 14464 18736 14495
rect 18874 14492 18880 14504
rect 18932 14492 18938 14544
rect 19352 14541 19380 14572
rect 19610 14560 19616 14572
rect 19668 14560 19674 14612
rect 19797 14603 19855 14609
rect 19797 14569 19809 14603
rect 19843 14569 19855 14603
rect 19797 14563 19855 14569
rect 22741 14603 22799 14609
rect 22741 14569 22753 14603
rect 22787 14600 22799 14603
rect 23290 14600 23296 14612
rect 22787 14572 23296 14600
rect 22787 14569 22799 14572
rect 22741 14563 22799 14569
rect 19337 14535 19395 14541
rect 19337 14501 19349 14535
rect 19383 14501 19395 14535
rect 19337 14495 19395 14501
rect 19426 14492 19432 14544
rect 19484 14532 19490 14544
rect 19812 14532 19840 14563
rect 23290 14560 23296 14572
rect 23348 14560 23354 14612
rect 23382 14560 23388 14612
rect 23440 14560 23446 14612
rect 24578 14560 24584 14612
rect 24636 14560 24642 14612
rect 22925 14535 22983 14541
rect 22925 14532 22937 14535
rect 19484 14504 19840 14532
rect 22020 14504 22937 14532
rect 19484 14492 19490 14504
rect 19889 14467 19947 14473
rect 19889 14464 19901 14467
rect 18708 14436 19901 14464
rect 18325 14427 18383 14433
rect 19889 14433 19901 14436
rect 19935 14464 19947 14467
rect 20346 14464 20352 14476
rect 19935 14436 20352 14464
rect 19935 14433 19947 14436
rect 19889 14427 19947 14433
rect 7929 14399 7987 14405
rect 7929 14396 7941 14399
rect 6972 14368 7941 14396
rect 6972 14356 6978 14368
rect 7929 14365 7941 14368
rect 7975 14365 7987 14399
rect 7929 14359 7987 14365
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14396 8171 14399
rect 9677 14399 9735 14405
rect 8159 14368 8248 14396
rect 8159 14365 8171 14368
rect 8113 14359 8171 14365
rect 2777 14331 2835 14337
rect 2777 14297 2789 14331
rect 2823 14328 2835 14331
rect 2823 14300 3188 14328
rect 2823 14297 2835 14300
rect 2777 14291 2835 14297
rect 3160 14272 3188 14300
rect 8220 14272 8248 14368
rect 9677 14365 9689 14399
rect 9723 14365 9735 14399
rect 9677 14359 9735 14365
rect 10045 14399 10103 14405
rect 10045 14365 10057 14399
rect 10091 14365 10103 14399
rect 10045 14359 10103 14365
rect 9950 14328 9956 14340
rect 8312 14300 9956 14328
rect 8312 14272 8340 14300
rect 9950 14288 9956 14300
rect 10008 14288 10014 14340
rect 3142 14220 3148 14272
rect 3200 14220 3206 14272
rect 3326 14220 3332 14272
rect 3384 14220 3390 14272
rect 8202 14220 8208 14272
rect 8260 14220 8266 14272
rect 8294 14220 8300 14272
rect 8352 14220 8358 14272
rect 9306 14220 9312 14272
rect 9364 14260 9370 14272
rect 9493 14263 9551 14269
rect 9493 14260 9505 14263
rect 9364 14232 9505 14260
rect 9364 14220 9370 14232
rect 9493 14229 9505 14232
rect 9539 14229 9551 14263
rect 9493 14223 9551 14229
rect 9858 14220 9864 14272
rect 9916 14220 9922 14272
rect 10060 14260 10088 14359
rect 10226 14356 10232 14408
rect 10284 14396 10290 14408
rect 10965 14399 11023 14405
rect 10284 14392 10916 14396
rect 10965 14392 10977 14399
rect 10284 14368 10977 14392
rect 10284 14356 10290 14368
rect 10888 14365 10977 14368
rect 11011 14365 11023 14399
rect 10888 14364 11023 14365
rect 10965 14359 11023 14364
rect 10410 14288 10416 14340
rect 10468 14328 10474 14340
rect 10597 14331 10655 14337
rect 10597 14328 10609 14331
rect 10468 14300 10609 14328
rect 10468 14288 10474 14300
rect 10597 14297 10609 14300
rect 10643 14297 10655 14331
rect 10597 14291 10655 14297
rect 10137 14263 10195 14269
rect 10137 14260 10149 14263
rect 10060 14232 10149 14260
rect 10137 14229 10149 14232
rect 10183 14229 10195 14263
rect 10137 14223 10195 14229
rect 10318 14220 10324 14272
rect 10376 14260 10382 14272
rect 10505 14263 10563 14269
rect 10505 14260 10517 14263
rect 10376 14232 10517 14260
rect 10376 14220 10382 14232
rect 10505 14229 10517 14232
rect 10551 14229 10563 14263
rect 10980 14260 11008 14359
rect 12250 14356 12256 14408
rect 12308 14396 12314 14408
rect 12308 14368 12374 14396
rect 12308 14356 12314 14368
rect 14090 14356 14096 14408
rect 14148 14356 14154 14408
rect 15470 14356 15476 14408
rect 15528 14356 15534 14408
rect 18340 14396 18368 14427
rect 20346 14424 20352 14436
rect 20404 14424 20410 14476
rect 21450 14424 21456 14476
rect 21508 14464 21514 14476
rect 22020 14464 22048 14504
rect 22925 14501 22937 14504
rect 22971 14501 22983 14535
rect 22925 14495 22983 14501
rect 21508 14436 22048 14464
rect 22097 14467 22155 14473
rect 21508 14424 21514 14436
rect 22097 14433 22109 14467
rect 22143 14464 22155 14467
rect 23474 14464 23480 14476
rect 22143 14436 23480 14464
rect 22143 14433 22155 14436
rect 22097 14427 22155 14433
rect 23474 14424 23480 14436
rect 23532 14424 23538 14476
rect 19705 14399 19763 14405
rect 19705 14396 19717 14399
rect 18340 14368 19717 14396
rect 19705 14365 19717 14368
rect 19751 14396 19763 14399
rect 19797 14399 19855 14405
rect 19797 14396 19809 14399
rect 19751 14368 19809 14396
rect 19751 14365 19763 14368
rect 19705 14359 19763 14365
rect 19797 14365 19809 14368
rect 19843 14365 19855 14399
rect 19797 14359 19855 14365
rect 22373 14399 22431 14405
rect 22373 14365 22385 14399
rect 22419 14365 22431 14399
rect 22373 14359 22431 14365
rect 11238 14288 11244 14340
rect 11296 14288 11302 14340
rect 19150 14288 19156 14340
rect 19208 14328 19214 14340
rect 19208 14300 20654 14328
rect 19208 14288 19214 14300
rect 21818 14288 21824 14340
rect 21876 14288 21882 14340
rect 11256 14260 11284 14288
rect 10980 14232 11284 14260
rect 10505 14223 10563 14229
rect 14458 14220 14464 14272
rect 14516 14260 14522 14272
rect 15841 14263 15899 14269
rect 15841 14260 15853 14263
rect 14516 14232 15853 14260
rect 14516 14220 14522 14232
rect 15841 14229 15853 14232
rect 15887 14229 15899 14263
rect 15841 14223 15899 14229
rect 19242 14220 19248 14272
rect 19300 14220 19306 14272
rect 20165 14263 20223 14269
rect 20165 14229 20177 14263
rect 20211 14260 20223 14263
rect 20254 14260 20260 14272
rect 20211 14232 20260 14260
rect 20211 14229 20223 14232
rect 20165 14223 20223 14229
rect 20254 14220 20260 14232
rect 20312 14220 20318 14272
rect 21634 14220 21640 14272
rect 21692 14260 21698 14272
rect 22189 14263 22247 14269
rect 22189 14260 22201 14263
rect 21692 14232 22201 14260
rect 21692 14220 21698 14232
rect 22189 14229 22201 14232
rect 22235 14229 22247 14263
rect 22388 14260 22416 14359
rect 22462 14356 22468 14408
rect 22520 14356 22526 14408
rect 22738 14356 22744 14408
rect 22796 14396 22802 14408
rect 22848 14405 23152 14406
rect 22848 14399 23167 14405
rect 22848 14396 23121 14399
rect 22796 14378 23121 14396
rect 22796 14368 22876 14378
rect 22796 14356 22802 14368
rect 23109 14365 23121 14378
rect 23155 14365 23167 14399
rect 23109 14359 23167 14365
rect 23198 14356 23204 14408
rect 23256 14356 23262 14408
rect 24210 14356 24216 14408
rect 24268 14396 24274 14408
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 24268 14368 24593 14396
rect 24268 14356 24274 14368
rect 24581 14365 24593 14368
rect 24627 14365 24639 14399
rect 24581 14359 24639 14365
rect 24670 14356 24676 14408
rect 24728 14356 24734 14408
rect 25038 14356 25044 14408
rect 25096 14356 25102 14408
rect 22756 14328 22784 14356
rect 22833 14331 22891 14337
rect 22833 14328 22845 14331
rect 22756 14300 22845 14328
rect 22833 14297 22845 14300
rect 22879 14297 22891 14331
rect 22833 14291 22891 14297
rect 23290 14288 23296 14340
rect 23348 14328 23354 14340
rect 23569 14331 23627 14337
rect 23569 14328 23581 14331
rect 23348 14300 23581 14328
rect 23348 14288 23354 14300
rect 23569 14297 23581 14300
rect 23615 14297 23627 14331
rect 23569 14291 23627 14297
rect 23382 14260 23388 14272
rect 22388 14232 23388 14260
rect 22189 14223 22247 14229
rect 23382 14220 23388 14232
rect 23440 14220 23446 14272
rect 24946 14220 24952 14272
rect 25004 14220 25010 14272
rect 25682 14220 25688 14272
rect 25740 14220 25746 14272
rect 1104 14170 26472 14192
rect 1104 14118 7252 14170
rect 7304 14118 7316 14170
rect 7368 14118 7380 14170
rect 7432 14118 7444 14170
rect 7496 14118 7508 14170
rect 7560 14118 13554 14170
rect 13606 14118 13618 14170
rect 13670 14118 13682 14170
rect 13734 14118 13746 14170
rect 13798 14118 13810 14170
rect 13862 14118 19856 14170
rect 19908 14118 19920 14170
rect 19972 14118 19984 14170
rect 20036 14118 20048 14170
rect 20100 14118 20112 14170
rect 20164 14118 26158 14170
rect 26210 14118 26222 14170
rect 26274 14118 26286 14170
rect 26338 14118 26350 14170
rect 26402 14118 26414 14170
rect 26466 14118 26472 14170
rect 1104 14096 26472 14118
rect 8294 14056 8300 14068
rect 6564 14028 8300 14056
rect 3053 13991 3111 13997
rect 3053 13957 3065 13991
rect 3099 13988 3111 13991
rect 3326 13988 3332 14000
rect 3099 13960 3332 13988
rect 3099 13957 3111 13960
rect 3053 13951 3111 13957
rect 3326 13948 3332 13960
rect 3384 13948 3390 14000
rect 5537 13991 5595 13997
rect 5537 13957 5549 13991
rect 5583 13988 5595 13991
rect 5905 13991 5963 13997
rect 5905 13988 5917 13991
rect 5583 13960 5917 13988
rect 5583 13957 5595 13960
rect 5537 13951 5595 13957
rect 5905 13957 5917 13960
rect 5951 13957 5963 13991
rect 5905 13951 5963 13957
rect 5997 13991 6055 13997
rect 5997 13957 6009 13991
rect 6043 13988 6055 13991
rect 6457 13991 6515 13997
rect 6457 13988 6469 13991
rect 6043 13960 6469 13988
rect 6043 13957 6055 13960
rect 5997 13951 6055 13957
rect 6457 13957 6469 13960
rect 6503 13957 6515 13991
rect 6457 13951 6515 13957
rect 2590 13880 2596 13932
rect 2648 13920 2654 13932
rect 2777 13923 2835 13929
rect 2777 13920 2789 13923
rect 2648 13892 2789 13920
rect 2648 13880 2654 13892
rect 2777 13889 2789 13892
rect 2823 13889 2835 13923
rect 4890 13920 4896 13932
rect 4186 13906 4896 13920
rect 2777 13883 2835 13889
rect 4172 13892 4896 13906
rect 3142 13812 3148 13864
rect 3200 13852 3206 13864
rect 4172 13852 4200 13892
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 4985 13923 5043 13929
rect 4985 13889 4997 13923
rect 5031 13920 5043 13923
rect 5074 13920 5080 13932
rect 5031 13892 5080 13920
rect 5031 13889 5043 13892
rect 4985 13883 5043 13889
rect 5074 13880 5080 13892
rect 5132 13880 5138 13932
rect 5813 13923 5871 13929
rect 5813 13889 5825 13923
rect 5859 13920 5871 13923
rect 5859 13892 6040 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 3200 13824 4200 13852
rect 3200 13812 3206 13824
rect 4798 13812 4804 13864
rect 4856 13852 4862 13864
rect 4856 13824 5764 13852
rect 4856 13812 4862 13824
rect 5626 13676 5632 13728
rect 5684 13676 5690 13728
rect 5736 13716 5764 13824
rect 6012 13796 6040 13892
rect 6178 13880 6184 13932
rect 6236 13880 6242 13932
rect 6564 13929 6592 14028
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 8938 14016 8944 14068
rect 8996 14056 9002 14068
rect 8996 14028 9536 14056
rect 8996 14016 9002 14028
rect 7742 13948 7748 14000
rect 7800 13948 7806 14000
rect 9122 13988 9128 14000
rect 8786 13960 9128 13988
rect 9122 13948 9128 13960
rect 9180 13948 9186 14000
rect 9217 13991 9275 13997
rect 9217 13957 9229 13991
rect 9263 13988 9275 13991
rect 9306 13988 9312 14000
rect 9263 13960 9312 13988
rect 9263 13957 9275 13960
rect 9217 13951 9275 13957
rect 9306 13948 9312 13960
rect 9364 13948 9370 14000
rect 6365 13923 6423 13929
rect 6365 13889 6377 13923
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 6543 13923 6601 13929
rect 6543 13889 6555 13923
rect 6589 13889 6601 13923
rect 6543 13883 6601 13889
rect 7193 13923 7251 13929
rect 7193 13889 7205 13923
rect 7239 13889 7251 13923
rect 7193 13883 7251 13889
rect 5994 13744 6000 13796
rect 6052 13784 6058 13796
rect 6380 13784 6408 13883
rect 6914 13812 6920 13864
rect 6972 13812 6978 13864
rect 7006 13812 7012 13864
rect 7064 13812 7070 13864
rect 7208 13784 7236 13883
rect 7760 13861 7788 13948
rect 7377 13855 7435 13861
rect 7377 13821 7389 13855
rect 7423 13852 7435 13855
rect 7745 13855 7803 13861
rect 7423 13824 7604 13852
rect 7423 13821 7435 13824
rect 7377 13815 7435 13821
rect 6052 13756 7236 13784
rect 7576 13784 7604 13824
rect 7745 13821 7757 13855
rect 7791 13821 7803 13855
rect 7745 13815 7803 13821
rect 8202 13812 8208 13864
rect 8260 13852 8266 13864
rect 9508 13861 9536 14028
rect 10594 14016 10600 14068
rect 10652 14056 10658 14068
rect 11517 14059 11575 14065
rect 11517 14056 11529 14059
rect 10652 14028 11529 14056
rect 10652 14016 10658 14028
rect 11517 14025 11529 14028
rect 11563 14025 11575 14059
rect 11517 14019 11575 14025
rect 14093 14059 14151 14065
rect 14093 14025 14105 14059
rect 14139 14056 14151 14059
rect 14182 14056 14188 14068
rect 14139 14028 14188 14056
rect 14139 14025 14151 14028
rect 14093 14019 14151 14025
rect 14182 14016 14188 14028
rect 14240 14016 14246 14068
rect 14458 14016 14464 14068
rect 14516 14016 14522 14068
rect 14553 14059 14611 14065
rect 14553 14025 14565 14059
rect 14599 14056 14611 14059
rect 15838 14056 15844 14068
rect 14599 14028 15844 14056
rect 14599 14025 14611 14028
rect 14553 14019 14611 14025
rect 15838 14016 15844 14028
rect 15896 14016 15902 14068
rect 16669 14059 16727 14065
rect 16669 14056 16681 14059
rect 16408 14028 16681 14056
rect 9858 13948 9864 14000
rect 9916 13948 9922 14000
rect 10134 13948 10140 14000
rect 10192 13988 10198 14000
rect 10192 13960 10350 13988
rect 10192 13948 10198 13960
rect 11146 13948 11152 14000
rect 11204 13988 11210 14000
rect 11885 13991 11943 13997
rect 11885 13988 11897 13991
rect 11204 13960 11897 13988
rect 11204 13948 11210 13960
rect 11885 13957 11897 13960
rect 11931 13957 11943 13991
rect 11885 13951 11943 13957
rect 11977 13991 12035 13997
rect 11977 13957 11989 13991
rect 12023 13988 12035 13991
rect 13906 13988 13912 14000
rect 12023 13960 13912 13988
rect 12023 13957 12035 13960
rect 11977 13951 12035 13957
rect 13906 13948 13912 13960
rect 13964 13948 13970 14000
rect 14200 13960 16344 13988
rect 14200 13920 14228 13960
rect 11992 13892 14228 13920
rect 9493 13855 9551 13861
rect 8260 13824 9444 13852
rect 8260 13812 8266 13824
rect 7576 13756 8248 13784
rect 6052 13744 6058 13756
rect 7374 13716 7380 13728
rect 5736 13688 7380 13716
rect 7374 13676 7380 13688
rect 7432 13716 7438 13728
rect 7926 13716 7932 13728
rect 7432 13688 7932 13716
rect 7432 13676 7438 13688
rect 7926 13676 7932 13688
rect 7984 13676 7990 13728
rect 8220 13716 8248 13756
rect 9122 13716 9128 13728
rect 8220 13688 9128 13716
rect 9122 13676 9128 13688
rect 9180 13676 9186 13728
rect 9416 13716 9444 13824
rect 9493 13821 9505 13855
rect 9539 13852 9551 13855
rect 9585 13855 9643 13861
rect 9585 13852 9597 13855
rect 9539 13824 9597 13852
rect 9539 13821 9551 13824
rect 9493 13815 9551 13821
rect 9585 13821 9597 13824
rect 9631 13852 9643 13855
rect 10226 13852 10232 13864
rect 9631 13824 10232 13852
rect 9631 13821 9643 13824
rect 9585 13815 9643 13821
rect 10226 13812 10232 13824
rect 10284 13812 10290 13864
rect 10318 13812 10324 13864
rect 10376 13852 10382 13864
rect 11333 13855 11391 13861
rect 11333 13852 11345 13855
rect 10376 13824 11345 13852
rect 10376 13812 10382 13824
rect 11333 13821 11345 13824
rect 11379 13821 11391 13855
rect 11992 13852 12020 13892
rect 14274 13880 14280 13932
rect 14332 13920 14338 13932
rect 14921 13923 14979 13929
rect 14921 13920 14933 13923
rect 14332 13892 14933 13920
rect 14332 13880 14338 13892
rect 14921 13889 14933 13892
rect 14967 13889 14979 13923
rect 14921 13883 14979 13889
rect 11333 13815 11391 13821
rect 11440 13824 12020 13852
rect 12161 13855 12219 13861
rect 11440 13716 11468 13824
rect 12161 13821 12173 13855
rect 12207 13852 12219 13855
rect 14645 13855 14703 13861
rect 12207 13824 12388 13852
rect 12207 13821 12219 13824
rect 12161 13815 12219 13821
rect 12360 13796 12388 13824
rect 14645 13821 14657 13855
rect 14691 13821 14703 13855
rect 16316 13852 16344 13960
rect 16408 13929 16436 14028
rect 16669 14025 16681 14028
rect 16715 14025 16727 14059
rect 16669 14019 16727 14025
rect 17129 14059 17187 14065
rect 17129 14025 17141 14059
rect 17175 14056 17187 14059
rect 17310 14056 17316 14068
rect 17175 14028 17316 14056
rect 17175 14025 17187 14028
rect 17129 14019 17187 14025
rect 17310 14016 17316 14028
rect 17368 14016 17374 14068
rect 18524 14028 19656 14056
rect 18049 13991 18107 13997
rect 18049 13957 18061 13991
rect 18095 13988 18107 13991
rect 18322 13988 18328 14000
rect 18095 13960 18328 13988
rect 18095 13957 18107 13960
rect 18049 13951 18107 13957
rect 18322 13948 18328 13960
rect 18380 13948 18386 14000
rect 16393 13923 16451 13929
rect 16393 13889 16405 13923
rect 16439 13889 16451 13923
rect 16393 13883 16451 13889
rect 17034 13880 17040 13932
rect 17092 13880 17098 13932
rect 18524 13920 18552 14028
rect 19150 13948 19156 14000
rect 19208 13948 19214 14000
rect 19628 13988 19656 14028
rect 19702 14016 19708 14068
rect 19760 14056 19766 14068
rect 21177 14059 21235 14065
rect 21177 14056 21189 14059
rect 19760 14028 21189 14056
rect 19760 14016 19766 14028
rect 21177 14025 21189 14028
rect 21223 14025 21235 14059
rect 21177 14019 21235 14025
rect 21818 14016 21824 14068
rect 21876 14056 21882 14068
rect 21919 14059 21977 14065
rect 21919 14056 21931 14059
rect 21876 14028 21931 14056
rect 21876 14016 21882 14028
rect 21919 14025 21931 14028
rect 21965 14025 21977 14059
rect 21919 14019 21977 14025
rect 22189 14059 22247 14065
rect 22189 14025 22201 14059
rect 22235 14025 22247 14059
rect 22189 14019 22247 14025
rect 23937 14059 23995 14065
rect 23937 14025 23949 14059
rect 23983 14056 23995 14059
rect 24578 14056 24584 14068
rect 23983 14028 24584 14056
rect 23983 14025 23995 14028
rect 23937 14019 23995 14025
rect 20806 13988 20812 14000
rect 19628 13960 20812 13988
rect 20806 13948 20812 13960
rect 20864 13948 20870 14000
rect 21450 13988 21456 14000
rect 21284 13960 21456 13988
rect 21284 13929 21312 13960
rect 21450 13948 21456 13960
rect 21508 13948 21514 14000
rect 21545 13991 21603 13997
rect 21545 13957 21557 13991
rect 21591 13988 21603 13991
rect 21726 13988 21732 14000
rect 21591 13960 21732 13988
rect 21591 13957 21603 13960
rect 21545 13951 21603 13957
rect 21726 13948 21732 13960
rect 21784 13988 21790 14000
rect 22005 13991 22063 13997
rect 22005 13988 22017 13991
rect 21784 13960 22017 13988
rect 21784 13948 21790 13960
rect 22005 13957 22017 13960
rect 22051 13957 22063 13991
rect 22005 13951 22063 13957
rect 17236 13892 18552 13920
rect 21085 13923 21143 13929
rect 17236 13852 17264 13892
rect 21085 13889 21097 13923
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 21269 13923 21327 13929
rect 21269 13889 21281 13923
rect 21315 13889 21327 13923
rect 21269 13883 21327 13889
rect 21361 13923 21419 13929
rect 21361 13889 21373 13923
rect 21407 13920 21419 13923
rect 21407 13892 21588 13920
rect 21407 13889 21419 13892
rect 21361 13883 21419 13889
rect 16316 13824 17264 13852
rect 17313 13855 17371 13861
rect 14645 13815 14703 13821
rect 17313 13821 17325 13855
rect 17359 13821 17371 13855
rect 17313 13815 17371 13821
rect 19797 13855 19855 13861
rect 19797 13821 19809 13855
rect 19843 13852 19855 13855
rect 20073 13855 20131 13861
rect 19843 13824 20024 13852
rect 19843 13821 19855 13824
rect 19797 13815 19855 13821
rect 12342 13744 12348 13796
rect 12400 13784 12406 13796
rect 14660 13784 14688 13815
rect 17328 13784 17356 13815
rect 17862 13784 17868 13796
rect 12400 13756 17868 13784
rect 12400 13744 12406 13756
rect 17862 13744 17868 13756
rect 17920 13744 17926 13796
rect 19996 13784 20024 13824
rect 20073 13821 20085 13855
rect 20119 13852 20131 13855
rect 20438 13852 20444 13864
rect 20119 13824 20444 13852
rect 20119 13821 20131 13824
rect 20073 13815 20131 13821
rect 20438 13812 20444 13824
rect 20496 13812 20502 13864
rect 21100 13852 21128 13883
rect 21560 13864 21588 13892
rect 21634 13880 21640 13932
rect 21692 13880 21698 13932
rect 21821 13923 21879 13929
rect 21821 13889 21833 13923
rect 21867 13889 21879 13923
rect 21821 13883 21879 13889
rect 22097 13923 22155 13929
rect 22097 13889 22109 13923
rect 22143 13920 22155 13923
rect 22204 13920 22232 14019
rect 24578 14016 24584 14028
rect 24636 14016 24642 14068
rect 23569 13991 23627 13997
rect 23569 13988 23581 13991
rect 22143 13892 22232 13920
rect 22296 13960 23581 13988
rect 22143 13889 22155 13892
rect 22097 13883 22155 13889
rect 21542 13852 21548 13864
rect 21100 13824 21548 13852
rect 21542 13812 21548 13824
rect 21600 13852 21606 13864
rect 21836 13852 21864 13883
rect 22296 13852 22324 13960
rect 23569 13957 23581 13960
rect 23615 13957 23627 13991
rect 23569 13951 23627 13957
rect 24026 13948 24032 14000
rect 24084 13988 24090 14000
rect 25409 13991 25467 13997
rect 24084 13960 24242 13988
rect 24084 13948 24090 13960
rect 25409 13957 25421 13991
rect 25455 13988 25467 13991
rect 25682 13988 25688 14000
rect 25455 13960 25688 13988
rect 25455 13957 25467 13960
rect 25409 13951 25467 13957
rect 25682 13948 25688 13960
rect 25740 13948 25746 14000
rect 22373 13923 22431 13929
rect 22373 13889 22385 13923
rect 22419 13920 22431 13923
rect 22738 13920 22744 13932
rect 22419 13892 22744 13920
rect 22419 13889 22431 13892
rect 22373 13883 22431 13889
rect 21600 13824 22324 13852
rect 21600 13812 21606 13824
rect 21361 13787 21419 13793
rect 21361 13784 21373 13787
rect 19996 13756 21373 13784
rect 21361 13753 21373 13756
rect 21407 13753 21419 13787
rect 21361 13747 21419 13753
rect 22186 13744 22192 13796
rect 22244 13784 22250 13796
rect 22388 13784 22416 13883
rect 22738 13880 22744 13892
rect 22796 13880 22802 13932
rect 22830 13880 22836 13932
rect 22888 13920 22894 13932
rect 23382 13920 23388 13932
rect 22888 13892 23388 13920
rect 22888 13880 22894 13892
rect 23382 13880 23388 13892
rect 23440 13880 23446 13932
rect 23753 13923 23811 13929
rect 23753 13889 23765 13923
rect 23799 13889 23811 13923
rect 23753 13883 23811 13889
rect 22462 13812 22468 13864
rect 22520 13852 22526 13864
rect 23198 13852 23204 13864
rect 22520 13824 23204 13852
rect 22520 13812 22526 13824
rect 23198 13812 23204 13824
rect 23256 13812 23262 13864
rect 23768 13852 23796 13883
rect 24394 13852 24400 13864
rect 23768 13824 24400 13852
rect 24394 13812 24400 13824
rect 24452 13812 24458 13864
rect 25682 13812 25688 13864
rect 25740 13812 25746 13864
rect 22244 13756 24440 13784
rect 22244 13744 22250 13756
rect 9416 13688 11468 13716
rect 15010 13676 15016 13728
rect 15068 13676 15074 13728
rect 16209 13719 16267 13725
rect 16209 13685 16221 13719
rect 16255 13716 16267 13719
rect 16298 13716 16304 13728
rect 16255 13688 16304 13716
rect 16255 13685 16267 13688
rect 16209 13679 16267 13685
rect 16298 13676 16304 13688
rect 16356 13676 16362 13728
rect 22462 13676 22468 13728
rect 22520 13716 22526 13728
rect 22646 13716 22652 13728
rect 22520 13688 22652 13716
rect 22520 13676 22526 13688
rect 22646 13676 22652 13688
rect 22704 13676 22710 13728
rect 22741 13719 22799 13725
rect 22741 13685 22753 13719
rect 22787 13716 22799 13719
rect 23382 13716 23388 13728
rect 22787 13688 23388 13716
rect 22787 13685 22799 13688
rect 22741 13679 22799 13685
rect 23382 13676 23388 13688
rect 23440 13676 23446 13728
rect 24412 13716 24440 13756
rect 25314 13716 25320 13728
rect 24412 13688 25320 13716
rect 25314 13676 25320 13688
rect 25372 13676 25378 13728
rect 1104 13626 26312 13648
rect 1104 13574 4101 13626
rect 4153 13574 4165 13626
rect 4217 13574 4229 13626
rect 4281 13574 4293 13626
rect 4345 13574 4357 13626
rect 4409 13574 10403 13626
rect 10455 13574 10467 13626
rect 10519 13574 10531 13626
rect 10583 13574 10595 13626
rect 10647 13574 10659 13626
rect 10711 13574 16705 13626
rect 16757 13574 16769 13626
rect 16821 13574 16833 13626
rect 16885 13574 16897 13626
rect 16949 13574 16961 13626
rect 17013 13574 23007 13626
rect 23059 13574 23071 13626
rect 23123 13574 23135 13626
rect 23187 13574 23199 13626
rect 23251 13574 23263 13626
rect 23315 13574 26312 13626
rect 1104 13552 26312 13574
rect 3881 13515 3939 13521
rect 3881 13481 3893 13515
rect 3927 13512 3939 13515
rect 4982 13512 4988 13524
rect 3927 13484 4988 13512
rect 3927 13481 3939 13484
rect 3881 13475 3939 13481
rect 4982 13472 4988 13484
rect 5040 13472 5046 13524
rect 5626 13472 5632 13524
rect 5684 13472 5690 13524
rect 5718 13472 5724 13524
rect 5776 13512 5782 13524
rect 5905 13515 5963 13521
rect 5905 13512 5917 13515
rect 5776 13484 5917 13512
rect 5776 13472 5782 13484
rect 5905 13481 5917 13484
rect 5951 13481 5963 13515
rect 5905 13475 5963 13481
rect 6086 13472 6092 13524
rect 6144 13512 6150 13524
rect 6362 13512 6368 13524
rect 6144 13484 6368 13512
rect 6144 13472 6150 13484
rect 6362 13472 6368 13484
rect 6420 13472 6426 13524
rect 6822 13472 6828 13524
rect 6880 13472 6886 13524
rect 11054 13512 11060 13524
rect 7208 13484 11060 13512
rect 3145 13447 3203 13453
rect 3145 13413 3157 13447
rect 3191 13444 3203 13447
rect 4338 13444 4344 13456
rect 3191 13416 4344 13444
rect 3191 13413 3203 13416
rect 3145 13407 3203 13413
rect 4338 13404 4344 13416
rect 4396 13404 4402 13456
rect 5353 13379 5411 13385
rect 5353 13345 5365 13379
rect 5399 13376 5411 13379
rect 5644 13376 5672 13472
rect 6178 13404 6184 13456
rect 6236 13444 6242 13456
rect 6454 13444 6460 13456
rect 6236 13416 6460 13444
rect 6236 13404 6242 13416
rect 6454 13404 6460 13416
rect 6512 13404 6518 13456
rect 7208 13453 7236 13484
rect 11054 13472 11060 13484
rect 11112 13472 11118 13524
rect 13906 13472 13912 13524
rect 13964 13512 13970 13524
rect 13964 13484 15424 13512
rect 13964 13472 13970 13484
rect 7193 13447 7251 13453
rect 7193 13413 7205 13447
rect 7239 13413 7251 13447
rect 7193 13407 7251 13413
rect 7374 13404 7380 13456
rect 7432 13404 7438 13456
rect 8478 13404 8484 13456
rect 8536 13444 8542 13456
rect 13173 13447 13231 13453
rect 13173 13444 13185 13447
rect 8536 13416 13185 13444
rect 8536 13404 8542 13416
rect 13173 13413 13185 13416
rect 13219 13413 13231 13447
rect 13173 13407 13231 13413
rect 14734 13404 14740 13456
rect 14792 13444 14798 13456
rect 14921 13447 14979 13453
rect 14921 13444 14933 13447
rect 14792 13416 14933 13444
rect 14792 13404 14798 13416
rect 14921 13413 14933 13416
rect 14967 13413 14979 13447
rect 14921 13407 14979 13413
rect 6549 13379 6607 13385
rect 6549 13376 6561 13379
rect 5399 13348 5672 13376
rect 5828 13348 6561 13376
rect 5399 13345 5411 13348
rect 5353 13339 5411 13345
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13277 1455 13311
rect 3142 13308 3148 13320
rect 2806 13280 3148 13308
rect 1397 13271 1455 13277
rect 1412 13240 1440 13271
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 5629 13311 5687 13317
rect 5629 13277 5641 13311
rect 5675 13277 5687 13311
rect 5629 13271 5687 13277
rect 1578 13240 1584 13252
rect 1412 13212 1584 13240
rect 1578 13200 1584 13212
rect 1636 13200 1642 13252
rect 1670 13200 1676 13252
rect 1728 13200 1734 13252
rect 4890 13200 4896 13252
rect 4948 13200 4954 13252
rect 5644 13240 5672 13271
rect 5718 13268 5724 13320
rect 5776 13308 5782 13320
rect 5828 13317 5856 13348
rect 6549 13345 6561 13348
rect 6595 13376 6607 13379
rect 6733 13379 6791 13385
rect 6733 13376 6745 13379
rect 6595 13348 6745 13376
rect 6595 13345 6607 13348
rect 6549 13339 6607 13345
rect 6733 13345 6745 13348
rect 6779 13376 6791 13379
rect 6914 13376 6920 13388
rect 6779 13348 6920 13376
rect 6779 13345 6791 13348
rect 6733 13339 6791 13345
rect 6914 13336 6920 13348
rect 6972 13376 6978 13388
rect 7561 13379 7619 13385
rect 7561 13376 7573 13379
rect 6972 13348 7328 13376
rect 6972 13336 6978 13348
rect 5813 13311 5871 13317
rect 5813 13308 5825 13311
rect 5776 13280 5825 13308
rect 5776 13268 5782 13280
rect 5813 13277 5825 13280
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 5994 13268 6000 13320
rect 6052 13308 6058 13320
rect 6089 13311 6147 13317
rect 6089 13308 6101 13311
rect 6052 13280 6101 13308
rect 6052 13268 6058 13280
rect 6089 13277 6101 13280
rect 6135 13277 6147 13311
rect 6089 13271 6147 13277
rect 5460 13212 5672 13240
rect 6104 13240 6132 13271
rect 6270 13268 6276 13320
rect 6328 13308 6334 13320
rect 6457 13311 6515 13317
rect 6457 13308 6469 13311
rect 6328 13280 6469 13308
rect 6328 13268 6334 13280
rect 6457 13277 6469 13280
rect 6503 13308 6515 13311
rect 6822 13308 6828 13320
rect 6503 13280 6828 13308
rect 6503 13277 6515 13280
rect 6457 13271 6515 13277
rect 6822 13268 6828 13280
rect 6880 13268 6886 13320
rect 7300 13317 7328 13348
rect 7484 13348 7573 13376
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13277 7067 13311
rect 7009 13271 7067 13277
rect 7285 13311 7343 13317
rect 7285 13277 7297 13311
rect 7331 13277 7343 13311
rect 7285 13271 7343 13277
rect 7024 13240 7052 13271
rect 7484 13240 7512 13348
rect 7561 13345 7573 13348
rect 7607 13345 7619 13379
rect 7561 13339 7619 13345
rect 7650 13336 7656 13388
rect 7708 13376 7714 13388
rect 11977 13379 12035 13385
rect 11977 13376 11989 13379
rect 7708 13348 11989 13376
rect 7708 13336 7714 13348
rect 11977 13345 11989 13348
rect 12023 13345 12035 13379
rect 14458 13376 14464 13388
rect 11977 13339 12035 13345
rect 13740 13348 14464 13376
rect 7742 13268 7748 13320
rect 7800 13308 7806 13320
rect 7837 13311 7895 13317
rect 7837 13308 7849 13311
rect 7800 13280 7849 13308
rect 7800 13268 7806 13280
rect 7837 13277 7849 13280
rect 7883 13277 7895 13311
rect 7837 13271 7895 13277
rect 8202 13268 8208 13320
rect 8260 13268 8266 13320
rect 8754 13268 8760 13320
rect 8812 13268 8818 13320
rect 12526 13268 12532 13320
rect 12584 13268 12590 13320
rect 13170 13268 13176 13320
rect 13228 13268 13234 13320
rect 13740 13317 13768 13348
rect 14458 13336 14464 13348
rect 14516 13376 14522 13388
rect 14645 13379 14703 13385
rect 14645 13376 14657 13379
rect 14516 13348 14657 13376
rect 14516 13336 14522 13348
rect 14645 13345 14657 13348
rect 14691 13345 14703 13379
rect 14645 13339 14703 13345
rect 15396 13320 15424 13484
rect 17034 13472 17040 13524
rect 17092 13512 17098 13524
rect 17770 13512 17776 13524
rect 17092 13484 17776 13512
rect 17092 13472 17098 13484
rect 17770 13472 17776 13484
rect 17828 13472 17834 13524
rect 21726 13472 21732 13524
rect 21784 13472 21790 13524
rect 22186 13512 22192 13524
rect 22066 13484 22192 13512
rect 16298 13336 16304 13388
rect 16356 13336 16362 13388
rect 18506 13376 18512 13388
rect 17420 13348 18512 13376
rect 13357 13311 13415 13317
rect 13357 13277 13369 13311
rect 13403 13277 13415 13311
rect 13357 13271 13415 13277
rect 13725 13311 13783 13317
rect 13725 13277 13737 13311
rect 13771 13277 13783 13311
rect 13725 13271 13783 13277
rect 13909 13311 13967 13317
rect 13909 13277 13921 13311
rect 13955 13308 13967 13311
rect 14274 13308 14280 13320
rect 13955 13280 14280 13308
rect 13955 13277 13967 13280
rect 13909 13271 13967 13277
rect 7653 13243 7711 13249
rect 7653 13240 7665 13243
rect 6104 13212 7665 13240
rect 5460 13184 5488 13212
rect 7653 13209 7665 13212
rect 7699 13209 7711 13243
rect 7653 13203 7711 13209
rect 9030 13200 9036 13252
rect 9088 13200 9094 13252
rect 9398 13200 9404 13252
rect 9456 13200 9462 13252
rect 12544 13240 12572 13268
rect 13372 13240 13400 13271
rect 14274 13268 14280 13280
rect 14332 13308 14338 13320
rect 14369 13311 14427 13317
rect 14369 13308 14381 13311
rect 14332 13280 14381 13308
rect 14332 13268 14338 13280
rect 14369 13277 14381 13280
rect 14415 13277 14427 13311
rect 14369 13271 14427 13277
rect 14844 13280 15332 13308
rect 14090 13240 14096 13252
rect 12544 13212 14096 13240
rect 14090 13200 14096 13212
rect 14148 13240 14154 13252
rect 14185 13243 14243 13249
rect 14185 13240 14197 13243
rect 14148 13212 14197 13240
rect 14148 13200 14154 13212
rect 14185 13209 14197 13212
rect 14231 13209 14243 13243
rect 14844 13240 14872 13280
rect 14185 13203 14243 13209
rect 14476 13212 14872 13240
rect 5442 13132 5448 13184
rect 5500 13132 5506 13184
rect 6270 13132 6276 13184
rect 6328 13132 6334 13184
rect 7561 13175 7619 13181
rect 7561 13141 7573 13175
rect 7607 13172 7619 13175
rect 8386 13172 8392 13184
rect 7607 13144 8392 13172
rect 7607 13141 7619 13144
rect 7561 13135 7619 13141
rect 8386 13132 8392 13144
rect 8444 13132 8450 13184
rect 12621 13175 12679 13181
rect 12621 13141 12633 13175
rect 12667 13172 12679 13175
rect 14476 13172 14504 13212
rect 14918 13200 14924 13252
rect 14976 13240 14982 13252
rect 15197 13243 15255 13249
rect 15197 13240 15209 13243
rect 14976 13212 15209 13240
rect 14976 13200 14982 13212
rect 15197 13209 15209 13212
rect 15243 13209 15255 13243
rect 15304 13240 15332 13280
rect 15378 13268 15384 13320
rect 15436 13268 15442 13320
rect 16022 13268 16028 13320
rect 16080 13268 16086 13320
rect 17420 13294 17448 13348
rect 18506 13336 18512 13348
rect 18564 13376 18570 13388
rect 19150 13376 19156 13388
rect 18564 13348 19156 13376
rect 18564 13336 18570 13348
rect 19150 13336 19156 13348
rect 19208 13336 19214 13388
rect 22066 13376 22094 13484
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 22281 13515 22339 13521
rect 22281 13481 22293 13515
rect 22327 13512 22339 13515
rect 22830 13512 22836 13524
rect 22327 13484 22836 13512
rect 22327 13481 22339 13484
rect 22281 13475 22339 13481
rect 22830 13472 22836 13484
rect 22888 13472 22894 13524
rect 24210 13472 24216 13524
rect 24268 13472 24274 13524
rect 24394 13472 24400 13524
rect 24452 13472 24458 13524
rect 24857 13515 24915 13521
rect 24857 13481 24869 13515
rect 24903 13512 24915 13515
rect 24946 13512 24952 13524
rect 24903 13484 24952 13512
rect 24903 13481 24915 13484
rect 24857 13475 24915 13481
rect 24946 13472 24952 13484
rect 25004 13472 25010 13524
rect 25038 13472 25044 13524
rect 25096 13472 25102 13524
rect 25682 13472 25688 13524
rect 25740 13472 25746 13524
rect 25700 13444 25728 13472
rect 24044 13416 25728 13444
rect 21928 13348 22094 13376
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 18598 13308 18604 13320
rect 18012 13280 18604 13308
rect 18012 13268 18018 13280
rect 18598 13268 18604 13280
rect 18656 13268 18662 13320
rect 21928 13317 21956 13348
rect 22462 13336 22468 13388
rect 22520 13376 22526 13388
rect 23474 13376 23480 13388
rect 22520 13348 23480 13376
rect 22520 13336 22526 13348
rect 23474 13336 23480 13348
rect 23532 13376 23538 13388
rect 24044 13376 24072 13416
rect 25866 13404 25872 13456
rect 25924 13404 25930 13456
rect 23532 13348 24072 13376
rect 24136 13348 25084 13376
rect 23532 13336 23538 13348
rect 21913 13311 21971 13317
rect 21913 13277 21925 13311
rect 21959 13277 21971 13311
rect 21913 13271 21971 13277
rect 22094 13268 22100 13320
rect 22152 13268 22158 13320
rect 24026 13308 24032 13320
rect 23874 13280 24032 13308
rect 24026 13268 24032 13280
rect 24084 13268 24090 13320
rect 22373 13243 22431 13249
rect 15304 13212 15976 13240
rect 15197 13203 15255 13209
rect 12667 13144 14504 13172
rect 14553 13175 14611 13181
rect 12667 13141 12679 13144
rect 12621 13135 12679 13141
rect 14553 13141 14565 13175
rect 14599 13172 14611 13175
rect 14734 13172 14740 13184
rect 14599 13144 14740 13172
rect 14599 13141 14611 13144
rect 14553 13135 14611 13141
rect 14734 13132 14740 13144
rect 14792 13132 14798 13184
rect 15102 13132 15108 13184
rect 15160 13132 15166 13184
rect 15562 13132 15568 13184
rect 15620 13132 15626 13184
rect 15948 13172 15976 13212
rect 22373 13209 22385 13243
rect 22419 13209 22431 13243
rect 22373 13203 22431 13209
rect 20714 13172 20720 13184
rect 15948 13144 20720 13172
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 22388 13172 22416 13203
rect 22738 13200 22744 13252
rect 22796 13200 22802 13252
rect 22554 13172 22560 13184
rect 22388 13144 22560 13172
rect 22554 13132 22560 13144
rect 22612 13172 22618 13184
rect 23382 13172 23388 13184
rect 22612 13144 23388 13172
rect 22612 13132 22618 13144
rect 23382 13132 23388 13144
rect 23440 13172 23446 13184
rect 24136 13172 24164 13348
rect 24673 13311 24731 13317
rect 24673 13277 24685 13311
rect 24719 13308 24731 13311
rect 24762 13308 24768 13320
rect 24719 13280 24768 13308
rect 24719 13277 24731 13280
rect 24673 13271 24731 13277
rect 24762 13268 24768 13280
rect 24820 13268 24826 13320
rect 24949 13311 25007 13317
rect 24949 13277 24961 13311
rect 24995 13277 25007 13311
rect 24949 13271 25007 13277
rect 23440 13144 24164 13172
rect 24964 13172 24992 13271
rect 25056 13249 25084 13348
rect 25130 13336 25136 13388
rect 25188 13336 25194 13388
rect 25314 13268 25320 13320
rect 25372 13268 25378 13320
rect 25682 13268 25688 13320
rect 25740 13268 25746 13320
rect 25041 13243 25099 13249
rect 25041 13209 25053 13243
rect 25087 13209 25099 13243
rect 25041 13203 25099 13209
rect 25501 13175 25559 13181
rect 25501 13172 25513 13175
rect 24964 13144 25513 13172
rect 23440 13132 23446 13144
rect 25501 13141 25513 13144
rect 25547 13141 25559 13175
rect 25501 13135 25559 13141
rect 1104 13082 26472 13104
rect 1104 13030 7252 13082
rect 7304 13030 7316 13082
rect 7368 13030 7380 13082
rect 7432 13030 7444 13082
rect 7496 13030 7508 13082
rect 7560 13030 13554 13082
rect 13606 13030 13618 13082
rect 13670 13030 13682 13082
rect 13734 13030 13746 13082
rect 13798 13030 13810 13082
rect 13862 13030 19856 13082
rect 19908 13030 19920 13082
rect 19972 13030 19984 13082
rect 20036 13030 20048 13082
rect 20100 13030 20112 13082
rect 20164 13030 26158 13082
rect 26210 13030 26222 13082
rect 26274 13030 26286 13082
rect 26338 13030 26350 13082
rect 26402 13030 26414 13082
rect 26466 13030 26472 13082
rect 1104 13008 26472 13030
rect 1578 12928 1584 12980
rect 1636 12928 1642 12980
rect 3145 12971 3203 12977
rect 3145 12937 3157 12971
rect 3191 12968 3203 12971
rect 7561 12971 7619 12977
rect 3191 12940 7512 12968
rect 3191 12937 3203 12940
rect 3145 12931 3203 12937
rect 1596 12900 1624 12928
rect 5718 12900 5724 12912
rect 1412 12872 1624 12900
rect 4264 12872 5724 12900
rect 1412 12841 1440 12872
rect 1397 12835 1455 12841
rect 1397 12801 1409 12835
rect 1443 12801 1455 12835
rect 3142 12832 3148 12844
rect 2806 12804 3148 12832
rect 1397 12795 1455 12801
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 4264 12841 4292 12872
rect 5718 12860 5724 12872
rect 5776 12900 5782 12912
rect 7484 12900 7512 12940
rect 7561 12937 7573 12971
rect 7607 12968 7619 12971
rect 9030 12968 9036 12980
rect 7607 12940 9036 12968
rect 7607 12937 7619 12940
rect 7561 12931 7619 12937
rect 9030 12928 9036 12940
rect 9088 12928 9094 12980
rect 9122 12928 9128 12980
rect 9180 12968 9186 12980
rect 9180 12940 10916 12968
rect 9180 12928 9186 12940
rect 7650 12900 7656 12912
rect 5776 12872 7420 12900
rect 7484 12872 7656 12900
rect 5776 12860 5782 12872
rect 4249 12835 4307 12841
rect 4249 12801 4261 12835
rect 4295 12801 4307 12835
rect 4249 12795 4307 12801
rect 4341 12835 4399 12841
rect 4341 12801 4353 12835
rect 4387 12832 4399 12835
rect 4430 12832 4436 12844
rect 4387 12804 4436 12832
rect 4387 12801 4399 12804
rect 4341 12795 4399 12801
rect 4430 12792 4436 12804
rect 4488 12792 4494 12844
rect 4525 12835 4583 12841
rect 4525 12801 4537 12835
rect 4571 12801 4583 12835
rect 4525 12795 4583 12801
rect 4801 12835 4859 12841
rect 4801 12801 4813 12835
rect 4847 12832 4859 12835
rect 5626 12832 5632 12844
rect 4847 12804 5632 12832
rect 4847 12801 4859 12804
rect 4801 12795 4859 12801
rect 1670 12724 1676 12776
rect 1728 12724 1734 12776
rect 4540 12696 4568 12795
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6012 12804 6561 12832
rect 4890 12724 4896 12776
rect 4948 12764 4954 12776
rect 5442 12764 5448 12776
rect 4948 12736 5448 12764
rect 4948 12724 4954 12736
rect 5442 12724 5448 12736
rect 5500 12764 5506 12776
rect 5537 12767 5595 12773
rect 5537 12764 5549 12767
rect 5500 12736 5549 12764
rect 5500 12724 5506 12736
rect 5537 12733 5549 12736
rect 5583 12733 5595 12767
rect 5537 12727 5595 12733
rect 6012 12708 6040 12804
rect 6549 12801 6561 12804
rect 6595 12832 6607 12835
rect 6638 12832 6644 12844
rect 6595 12804 6644 12832
rect 6595 12801 6607 12804
rect 6549 12795 6607 12801
rect 6638 12792 6644 12804
rect 6696 12792 6702 12844
rect 6840 12841 6868 12872
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 6917 12835 6975 12841
rect 6917 12801 6929 12835
rect 6963 12801 6975 12835
rect 6917 12795 6975 12801
rect 7101 12835 7159 12841
rect 7101 12801 7113 12835
rect 7147 12801 7159 12835
rect 7392 12832 7420 12872
rect 7650 12860 7656 12872
rect 7708 12860 7714 12912
rect 8202 12900 8208 12912
rect 7944 12872 8208 12900
rect 7742 12832 7748 12844
rect 7392 12804 7748 12832
rect 7101 12795 7159 12801
rect 6362 12724 6368 12776
rect 6420 12764 6426 12776
rect 6932 12764 6960 12795
rect 6420 12736 6960 12764
rect 6420 12724 6426 12736
rect 5994 12696 6000 12708
rect 4540 12668 6000 12696
rect 5994 12656 6000 12668
rect 6052 12656 6058 12708
rect 6733 12699 6791 12705
rect 6733 12696 6745 12699
rect 6104 12668 6745 12696
rect 4709 12631 4767 12637
rect 4709 12597 4721 12631
rect 4755 12628 4767 12631
rect 5718 12628 5724 12640
rect 4755 12600 5724 12628
rect 4755 12597 4767 12600
rect 4709 12591 4767 12597
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 5810 12588 5816 12640
rect 5868 12628 5874 12640
rect 6104 12628 6132 12668
rect 6733 12665 6745 12668
rect 6779 12665 6791 12699
rect 6733 12659 6791 12665
rect 6822 12656 6828 12708
rect 6880 12696 6886 12708
rect 7116 12696 7144 12795
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 7944 12841 7972 12872
rect 8202 12860 8208 12872
rect 8260 12860 8266 12912
rect 9582 12900 9588 12912
rect 9522 12872 9588 12900
rect 9582 12860 9588 12872
rect 9640 12860 9646 12912
rect 7929 12835 7987 12841
rect 7929 12801 7941 12835
rect 7975 12801 7987 12835
rect 7929 12795 7987 12801
rect 8018 12792 8024 12844
rect 8076 12792 8082 12844
rect 10888 12841 10916 12940
rect 12066 12928 12072 12980
rect 12124 12968 12130 12980
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 12124 12940 12173 12968
rect 12124 12928 12130 12940
rect 12161 12937 12173 12940
rect 12207 12937 12219 12971
rect 12161 12931 12219 12937
rect 12526 12928 12532 12980
rect 12584 12928 12590 12980
rect 13170 12928 13176 12980
rect 13228 12928 13234 12980
rect 13906 12968 13912 12980
rect 13372 12940 13912 12968
rect 11330 12900 11336 12912
rect 11164 12872 11336 12900
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12801 10931 12835
rect 10873 12795 10931 12801
rect 10962 12792 10968 12844
rect 11020 12792 11026 12844
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12764 7895 12767
rect 7883 12736 8156 12764
rect 7883 12733 7895 12736
rect 7837 12727 7895 12733
rect 6880 12668 7144 12696
rect 6880 12656 6886 12668
rect 5868 12600 6132 12628
rect 5868 12588 5874 12600
rect 6362 12588 6368 12640
rect 6420 12588 6426 12640
rect 7006 12588 7012 12640
rect 7064 12588 7070 12640
rect 7116 12628 7144 12668
rect 7745 12631 7803 12637
rect 7745 12628 7757 12631
rect 7116 12600 7757 12628
rect 7745 12597 7757 12600
rect 7791 12597 7803 12631
rect 8128 12628 8156 12736
rect 8294 12724 8300 12776
rect 8352 12724 8358 12776
rect 9490 12724 9496 12776
rect 9548 12764 9554 12776
rect 11164 12773 11192 12872
rect 11330 12860 11336 12872
rect 11388 12900 11394 12912
rect 11388 12872 12756 12900
rect 11388 12860 11394 12872
rect 11241 12835 11299 12841
rect 11241 12801 11253 12835
rect 11287 12801 11299 12835
rect 11241 12795 11299 12801
rect 11149 12767 11207 12773
rect 11149 12764 11161 12767
rect 9548 12736 11161 12764
rect 9548 12724 9554 12736
rect 11149 12733 11161 12736
rect 11195 12733 11207 12767
rect 11256 12764 11284 12795
rect 12066 12792 12072 12844
rect 12124 12792 12130 12844
rect 12434 12764 12440 12776
rect 11256 12736 12440 12764
rect 11149 12727 11207 12733
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 12618 12724 12624 12776
rect 12676 12724 12682 12776
rect 12728 12773 12756 12872
rect 13372 12841 13400 12940
rect 13906 12928 13912 12940
rect 13964 12928 13970 12980
rect 14553 12971 14611 12977
rect 14553 12937 14565 12971
rect 14599 12968 14611 12971
rect 14918 12968 14924 12980
rect 14599 12940 14924 12968
rect 14599 12937 14611 12940
rect 14553 12931 14611 12937
rect 14918 12928 14924 12940
rect 14976 12928 14982 12980
rect 15102 12928 15108 12980
rect 15160 12928 15166 12980
rect 15562 12928 15568 12980
rect 15620 12968 15626 12980
rect 22465 12971 22523 12977
rect 15620 12940 22094 12968
rect 15620 12928 15626 12940
rect 13648 12872 14412 12900
rect 13648 12841 13676 12872
rect 13357 12835 13415 12841
rect 13357 12801 13369 12835
rect 13403 12801 13415 12835
rect 13357 12795 13415 12801
rect 13633 12835 13691 12841
rect 13633 12801 13645 12835
rect 13679 12801 13691 12835
rect 13633 12795 13691 12801
rect 13817 12835 13875 12841
rect 13817 12801 13829 12835
rect 13863 12832 13875 12835
rect 13992 12835 14050 12841
rect 13863 12804 13952 12832
rect 13863 12801 13875 12804
rect 13817 12795 13875 12801
rect 13924 12776 13952 12804
rect 13992 12801 14004 12835
rect 14038 12801 14050 12835
rect 13992 12795 14050 12801
rect 12713 12767 12771 12773
rect 12713 12733 12725 12767
rect 12759 12733 12771 12767
rect 12713 12727 12771 12733
rect 13906 12724 13912 12776
rect 13964 12724 13970 12776
rect 9766 12656 9772 12708
rect 9824 12696 9830 12708
rect 9824 12668 12434 12696
rect 9824 12656 9830 12668
rect 8754 12628 8760 12640
rect 8128 12600 8760 12628
rect 7745 12591 7803 12597
rect 8754 12588 8760 12600
rect 8812 12588 8818 12640
rect 10689 12631 10747 12637
rect 10689 12597 10701 12631
rect 10735 12628 10747 12631
rect 10778 12628 10784 12640
rect 10735 12600 10784 12628
rect 10735 12597 10747 12600
rect 10689 12591 10747 12597
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 11882 12588 11888 12640
rect 11940 12588 11946 12640
rect 12406 12628 12434 12668
rect 13170 12656 13176 12708
rect 13228 12696 13234 12708
rect 14007 12696 14035 12795
rect 14090 12792 14096 12844
rect 14148 12792 14154 12844
rect 14384 12841 14412 12872
rect 14369 12835 14427 12841
rect 14369 12801 14381 12835
rect 14415 12832 14427 12835
rect 14550 12832 14556 12844
rect 14415 12804 14556 12832
rect 14415 12801 14427 12804
rect 14369 12795 14427 12801
rect 14550 12792 14556 12804
rect 14608 12832 14614 12844
rect 14645 12835 14703 12841
rect 14645 12832 14657 12835
rect 14608 12804 14657 12832
rect 14608 12792 14614 12804
rect 14645 12801 14657 12804
rect 14691 12801 14703 12835
rect 14645 12795 14703 12801
rect 14660 12764 14688 12795
rect 14918 12792 14924 12844
rect 14976 12792 14982 12844
rect 15120 12841 15148 12928
rect 15381 12903 15439 12909
rect 15381 12869 15393 12903
rect 15427 12900 15439 12903
rect 15654 12900 15660 12912
rect 15427 12872 15660 12900
rect 15427 12869 15439 12872
rect 15381 12863 15439 12869
rect 15654 12860 15660 12872
rect 15712 12860 15718 12912
rect 15746 12860 15752 12912
rect 15804 12900 15810 12912
rect 18506 12900 18512 12912
rect 15804 12872 16252 12900
rect 18446 12872 18512 12900
rect 15804 12860 15810 12872
rect 15105 12835 15163 12841
rect 15105 12801 15117 12835
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 15470 12792 15476 12844
rect 15528 12832 15534 12844
rect 16224 12841 16252 12872
rect 18506 12860 18512 12872
rect 18564 12860 18570 12912
rect 20254 12860 20260 12912
rect 20312 12860 20318 12912
rect 15565 12835 15623 12841
rect 15565 12832 15577 12835
rect 15528 12804 15577 12832
rect 15528 12792 15534 12804
rect 15565 12801 15577 12804
rect 15611 12801 15623 12835
rect 15565 12795 15623 12801
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12801 15991 12835
rect 15933 12795 15991 12801
rect 16209 12835 16267 12841
rect 16209 12801 16221 12835
rect 16255 12801 16267 12835
rect 16209 12795 16267 12801
rect 15749 12767 15807 12773
rect 15749 12764 15761 12767
rect 14660 12736 15761 12764
rect 15749 12733 15761 12736
rect 15795 12733 15807 12767
rect 15948 12764 15976 12795
rect 16390 12792 16396 12844
rect 16448 12792 16454 12844
rect 19889 12835 19947 12841
rect 19889 12801 19901 12835
rect 19935 12801 19947 12835
rect 19889 12795 19947 12801
rect 19981 12835 20039 12841
rect 19981 12801 19993 12835
rect 20027 12832 20039 12835
rect 20272 12832 20300 12860
rect 20530 12832 20536 12844
rect 20027 12804 20536 12832
rect 20027 12801 20039 12804
rect 19981 12795 20039 12801
rect 16301 12767 16359 12773
rect 16301 12764 16313 12767
rect 15948 12736 16313 12764
rect 15749 12727 15807 12733
rect 16301 12733 16313 12736
rect 16347 12733 16359 12767
rect 16301 12727 16359 12733
rect 16945 12767 17003 12773
rect 16945 12733 16957 12767
rect 16991 12733 17003 12767
rect 16945 12727 17003 12733
rect 14458 12696 14464 12708
rect 13228 12668 14464 12696
rect 13228 12656 13234 12668
rect 14458 12656 14464 12668
rect 14516 12656 14522 12708
rect 15930 12656 15936 12708
rect 15988 12656 15994 12708
rect 13814 12628 13820 12640
rect 12406 12600 13820 12628
rect 13814 12588 13820 12600
rect 13872 12628 13878 12640
rect 14274 12628 14280 12640
rect 13872 12600 14280 12628
rect 13872 12588 13878 12600
rect 14274 12588 14280 12600
rect 14332 12588 14338 12640
rect 16298 12588 16304 12640
rect 16356 12628 16362 12640
rect 16960 12628 16988 12727
rect 17218 12724 17224 12776
rect 17276 12724 17282 12776
rect 18693 12767 18751 12773
rect 18693 12733 18705 12767
rect 18739 12764 18751 12767
rect 19337 12767 19395 12773
rect 19337 12764 19349 12767
rect 18739 12736 19349 12764
rect 18739 12733 18751 12736
rect 18693 12727 18751 12733
rect 19337 12733 19349 12736
rect 19383 12764 19395 12767
rect 19610 12764 19616 12776
rect 19383 12736 19616 12764
rect 19383 12733 19395 12736
rect 19337 12727 19395 12733
rect 19610 12724 19616 12736
rect 19668 12724 19674 12776
rect 19904 12764 19932 12795
rect 20530 12792 20536 12804
rect 20588 12792 20594 12844
rect 22066 12832 22094 12940
rect 22465 12937 22477 12971
rect 22511 12968 22523 12971
rect 22738 12968 22744 12980
rect 22511 12940 22744 12968
rect 22511 12937 22523 12940
rect 22465 12931 22523 12937
rect 22738 12928 22744 12940
rect 22796 12928 22802 12980
rect 24670 12928 24676 12980
rect 24728 12968 24734 12980
rect 25225 12971 25283 12977
rect 25225 12968 25237 12971
rect 24728 12940 25237 12968
rect 24728 12928 24734 12940
rect 25225 12937 25237 12940
rect 25271 12937 25283 12971
rect 25225 12931 25283 12937
rect 23750 12860 23756 12912
rect 23808 12860 23814 12912
rect 24026 12860 24032 12912
rect 24084 12900 24090 12912
rect 24084 12872 24242 12900
rect 24084 12860 24090 12872
rect 22066 12804 23152 12832
rect 20346 12764 20352 12776
rect 19904 12736 20352 12764
rect 20346 12724 20352 12736
rect 20404 12724 20410 12776
rect 23017 12767 23075 12773
rect 23017 12733 23029 12767
rect 23063 12733 23075 12767
rect 23124 12764 23152 12804
rect 23474 12792 23480 12844
rect 23532 12792 23538 12844
rect 25222 12764 25228 12776
rect 23124 12736 25228 12764
rect 23017 12727 23075 12733
rect 18414 12628 18420 12640
rect 16356 12600 18420 12628
rect 16356 12588 16362 12600
rect 18414 12588 18420 12600
rect 18472 12588 18478 12640
rect 18782 12588 18788 12640
rect 18840 12588 18846 12640
rect 20165 12631 20223 12637
rect 20165 12597 20177 12631
rect 20211 12628 20223 12631
rect 20990 12628 20996 12640
rect 20211 12600 20996 12628
rect 20211 12597 20223 12600
rect 20165 12591 20223 12597
rect 20990 12588 20996 12600
rect 21048 12588 21054 12640
rect 22094 12588 22100 12640
rect 22152 12628 22158 12640
rect 23032 12628 23060 12727
rect 25222 12724 25228 12736
rect 25280 12724 25286 12776
rect 23290 12628 23296 12640
rect 22152 12600 23296 12628
rect 22152 12588 22158 12600
rect 23290 12588 23296 12600
rect 23348 12628 23354 12640
rect 25130 12628 25136 12640
rect 23348 12600 25136 12628
rect 23348 12588 23354 12600
rect 25130 12588 25136 12600
rect 25188 12588 25194 12640
rect 1104 12538 26312 12560
rect 1104 12486 4101 12538
rect 4153 12486 4165 12538
rect 4217 12486 4229 12538
rect 4281 12486 4293 12538
rect 4345 12486 4357 12538
rect 4409 12486 10403 12538
rect 10455 12486 10467 12538
rect 10519 12486 10531 12538
rect 10583 12486 10595 12538
rect 10647 12486 10659 12538
rect 10711 12486 16705 12538
rect 16757 12486 16769 12538
rect 16821 12486 16833 12538
rect 16885 12486 16897 12538
rect 16949 12486 16961 12538
rect 17013 12486 23007 12538
rect 23059 12486 23071 12538
rect 23123 12486 23135 12538
rect 23187 12486 23199 12538
rect 23251 12486 23263 12538
rect 23315 12486 26312 12538
rect 1104 12464 26312 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 1670 12424 1676 12436
rect 1627 12396 1676 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 1670 12384 1676 12396
rect 1728 12384 1734 12436
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 8941 12427 8999 12433
rect 8941 12424 8953 12427
rect 8352 12396 8953 12424
rect 8352 12384 8358 12396
rect 8941 12393 8953 12396
rect 8987 12393 8999 12427
rect 8941 12387 8999 12393
rect 9048 12396 11836 12424
rect 5718 12316 5724 12368
rect 5776 12356 5782 12368
rect 6641 12359 6699 12365
rect 6641 12356 6653 12359
rect 5776 12328 6653 12356
rect 5776 12316 5782 12328
rect 6641 12325 6653 12328
rect 6687 12325 6699 12359
rect 6641 12319 6699 12325
rect 7834 12316 7840 12368
rect 7892 12356 7898 12368
rect 9048 12356 9076 12396
rect 7892 12328 9076 12356
rect 11808 12356 11836 12396
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 12621 12427 12679 12433
rect 12621 12424 12633 12427
rect 12492 12396 12633 12424
rect 12492 12384 12498 12396
rect 12621 12393 12633 12396
rect 12667 12393 12679 12427
rect 12621 12387 12679 12393
rect 12710 12384 12716 12436
rect 12768 12424 12774 12436
rect 13357 12427 13415 12433
rect 13357 12424 13369 12427
rect 12768 12396 13369 12424
rect 12768 12384 12774 12396
rect 13357 12393 13369 12396
rect 13403 12393 13415 12427
rect 15565 12427 15623 12433
rect 15565 12424 15577 12427
rect 13357 12387 13415 12393
rect 14844 12396 15577 12424
rect 11808 12328 13584 12356
rect 7892 12316 7898 12328
rect 3694 12248 3700 12300
rect 3752 12288 3758 12300
rect 4341 12291 4399 12297
rect 4341 12288 4353 12291
rect 3752 12260 4353 12288
rect 3752 12248 3758 12260
rect 4341 12257 4353 12260
rect 4387 12257 4399 12291
rect 4341 12251 4399 12257
rect 4706 12248 4712 12300
rect 4764 12248 4770 12300
rect 6086 12248 6092 12300
rect 6144 12288 6150 12300
rect 6144 12260 6316 12288
rect 6144 12248 6150 12260
rect 934 12180 940 12232
rect 992 12220 998 12232
rect 1397 12223 1455 12229
rect 1397 12220 1409 12223
rect 992 12192 1409 12220
rect 992 12180 998 12192
rect 1397 12189 1409 12192
rect 1443 12189 1455 12223
rect 1397 12183 1455 12189
rect 1765 12223 1823 12229
rect 1765 12189 1777 12223
rect 1811 12189 1823 12223
rect 1765 12183 1823 12189
rect 1780 12152 1808 12183
rect 5534 12180 5540 12232
rect 5592 12180 5598 12232
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 6288 12229 6316 12260
rect 6730 12248 6736 12300
rect 6788 12288 6794 12300
rect 9585 12291 9643 12297
rect 6788 12260 7052 12288
rect 6788 12248 6794 12260
rect 6181 12223 6239 12229
rect 6181 12220 6193 12223
rect 5960 12192 6193 12220
rect 5960 12180 5966 12192
rect 6181 12189 6193 12192
rect 6227 12189 6239 12223
rect 6181 12183 6239 12189
rect 6273 12223 6331 12229
rect 6273 12189 6285 12223
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 1412 12124 1808 12152
rect 1412 12096 1440 12124
rect 2038 12112 2044 12164
rect 2096 12112 2102 12164
rect 2774 12112 2780 12164
rect 2832 12112 2838 12164
rect 3970 12152 3976 12164
rect 3528 12124 3976 12152
rect 1394 12044 1400 12096
rect 1452 12044 1458 12096
rect 3528 12093 3556 12124
rect 3970 12112 3976 12124
rect 4028 12152 4034 12164
rect 4157 12155 4215 12161
rect 4157 12152 4169 12155
rect 4028 12124 4169 12152
rect 4028 12112 4034 12124
rect 4157 12121 4169 12124
rect 4203 12121 4215 12155
rect 4157 12115 4215 12121
rect 6362 12112 6368 12164
rect 6420 12112 6426 12164
rect 6564 12152 6592 12183
rect 6638 12180 6644 12232
rect 6696 12220 6702 12232
rect 6825 12223 6883 12229
rect 6825 12220 6837 12223
rect 6696 12192 6837 12220
rect 6696 12180 6702 12192
rect 6825 12189 6837 12192
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 6914 12180 6920 12232
rect 6972 12180 6978 12232
rect 7024 12229 7052 12260
rect 9585 12257 9597 12291
rect 9631 12288 9643 12291
rect 9766 12288 9772 12300
rect 9631 12260 9772 12288
rect 9631 12257 9643 12260
rect 9585 12251 9643 12257
rect 9766 12248 9772 12260
rect 9824 12248 9830 12300
rect 10226 12248 10232 12300
rect 10284 12288 10290 12300
rect 10505 12291 10563 12297
rect 10505 12288 10517 12291
rect 10284 12260 10517 12288
rect 10284 12248 10290 12260
rect 10505 12257 10517 12260
rect 10551 12288 10563 12291
rect 11146 12288 11152 12300
rect 10551 12260 11152 12288
rect 10551 12257 10563 12260
rect 10505 12251 10563 12257
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 12529 12291 12587 12297
rect 12529 12257 12541 12291
rect 12575 12288 12587 12291
rect 13170 12288 13176 12300
rect 12575 12260 13176 12288
rect 12575 12257 12587 12260
rect 12529 12251 12587 12257
rect 13170 12248 13176 12260
rect 13228 12248 13234 12300
rect 7009 12223 7067 12229
rect 7009 12189 7021 12223
rect 7055 12189 7067 12223
rect 7009 12183 7067 12189
rect 7098 12180 7104 12232
rect 7156 12220 7162 12232
rect 7193 12223 7251 12229
rect 7193 12220 7205 12223
rect 7156 12192 7205 12220
rect 7156 12180 7162 12192
rect 7193 12189 7205 12192
rect 7239 12189 7251 12223
rect 7193 12183 7251 12189
rect 8386 12180 8392 12232
rect 8444 12220 8450 12232
rect 9066 12223 9124 12229
rect 9066 12220 9078 12223
rect 8444 12192 9078 12220
rect 8444 12180 8450 12192
rect 9066 12189 9078 12192
rect 9112 12189 9124 12223
rect 9066 12183 9124 12189
rect 9398 12180 9404 12232
rect 9456 12220 9462 12232
rect 9493 12223 9551 12229
rect 9493 12220 9505 12223
rect 9456 12192 9505 12220
rect 9456 12180 9462 12192
rect 9493 12189 9505 12192
rect 9539 12189 9551 12223
rect 9493 12183 9551 12189
rect 10134 12180 10140 12232
rect 10192 12180 10198 12232
rect 13556 12229 13584 12328
rect 14090 12316 14096 12368
rect 14148 12316 14154 12368
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 14108 12288 14136 12316
rect 13872 12260 14035 12288
rect 14108 12260 14320 12288
rect 13872 12248 13878 12260
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12189 13599 12223
rect 13541 12183 13599 12189
rect 13633 12223 13691 12229
rect 13633 12189 13645 12223
rect 13679 12189 13691 12223
rect 13633 12183 13691 12189
rect 6564 12124 6960 12152
rect 6932 12096 6960 12124
rect 3513 12087 3571 12093
rect 3513 12053 3525 12087
rect 3559 12053 3571 12087
rect 3513 12047 3571 12053
rect 3602 12044 3608 12096
rect 3660 12084 3666 12096
rect 3789 12087 3847 12093
rect 3789 12084 3801 12087
rect 3660 12056 3801 12084
rect 3660 12044 3666 12056
rect 3789 12053 3801 12056
rect 3835 12053 3847 12087
rect 3789 12047 3847 12053
rect 4249 12087 4307 12093
rect 4249 12053 4261 12087
rect 4295 12084 4307 12087
rect 5997 12087 6055 12093
rect 5997 12084 6009 12087
rect 4295 12056 6009 12084
rect 4295 12053 4307 12056
rect 4249 12047 4307 12053
rect 5997 12053 6009 12056
rect 6043 12053 6055 12087
rect 5997 12047 6055 12053
rect 6914 12044 6920 12096
rect 6972 12044 6978 12096
rect 9122 12044 9128 12096
rect 9180 12044 9186 12096
rect 10152 12084 10180 12180
rect 10778 12112 10784 12164
rect 10836 12112 10842 12164
rect 11164 12124 11270 12152
rect 11164 12084 11192 12124
rect 12986 12112 12992 12164
rect 13044 12152 13050 12164
rect 13648 12152 13676 12183
rect 13906 12180 13912 12232
rect 13964 12180 13970 12232
rect 14007 12220 14035 12260
rect 14292 12229 14320 12260
rect 14458 12248 14464 12300
rect 14516 12248 14522 12300
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 14007 12192 14105 12220
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 13044 12124 13676 12152
rect 13725 12155 13783 12161
rect 13044 12112 13050 12124
rect 13725 12121 13737 12155
rect 13771 12152 13783 12155
rect 14476 12152 14504 12248
rect 14844 12232 14872 12396
rect 15565 12393 15577 12396
rect 15611 12393 15623 12427
rect 15565 12387 15623 12393
rect 17218 12384 17224 12436
rect 17276 12424 17282 12436
rect 17313 12427 17371 12433
rect 17313 12424 17325 12427
rect 17276 12396 17325 12424
rect 17276 12384 17282 12396
rect 17313 12393 17325 12396
rect 17359 12393 17371 12427
rect 20898 12424 20904 12436
rect 17313 12387 17371 12393
rect 17420 12396 20904 12424
rect 15105 12291 15163 12297
rect 15105 12257 15117 12291
rect 15151 12288 15163 12291
rect 15286 12288 15292 12300
rect 15151 12260 15292 12288
rect 15151 12257 15163 12260
rect 15105 12251 15163 12257
rect 15286 12248 15292 12260
rect 15344 12248 15350 12300
rect 15654 12248 15660 12300
rect 15712 12288 15718 12300
rect 17420 12288 17448 12396
rect 20898 12384 20904 12396
rect 20956 12384 20962 12436
rect 22094 12384 22100 12436
rect 22152 12424 22158 12436
rect 22189 12427 22247 12433
rect 22189 12424 22201 12427
rect 22152 12396 22201 12424
rect 22152 12384 22158 12396
rect 22189 12393 22201 12396
rect 22235 12393 22247 12427
rect 22189 12387 22247 12393
rect 17696 12328 18184 12356
rect 17696 12300 17724 12328
rect 15712 12260 17448 12288
rect 15712 12248 15718 12260
rect 17678 12248 17684 12300
rect 17736 12248 17742 12300
rect 18046 12248 18052 12300
rect 18104 12248 18110 12300
rect 18156 12297 18184 12328
rect 18141 12291 18199 12297
rect 18141 12257 18153 12291
rect 18187 12257 18199 12291
rect 22462 12288 22468 12300
rect 18141 12251 18199 12257
rect 20456 12260 22468 12288
rect 14645 12223 14703 12229
rect 14543 12201 14601 12207
rect 14543 12167 14555 12201
rect 14589 12167 14601 12201
rect 14645 12189 14657 12223
rect 14691 12189 14703 12223
rect 14645 12183 14703 12189
rect 14543 12164 14601 12167
rect 14543 12161 14556 12164
rect 13771 12124 14504 12152
rect 13771 12121 13783 12124
rect 13725 12115 13783 12121
rect 14550 12112 14556 12161
rect 14608 12112 14614 12164
rect 14660 12152 14688 12183
rect 14826 12180 14832 12232
rect 14884 12180 14890 12232
rect 14918 12180 14924 12232
rect 14976 12220 14982 12232
rect 15197 12223 15255 12229
rect 15197 12220 15209 12223
rect 14976 12192 15209 12220
rect 14976 12180 14982 12192
rect 15197 12189 15209 12192
rect 15243 12189 15255 12223
rect 15197 12183 15255 12189
rect 17497 12223 17555 12229
rect 17497 12189 17509 12223
rect 17543 12220 17555 12223
rect 17957 12223 18015 12229
rect 17543 12192 17632 12220
rect 17543 12189 17555 12192
rect 17497 12183 17555 12189
rect 15010 12152 15016 12164
rect 14660 12124 15016 12152
rect 15010 12112 15016 12124
rect 15068 12152 15074 12164
rect 15378 12152 15384 12164
rect 15068 12124 15384 12152
rect 15068 12112 15074 12124
rect 15378 12112 15384 12124
rect 15436 12112 15442 12164
rect 12342 12084 12348 12096
rect 10152 12056 12348 12084
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 14461 12087 14519 12093
rect 14461 12053 14473 12087
rect 14507 12084 14519 12087
rect 14918 12084 14924 12096
rect 14507 12056 14924 12084
rect 14507 12053 14519 12056
rect 14461 12047 14519 12053
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 15562 12044 15568 12096
rect 15620 12044 15626 12096
rect 15746 12044 15752 12096
rect 15804 12044 15810 12096
rect 17604 12093 17632 12192
rect 17957 12189 17969 12223
rect 18003 12220 18015 12223
rect 18782 12220 18788 12232
rect 18003 12192 18788 12220
rect 18003 12189 18015 12192
rect 17957 12183 18015 12189
rect 18782 12180 18788 12192
rect 18840 12180 18846 12232
rect 20162 12180 20168 12232
rect 20220 12180 20226 12232
rect 20254 12180 20260 12232
rect 20312 12220 20318 12232
rect 20456 12229 20484 12260
rect 22462 12248 22468 12260
rect 22520 12248 22526 12300
rect 20441 12223 20499 12229
rect 20441 12220 20453 12223
rect 20312 12192 20453 12220
rect 20312 12180 20318 12192
rect 20441 12189 20453 12192
rect 20487 12189 20499 12223
rect 20441 12183 20499 12189
rect 20180 12152 20208 12180
rect 20346 12152 20352 12164
rect 17972 12124 20116 12152
rect 20180 12124 20352 12152
rect 17972 12096 18000 12124
rect 17589 12087 17647 12093
rect 17589 12053 17601 12087
rect 17635 12053 17647 12087
rect 17589 12047 17647 12053
rect 17954 12044 17960 12096
rect 18012 12044 18018 12096
rect 18966 12044 18972 12096
rect 19024 12084 19030 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 19024 12056 19625 12084
rect 19024 12044 19030 12056
rect 19613 12053 19625 12056
rect 19659 12053 19671 12087
rect 20088 12084 20116 12124
rect 20346 12112 20352 12124
rect 20404 12112 20410 12164
rect 20714 12112 20720 12164
rect 20772 12112 20778 12164
rect 20824 12124 21206 12152
rect 20824 12084 20852 12124
rect 20088 12056 20852 12084
rect 19613 12047 19671 12053
rect 1104 11994 26472 12016
rect 1104 11942 7252 11994
rect 7304 11942 7316 11994
rect 7368 11942 7380 11994
rect 7432 11942 7444 11994
rect 7496 11942 7508 11994
rect 7560 11942 13554 11994
rect 13606 11942 13618 11994
rect 13670 11942 13682 11994
rect 13734 11942 13746 11994
rect 13798 11942 13810 11994
rect 13862 11942 19856 11994
rect 19908 11942 19920 11994
rect 19972 11942 19984 11994
rect 20036 11942 20048 11994
rect 20100 11942 20112 11994
rect 20164 11942 26158 11994
rect 26210 11942 26222 11994
rect 26274 11942 26286 11994
rect 26338 11942 26350 11994
rect 26402 11942 26414 11994
rect 26466 11942 26472 11994
rect 1104 11920 26472 11942
rect 2038 11840 2044 11892
rect 2096 11880 2102 11892
rect 2685 11883 2743 11889
rect 2685 11880 2697 11883
rect 2096 11852 2697 11880
rect 2096 11840 2102 11852
rect 2685 11849 2697 11852
rect 2731 11849 2743 11883
rect 3602 11880 3608 11892
rect 2685 11843 2743 11849
rect 2884 11852 3608 11880
rect 2774 11704 2780 11756
rect 2832 11704 2838 11756
rect 2884 11753 2912 11852
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 5629 11883 5687 11889
rect 5629 11880 5641 11883
rect 4540 11852 5641 11880
rect 4540 11821 4568 11852
rect 5629 11849 5641 11852
rect 5675 11849 5687 11883
rect 5629 11843 5687 11849
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 10318 11880 10324 11892
rect 9824 11852 10324 11880
rect 9824 11840 9830 11852
rect 10318 11840 10324 11852
rect 10376 11840 10382 11892
rect 13998 11880 14004 11892
rect 10796 11852 14004 11880
rect 10796 11824 10824 11852
rect 13998 11840 14004 11852
rect 14056 11840 14062 11892
rect 14182 11840 14188 11892
rect 14240 11880 14246 11892
rect 14369 11883 14427 11889
rect 14369 11880 14381 11883
rect 14240 11852 14381 11880
rect 14240 11840 14246 11852
rect 14369 11849 14381 11852
rect 14415 11849 14427 11883
rect 14369 11843 14427 11849
rect 15010 11840 15016 11892
rect 15068 11880 15074 11892
rect 15068 11852 15328 11880
rect 15068 11840 15074 11852
rect 4525 11815 4583 11821
rect 4525 11781 4537 11815
rect 4571 11781 4583 11815
rect 4890 11812 4896 11824
rect 4525 11775 4583 11781
rect 4816 11784 4896 11812
rect 4816 11753 4844 11784
rect 4890 11772 4896 11784
rect 4948 11772 4954 11824
rect 5534 11772 5540 11824
rect 5592 11812 5598 11824
rect 10413 11815 10471 11821
rect 10413 11812 10425 11815
rect 5592 11784 10425 11812
rect 5592 11772 5598 11784
rect 10413 11781 10425 11784
rect 10459 11812 10471 11815
rect 10778 11812 10784 11824
rect 10459 11784 10784 11812
rect 10459 11781 10471 11784
rect 10413 11775 10471 11781
rect 10778 11772 10784 11784
rect 10836 11772 10842 11824
rect 11146 11772 11152 11824
rect 11204 11812 11210 11824
rect 11204 11784 11652 11812
rect 11204 11772 11210 11784
rect 11624 11756 11652 11784
rect 11882 11772 11888 11824
rect 11940 11772 11946 11824
rect 12342 11772 12348 11824
rect 12400 11772 12406 11824
rect 13170 11772 13176 11824
rect 13228 11812 13234 11824
rect 13725 11815 13783 11821
rect 13725 11812 13737 11815
rect 13228 11784 13737 11812
rect 13228 11772 13234 11784
rect 13725 11781 13737 11784
rect 13771 11781 13783 11815
rect 13725 11775 13783 11781
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11713 2927 11747
rect 4801 11747 4859 11753
rect 2869 11707 2927 11713
rect 2792 11676 2820 11704
rect 3436 11676 3464 11730
rect 4801 11713 4813 11747
rect 4847 11713 4859 11747
rect 4801 11707 4859 11713
rect 5810 11704 5816 11756
rect 5868 11704 5874 11756
rect 5902 11704 5908 11756
rect 5960 11704 5966 11756
rect 6181 11747 6239 11753
rect 6181 11713 6193 11747
rect 6227 11713 6239 11747
rect 6181 11707 6239 11713
rect 6457 11747 6515 11753
rect 6457 11713 6469 11747
rect 6503 11713 6515 11747
rect 6457 11707 6515 11713
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11744 6607 11747
rect 6638 11744 6644 11756
rect 6595 11716 6644 11744
rect 6595 11713 6607 11716
rect 6549 11707 6607 11713
rect 2792 11648 3464 11676
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11645 4951 11679
rect 4893 11639 4951 11645
rect 5537 11679 5595 11685
rect 5537 11645 5549 11679
rect 5583 11676 5595 11679
rect 6196 11676 6224 11707
rect 5583 11648 6224 11676
rect 6472 11676 6500 11707
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11744 6791 11747
rect 7006 11744 7012 11756
rect 6779 11716 7012 11744
rect 6779 11713 6791 11716
rect 6733 11707 6791 11713
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 9858 11704 9864 11756
rect 9916 11704 9922 11756
rect 10045 11747 10103 11753
rect 10045 11713 10057 11747
rect 10091 11713 10103 11747
rect 10045 11707 10103 11713
rect 7190 11676 7196 11688
rect 6472 11648 7196 11676
rect 5583 11645 5595 11648
rect 5537 11639 5595 11645
rect 3053 11543 3111 11549
rect 3053 11509 3065 11543
rect 3099 11540 3111 11543
rect 3878 11540 3884 11552
rect 3099 11512 3884 11540
rect 3099 11509 3111 11512
rect 3053 11503 3111 11509
rect 3878 11500 3884 11512
rect 3936 11540 3942 11552
rect 4908 11540 4936 11639
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 10060 11676 10088 11707
rect 10318 11704 10324 11756
rect 10376 11742 10382 11756
rect 10376 11714 10419 11742
rect 10376 11704 10382 11714
rect 11606 11704 11612 11756
rect 11664 11704 11670 11756
rect 13630 11704 13636 11756
rect 13688 11704 13694 11756
rect 13740 11744 13768 11775
rect 13814 11772 13820 11824
rect 13872 11812 13878 11824
rect 13909 11815 13967 11821
rect 13909 11812 13921 11815
rect 13872 11784 13921 11812
rect 13872 11772 13878 11784
rect 13909 11781 13921 11784
rect 13955 11781 13967 11815
rect 14553 11815 14611 11821
rect 14553 11812 14565 11815
rect 13909 11775 13967 11781
rect 14016 11784 14565 11812
rect 14016 11744 14044 11784
rect 14553 11781 14565 11784
rect 14599 11812 14611 11815
rect 14826 11812 14832 11824
rect 14599 11784 14832 11812
rect 14599 11781 14611 11784
rect 14553 11775 14611 11781
rect 14826 11772 14832 11784
rect 14884 11772 14890 11824
rect 14936 11784 15148 11812
rect 13740 11716 14044 11744
rect 14090 11704 14096 11756
rect 14148 11744 14154 11756
rect 14277 11747 14335 11753
rect 14277 11744 14289 11747
rect 14148 11716 14289 11744
rect 14148 11704 14154 11716
rect 14277 11713 14289 11716
rect 14323 11713 14335 11747
rect 14277 11707 14335 11713
rect 14642 11704 14648 11756
rect 14700 11744 14706 11756
rect 14936 11753 14964 11784
rect 14921 11747 14979 11753
rect 14921 11744 14933 11747
rect 14700 11716 14933 11744
rect 14700 11704 14706 11716
rect 14921 11713 14933 11716
rect 14967 11713 14979 11747
rect 14921 11707 14979 11713
rect 15010 11704 15016 11756
rect 15068 11704 15074 11756
rect 9784 11648 10088 11676
rect 13357 11679 13415 11685
rect 9398 11608 9404 11620
rect 6104 11580 9404 11608
rect 3936 11512 4936 11540
rect 3936 11500 3942 11512
rect 5534 11500 5540 11552
rect 5592 11540 5598 11552
rect 6104 11549 6132 11580
rect 9398 11568 9404 11580
rect 9456 11568 9462 11620
rect 6089 11543 6147 11549
rect 6089 11540 6101 11543
rect 5592 11512 6101 11540
rect 5592 11500 5598 11512
rect 6089 11509 6101 11512
rect 6135 11509 6147 11543
rect 6089 11503 6147 11509
rect 6730 11500 6736 11552
rect 6788 11500 6794 11552
rect 9582 11500 9588 11552
rect 9640 11540 9646 11552
rect 9784 11540 9812 11648
rect 13357 11645 13369 11679
rect 13403 11676 13415 11679
rect 14108 11676 14136 11704
rect 13403 11648 14136 11676
rect 13403 11645 13415 11648
rect 13357 11639 13415 11645
rect 14550 11636 14556 11688
rect 14608 11676 14614 11688
rect 15028 11676 15056 11704
rect 14608 11648 15056 11676
rect 15120 11676 15148 11784
rect 15300 11753 15328 11852
rect 15378 11840 15384 11892
rect 15436 11840 15442 11892
rect 15657 11883 15715 11889
rect 15657 11849 15669 11883
rect 15703 11880 15715 11883
rect 16298 11880 16304 11892
rect 15703 11852 16304 11880
rect 15703 11849 15715 11852
rect 15657 11843 15715 11849
rect 16298 11840 16304 11852
rect 16356 11840 16362 11892
rect 19076 11852 19840 11880
rect 15396 11812 15424 11840
rect 18230 11812 18236 11824
rect 15396 11784 15792 11812
rect 15289 11747 15347 11753
rect 15289 11713 15301 11747
rect 15335 11713 15347 11747
rect 15289 11707 15347 11713
rect 15378 11704 15384 11756
rect 15436 11704 15442 11756
rect 15470 11704 15476 11756
rect 15528 11704 15534 11756
rect 15764 11753 15792 11784
rect 17236 11784 18236 11812
rect 17236 11756 17264 11784
rect 18230 11772 18236 11784
rect 18288 11812 18294 11824
rect 19076 11812 19104 11852
rect 18288 11784 19182 11812
rect 18288 11772 18294 11784
rect 15749 11747 15807 11753
rect 15749 11713 15761 11747
rect 15795 11713 15807 11747
rect 15749 11707 15807 11713
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 15488 11676 15516 11704
rect 15657 11679 15715 11685
rect 15657 11676 15669 11679
rect 15120 11648 15669 11676
rect 14608 11636 14614 11648
rect 15657 11645 15669 11648
rect 15703 11676 15715 11679
rect 15948 11676 15976 11707
rect 17218 11704 17224 11756
rect 17276 11704 17282 11756
rect 18414 11704 18420 11756
rect 18472 11704 18478 11756
rect 19812 11744 19840 11852
rect 24762 11840 24768 11892
rect 24820 11880 24826 11892
rect 24949 11883 25007 11889
rect 24949 11880 24961 11883
rect 24820 11852 24961 11880
rect 24820 11840 24826 11852
rect 24949 11849 24961 11852
rect 24995 11849 25007 11883
rect 24949 11843 25007 11849
rect 25225 11883 25283 11889
rect 25225 11849 25237 11883
rect 25271 11880 25283 11883
rect 25682 11880 25688 11892
rect 25271 11852 25688 11880
rect 25271 11849 25283 11852
rect 25225 11843 25283 11849
rect 25682 11840 25688 11852
rect 25740 11840 25746 11892
rect 22278 11772 22284 11824
rect 22336 11812 22342 11824
rect 22738 11812 22744 11824
rect 22336 11784 22744 11812
rect 22336 11772 22342 11784
rect 22738 11772 22744 11784
rect 22796 11772 22802 11824
rect 24026 11772 24032 11824
rect 24084 11772 24090 11824
rect 20349 11747 20407 11753
rect 20349 11744 20361 11747
rect 19812 11730 20361 11744
rect 19826 11716 20361 11730
rect 20349 11713 20361 11716
rect 20395 11713 20407 11747
rect 20349 11707 20407 11713
rect 20530 11704 20536 11756
rect 20588 11744 20594 11756
rect 21269 11747 21327 11753
rect 21269 11744 21281 11747
rect 20588 11716 21281 11744
rect 20588 11704 20594 11716
rect 21269 11713 21281 11716
rect 21315 11713 21327 11747
rect 21269 11707 21327 11713
rect 21453 11747 21511 11753
rect 21453 11713 21465 11747
rect 21499 11744 21511 11747
rect 21821 11747 21879 11753
rect 21821 11744 21833 11747
rect 21499 11716 21833 11744
rect 21499 11713 21511 11716
rect 21453 11707 21511 11713
rect 21821 11713 21833 11716
rect 21867 11713 21879 11747
rect 21821 11707 21879 11713
rect 22094 11704 22100 11756
rect 22152 11704 22158 11756
rect 22462 11704 22468 11756
rect 22520 11744 22526 11756
rect 23201 11747 23259 11753
rect 23201 11744 23213 11747
rect 22520 11716 23213 11744
rect 22520 11704 22526 11716
rect 23201 11713 23213 11716
rect 23247 11713 23259 11747
rect 23201 11707 23259 11713
rect 25041 11747 25099 11753
rect 25041 11713 25053 11747
rect 25087 11713 25099 11747
rect 25041 11707 25099 11713
rect 15703 11648 15976 11676
rect 15703 11645 15715 11648
rect 15657 11639 15715 11645
rect 16390 11636 16396 11688
rect 16448 11636 16454 11688
rect 18690 11636 18696 11688
rect 18748 11636 18754 11688
rect 20806 11636 20812 11688
rect 20864 11636 20870 11688
rect 21085 11679 21143 11685
rect 21085 11645 21097 11679
rect 21131 11645 21143 11679
rect 21085 11639 21143 11645
rect 9861 11611 9919 11617
rect 9861 11577 9873 11611
rect 9907 11608 9919 11611
rect 11238 11608 11244 11620
rect 9907 11580 11244 11608
rect 9907 11577 9919 11580
rect 9861 11571 9919 11577
rect 11238 11568 11244 11580
rect 11296 11568 11302 11620
rect 13909 11611 13967 11617
rect 13909 11577 13921 11611
rect 13955 11608 13967 11611
rect 15473 11611 15531 11617
rect 15473 11608 15485 11611
rect 13955 11580 15485 11608
rect 13955 11577 13967 11580
rect 13909 11571 13967 11577
rect 15473 11577 15485 11580
rect 15519 11577 15531 11611
rect 16408 11608 16436 11636
rect 21100 11608 21128 11639
rect 23474 11636 23480 11688
rect 23532 11636 23538 11688
rect 15473 11571 15531 11577
rect 15580 11580 16436 11608
rect 20916 11580 21128 11608
rect 10229 11543 10287 11549
rect 10229 11540 10241 11543
rect 9640 11512 10241 11540
rect 9640 11500 9646 11512
rect 10229 11509 10241 11512
rect 10275 11509 10287 11543
rect 10229 11503 10287 11509
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 14553 11543 14611 11549
rect 14553 11540 14565 11543
rect 13872 11512 14565 11540
rect 13872 11500 13878 11512
rect 14553 11509 14565 11512
rect 14599 11540 14611 11543
rect 15580 11540 15608 11580
rect 20916 11552 20944 11580
rect 14599 11512 15608 11540
rect 14599 11509 14611 11512
rect 14553 11503 14611 11509
rect 15838 11500 15844 11552
rect 15896 11500 15902 11552
rect 20165 11543 20223 11549
rect 20165 11509 20177 11543
rect 20211 11540 20223 11543
rect 20346 11540 20352 11552
rect 20211 11512 20352 11540
rect 20211 11509 20223 11512
rect 20165 11503 20223 11509
rect 20346 11500 20352 11512
rect 20404 11500 20410 11552
rect 20898 11500 20904 11552
rect 20956 11500 20962 11552
rect 22002 11500 22008 11552
rect 22060 11500 22066 11552
rect 22281 11543 22339 11549
rect 22281 11509 22293 11543
rect 22327 11540 22339 11543
rect 22554 11540 22560 11552
rect 22327 11512 22560 11540
rect 22327 11509 22339 11512
rect 22281 11503 22339 11509
rect 22554 11500 22560 11512
rect 22612 11500 22618 11552
rect 22830 11500 22836 11552
rect 22888 11540 22894 11552
rect 25056 11540 25084 11707
rect 22888 11512 25084 11540
rect 22888 11500 22894 11512
rect 1104 11450 26312 11472
rect 1104 11398 4101 11450
rect 4153 11398 4165 11450
rect 4217 11398 4229 11450
rect 4281 11398 4293 11450
rect 4345 11398 4357 11450
rect 4409 11398 10403 11450
rect 10455 11398 10467 11450
rect 10519 11398 10531 11450
rect 10583 11398 10595 11450
rect 10647 11398 10659 11450
rect 10711 11398 16705 11450
rect 16757 11398 16769 11450
rect 16821 11398 16833 11450
rect 16885 11398 16897 11450
rect 16949 11398 16961 11450
rect 17013 11398 23007 11450
rect 23059 11398 23071 11450
rect 23123 11398 23135 11450
rect 23187 11398 23199 11450
rect 23251 11398 23263 11450
rect 23315 11398 26312 11450
rect 1104 11376 26312 11398
rect 3694 11296 3700 11348
rect 3752 11336 3758 11348
rect 5534 11336 5540 11348
rect 3752 11308 5540 11336
rect 3752 11296 3758 11308
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 5902 11296 5908 11348
rect 5960 11336 5966 11348
rect 6273 11339 6331 11345
rect 6273 11336 6285 11339
rect 5960 11308 6285 11336
rect 5960 11296 5966 11308
rect 6273 11305 6285 11308
rect 6319 11305 6331 11339
rect 6273 11299 6331 11305
rect 6730 11296 6736 11348
rect 6788 11296 6794 11348
rect 6914 11296 6920 11348
rect 6972 11336 6978 11348
rect 7929 11339 7987 11345
rect 7929 11336 7941 11339
rect 6972 11308 7941 11336
rect 6972 11296 6978 11308
rect 7929 11305 7941 11308
rect 7975 11305 7987 11339
rect 7929 11299 7987 11305
rect 8941 11339 8999 11345
rect 8941 11305 8953 11339
rect 8987 11336 8999 11339
rect 9122 11336 9128 11348
rect 8987 11308 9128 11336
rect 8987 11305 8999 11308
rect 8941 11299 8999 11305
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 10778 11296 10784 11348
rect 10836 11296 10842 11348
rect 10873 11339 10931 11345
rect 10873 11305 10885 11339
rect 10919 11336 10931 11339
rect 18601 11339 18659 11345
rect 10919 11308 11744 11336
rect 10919 11305 10931 11308
rect 10873 11299 10931 11305
rect 3786 11268 3792 11280
rect 2746 11240 3792 11268
rect 1394 11024 1400 11076
rect 1452 11064 1458 11076
rect 2746 11064 2774 11240
rect 3786 11228 3792 11240
rect 3844 11268 3850 11280
rect 4890 11268 4896 11280
rect 3844 11240 4896 11268
rect 3844 11228 3850 11240
rect 4890 11228 4896 11240
rect 4948 11228 4954 11280
rect 6641 11271 6699 11277
rect 6641 11237 6653 11271
rect 6687 11268 6699 11271
rect 6748 11268 6776 11296
rect 6687 11240 6776 11268
rect 6687 11237 6699 11240
rect 6641 11231 6699 11237
rect 7098 11228 7104 11280
rect 7156 11268 7162 11280
rect 7193 11271 7251 11277
rect 7193 11268 7205 11271
rect 7156 11240 7205 11268
rect 7156 11228 7162 11240
rect 7193 11237 7205 11240
rect 7239 11237 7251 11271
rect 7193 11231 7251 11237
rect 7760 11240 10456 11268
rect 4706 11160 4712 11212
rect 4764 11200 4770 11212
rect 5629 11203 5687 11209
rect 5629 11200 5641 11203
rect 4764 11172 5641 11200
rect 4764 11160 4770 11172
rect 5629 11169 5641 11172
rect 5675 11169 5687 11203
rect 5629 11163 5687 11169
rect 6086 11160 6092 11212
rect 6144 11160 6150 11212
rect 6549 11203 6607 11209
rect 6549 11169 6561 11203
rect 6595 11169 6607 11203
rect 6549 11163 6607 11169
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 3142 11132 3148 11144
rect 3099 11104 3148 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 5810 11092 5816 11144
rect 5868 11092 5874 11144
rect 5902 11092 5908 11144
rect 5960 11092 5966 11144
rect 5997 11135 6055 11141
rect 5997 11101 6009 11135
rect 6043 11101 6055 11135
rect 5997 11095 6055 11101
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11101 6515 11135
rect 6564 11132 6592 11163
rect 6638 11132 6644 11144
rect 6564 11104 6644 11132
rect 6457 11095 6515 11101
rect 1452 11036 2774 11064
rect 1452 11024 1458 11036
rect 6012 11008 6040 11095
rect 6472 11064 6500 11095
rect 6638 11092 6644 11104
rect 6696 11092 6702 11144
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11132 6791 11135
rect 7116 11132 7144 11228
rect 7558 11132 7564 11144
rect 6779 11104 7144 11132
rect 7208 11104 7564 11132
rect 6779 11101 6791 11104
rect 6733 11095 6791 11101
rect 7208 11064 7236 11104
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 6472 11036 7236 11064
rect 3602 10956 3608 11008
rect 3660 10956 3666 11008
rect 5994 10956 6000 11008
rect 6052 10996 6058 11008
rect 6362 10996 6368 11008
rect 6052 10968 6368 10996
rect 6052 10956 6058 10968
rect 6362 10956 6368 10968
rect 6420 10996 6426 11008
rect 7101 10999 7159 11005
rect 7101 10996 7113 10999
rect 6420 10968 7113 10996
rect 6420 10956 6426 10968
rect 7101 10965 7113 10968
rect 7147 10996 7159 10999
rect 7760 10996 7788 11240
rect 10428 11212 10456 11240
rect 7926 11160 7932 11212
rect 7984 11200 7990 11212
rect 8113 11203 8171 11209
rect 8113 11200 8125 11203
rect 7984 11172 8125 11200
rect 7984 11160 7990 11172
rect 8113 11169 8125 11172
rect 8159 11169 8171 11203
rect 8570 11200 8576 11212
rect 8113 11163 8171 11169
rect 8220 11172 8576 11200
rect 8220 11141 8248 11172
rect 8570 11160 8576 11172
rect 8628 11200 8634 11212
rect 8938 11200 8944 11212
rect 8628 11172 8944 11200
rect 8628 11160 8634 11172
rect 8938 11160 8944 11172
rect 8996 11200 9002 11212
rect 8996 11172 9260 11200
rect 8996 11160 9002 11172
rect 9232 11141 9260 11172
rect 10410 11160 10416 11212
rect 10468 11160 10474 11212
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11101 8263 11135
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 8205 11095 8263 11101
rect 8864 11104 9137 11132
rect 8864 11008 8892 11104
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11101 9551 11135
rect 9493 11095 9551 11101
rect 9306 11024 9312 11076
rect 9364 11024 9370 11076
rect 7147 10968 7788 10996
rect 7147 10965 7159 10968
rect 7101 10959 7159 10965
rect 8846 10956 8852 11008
rect 8904 10956 8910 11008
rect 9122 10956 9128 11008
rect 9180 10996 9186 11008
rect 9508 10996 9536 11095
rect 9582 11092 9588 11144
rect 9640 11092 9646 11144
rect 10796 11141 10824 11296
rect 11238 11160 11244 11212
rect 11296 11160 11302 11212
rect 11330 11160 11336 11212
rect 11388 11160 11394 11212
rect 11606 11160 11612 11212
rect 11664 11160 11670 11212
rect 11716 11200 11744 11308
rect 18601 11305 18613 11339
rect 18647 11336 18659 11339
rect 18690 11336 18696 11348
rect 18647 11308 18696 11336
rect 18647 11305 18659 11308
rect 18601 11299 18659 11305
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 23474 11296 23480 11348
rect 23532 11336 23538 11348
rect 24397 11339 24455 11345
rect 24397 11336 24409 11339
rect 23532 11308 24409 11336
rect 23532 11296 23538 11308
rect 24397 11305 24409 11308
rect 24443 11305 24455 11339
rect 24397 11299 24455 11305
rect 25314 11296 25320 11348
rect 25372 11296 25378 11348
rect 25133 11271 25191 11277
rect 25133 11237 25145 11271
rect 25179 11237 25191 11271
rect 25133 11231 25191 11237
rect 11885 11203 11943 11209
rect 11885 11200 11897 11203
rect 11716 11172 11897 11200
rect 11885 11169 11897 11172
rect 11931 11169 11943 11203
rect 11885 11163 11943 11169
rect 14642 11160 14648 11212
rect 14700 11200 14706 11212
rect 14737 11203 14795 11209
rect 14737 11200 14749 11203
rect 14700 11172 14749 11200
rect 14700 11160 14706 11172
rect 14737 11169 14749 11172
rect 14783 11169 14795 11203
rect 14737 11163 14795 11169
rect 17402 11160 17408 11212
rect 17460 11200 17466 11212
rect 17957 11203 18015 11209
rect 17957 11200 17969 11203
rect 17460 11172 17969 11200
rect 17460 11160 17466 11172
rect 17957 11169 17969 11172
rect 18003 11169 18015 11203
rect 17957 11163 18015 11169
rect 18414 11160 18420 11212
rect 18472 11200 18478 11212
rect 19245 11203 19303 11209
rect 19245 11200 19257 11203
rect 18472 11172 19257 11200
rect 18472 11160 18478 11172
rect 19245 11169 19257 11172
rect 19291 11169 19303 11203
rect 19245 11163 19303 11169
rect 21082 11160 21088 11212
rect 21140 11160 21146 11212
rect 21542 11160 21548 11212
rect 21600 11200 21606 11212
rect 22002 11200 22008 11212
rect 21600 11172 22008 11200
rect 21600 11160 21606 11172
rect 22002 11160 22008 11172
rect 22060 11200 22066 11212
rect 22186 11200 22192 11212
rect 22060 11172 22192 11200
rect 22060 11160 22066 11172
rect 22186 11160 22192 11172
rect 22244 11160 22250 11212
rect 22462 11160 22468 11212
rect 22520 11200 22526 11212
rect 22833 11203 22891 11209
rect 22833 11200 22845 11203
rect 22520 11172 22845 11200
rect 22520 11160 22526 11172
rect 22833 11169 22845 11172
rect 22879 11200 22891 11203
rect 23661 11203 23719 11209
rect 23661 11200 23673 11203
rect 22879 11172 23673 11200
rect 22879 11169 22891 11172
rect 22833 11163 22891 11169
rect 23661 11169 23673 11172
rect 23707 11169 23719 11203
rect 23661 11163 23719 11169
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11101 10839 11135
rect 10781 11095 10839 11101
rect 11054 11092 11060 11144
rect 11112 11092 11118 11144
rect 11149 11135 11207 11141
rect 11149 11101 11161 11135
rect 11195 11132 11207 11135
rect 11256 11132 11284 11160
rect 11195 11104 11284 11132
rect 11425 11135 11483 11141
rect 11195 11101 11207 11104
rect 11149 11095 11207 11101
rect 11425 11101 11437 11135
rect 11471 11132 11483 11135
rect 14458 11132 14464 11144
rect 11471 11104 11560 11132
rect 11471 11101 11483 11104
rect 11425 11095 11483 11101
rect 10042 11024 10048 11076
rect 10100 11024 10106 11076
rect 9180 10968 9536 10996
rect 9180 10956 9186 10968
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 10778 10996 10784 11008
rect 9732 10968 10784 10996
rect 9732 10956 9738 10968
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 11532 10996 11560 11104
rect 13648 11104 14464 11132
rect 12342 11024 12348 11076
rect 12400 11024 12406 11076
rect 13648 11073 13676 11104
rect 14458 11092 14464 11104
rect 14516 11092 14522 11144
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11132 14611 11135
rect 15746 11132 15752 11144
rect 14599 11104 15752 11132
rect 14599 11101 14611 11104
rect 14553 11095 14611 11101
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 17221 11135 17279 11141
rect 17221 11101 17233 11135
rect 17267 11132 17279 11135
rect 17494 11132 17500 11144
rect 17267 11104 17500 11132
rect 17267 11101 17279 11104
rect 17221 11095 17279 11101
rect 17494 11092 17500 11104
rect 17552 11092 17558 11144
rect 18785 11135 18843 11141
rect 18785 11101 18797 11135
rect 18831 11101 18843 11135
rect 18785 11095 18843 11101
rect 13633 11067 13691 11073
rect 13633 11033 13645 11067
rect 13679 11033 13691 11067
rect 13633 11027 13691 11033
rect 13648 10996 13676 11027
rect 14182 11024 14188 11076
rect 14240 11064 14246 11076
rect 14737 11067 14795 11073
rect 14737 11064 14749 11067
rect 14240 11036 14749 11064
rect 14240 11024 14246 11036
rect 14737 11033 14749 11036
rect 14783 11033 14795 11067
rect 18800 11064 18828 11095
rect 18966 11092 18972 11144
rect 19024 11092 19030 11144
rect 19061 11135 19119 11141
rect 19061 11101 19073 11135
rect 19107 11101 19119 11135
rect 20806 11132 20812 11144
rect 20654 11104 20812 11132
rect 19061 11095 19119 11101
rect 19076 11064 19104 11095
rect 20806 11092 20812 11104
rect 20864 11132 20870 11144
rect 21450 11132 21456 11144
rect 20864 11104 21456 11132
rect 20864 11092 20870 11104
rect 21450 11092 21456 11104
rect 21508 11092 21514 11144
rect 23382 11092 23388 11144
rect 23440 11132 23446 11144
rect 24949 11135 25007 11141
rect 24949 11132 24961 11135
rect 23440 11104 24961 11132
rect 23440 11092 23446 11104
rect 24949 11101 24961 11104
rect 24995 11101 25007 11135
rect 24949 11095 25007 11101
rect 19242 11064 19248 11076
rect 18800 11036 19012 11064
rect 19076 11036 19248 11064
rect 14737 11027 14795 11033
rect 11532 10968 13676 10996
rect 17034 10956 17040 11008
rect 17092 10956 17098 11008
rect 17310 10956 17316 11008
rect 17368 10956 17374 11008
rect 18984 10996 19012 11036
rect 19242 11024 19248 11036
rect 19300 11024 19306 11076
rect 19518 11024 19524 11076
rect 19576 11024 19582 11076
rect 22278 11024 22284 11076
rect 22336 11064 22342 11076
rect 22557 11067 22615 11073
rect 22557 11064 22569 11067
rect 22336 11036 22569 11064
rect 22336 11024 22342 11036
rect 22557 11033 22569 11036
rect 22603 11033 22615 11067
rect 22557 11027 22615 11033
rect 22646 11024 22652 11076
rect 22704 11064 22710 11076
rect 22925 11067 22983 11073
rect 22925 11064 22937 11067
rect 22704 11036 22937 11064
rect 22704 11024 22710 11036
rect 22925 11033 22937 11036
rect 22971 11033 22983 11067
rect 25148 11064 25176 11231
rect 25682 11092 25688 11144
rect 25740 11092 25746 11144
rect 22925 11027 22983 11033
rect 23584 11036 25176 11064
rect 19702 10996 19708 11008
rect 18984 10968 19708 10996
rect 19702 10956 19708 10968
rect 19760 10956 19766 11008
rect 20898 10956 20904 11008
rect 20956 10996 20962 11008
rect 20993 10999 21051 11005
rect 20993 10996 21005 10999
rect 20956 10968 21005 10996
rect 20956 10956 20962 10968
rect 20993 10965 21005 10968
rect 21039 10965 21051 10999
rect 20993 10959 21051 10965
rect 21266 10956 21272 11008
rect 21324 10996 21330 11008
rect 23584 10996 23612 11036
rect 21324 10968 23612 10996
rect 21324 10956 21330 10968
rect 24394 10956 24400 11008
rect 24452 10996 24458 11008
rect 25317 10999 25375 11005
rect 25317 10996 25329 10999
rect 24452 10968 25329 10996
rect 24452 10956 24458 10968
rect 25317 10965 25329 10968
rect 25363 10965 25375 10999
rect 25317 10959 25375 10965
rect 1104 10906 26472 10928
rect 1104 10854 7252 10906
rect 7304 10854 7316 10906
rect 7368 10854 7380 10906
rect 7432 10854 7444 10906
rect 7496 10854 7508 10906
rect 7560 10854 13554 10906
rect 13606 10854 13618 10906
rect 13670 10854 13682 10906
rect 13734 10854 13746 10906
rect 13798 10854 13810 10906
rect 13862 10854 19856 10906
rect 19908 10854 19920 10906
rect 19972 10854 19984 10906
rect 20036 10854 20048 10906
rect 20100 10854 20112 10906
rect 20164 10854 26158 10906
rect 26210 10854 26222 10906
rect 26274 10854 26286 10906
rect 26338 10854 26350 10906
rect 26402 10854 26414 10906
rect 26466 10854 26472 10906
rect 1104 10832 26472 10854
rect 3142 10792 3148 10804
rect 1504 10764 3148 10792
rect 1504 10733 1532 10764
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 5902 10752 5908 10804
rect 5960 10792 5966 10804
rect 6365 10795 6423 10801
rect 6365 10792 6377 10795
rect 5960 10764 6377 10792
rect 5960 10752 5966 10764
rect 6365 10761 6377 10764
rect 6411 10761 6423 10795
rect 6365 10755 6423 10761
rect 6730 10752 6736 10804
rect 6788 10792 6794 10804
rect 7098 10801 7104 10804
rect 7085 10795 7104 10801
rect 6788 10764 7052 10792
rect 6788 10752 6794 10764
rect 1489 10727 1547 10733
rect 1489 10693 1501 10727
rect 1535 10693 1547 10727
rect 1489 10687 1547 10693
rect 2774 10684 2780 10736
rect 2832 10684 2838 10736
rect 3237 10727 3295 10733
rect 3237 10693 3249 10727
rect 3283 10724 3295 10727
rect 4065 10727 4123 10733
rect 4065 10724 4077 10727
rect 3283 10696 4077 10724
rect 3283 10693 3295 10696
rect 3237 10687 3295 10693
rect 4065 10693 4077 10696
rect 4111 10693 4123 10727
rect 5994 10724 6000 10736
rect 4065 10687 4123 10693
rect 5828 10696 6000 10724
rect 3513 10659 3571 10665
rect 3513 10625 3525 10659
rect 3559 10656 3571 10659
rect 3786 10656 3792 10668
rect 3559 10628 3792 10656
rect 3559 10625 3571 10628
rect 3513 10619 3571 10625
rect 3786 10616 3792 10628
rect 3844 10616 3850 10668
rect 3881 10659 3939 10665
rect 3881 10625 3893 10659
rect 3927 10656 3939 10659
rect 4706 10656 4712 10668
rect 3927 10628 4712 10656
rect 3927 10625 3939 10628
rect 3881 10619 3939 10625
rect 4706 10616 4712 10628
rect 4764 10616 4770 10668
rect 5828 10665 5856 10696
rect 5994 10684 6000 10696
rect 6052 10684 6058 10736
rect 6086 10684 6092 10736
rect 6144 10724 6150 10736
rect 7024 10724 7052 10764
rect 7085 10761 7097 10795
rect 7156 10792 7162 10804
rect 7558 10792 7564 10804
rect 7156 10764 7564 10792
rect 7085 10755 7104 10761
rect 7098 10752 7104 10755
rect 7156 10752 7162 10764
rect 7558 10752 7564 10764
rect 7616 10752 7622 10804
rect 8662 10752 8668 10804
rect 8720 10792 8726 10804
rect 8720 10764 8892 10792
rect 8720 10752 8726 10764
rect 7285 10727 7343 10733
rect 7285 10724 7297 10727
rect 6144 10696 6960 10724
rect 7024 10696 7297 10724
rect 6144 10684 6150 10696
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10656 5963 10659
rect 6454 10656 6460 10668
rect 5951 10628 6460 10656
rect 5951 10625 5963 10628
rect 5905 10619 5963 10625
rect 6454 10616 6460 10628
rect 6512 10616 6518 10668
rect 6564 10665 6592 10696
rect 6932 10668 6960 10696
rect 7285 10693 7297 10696
rect 7331 10724 7343 10727
rect 8757 10727 8815 10733
rect 8757 10724 8769 10727
rect 7331 10696 7512 10724
rect 7331 10693 7343 10696
rect 7285 10687 7343 10693
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 3602 10548 3608 10600
rect 3660 10548 3666 10600
rect 5626 10548 5632 10600
rect 5684 10548 5690 10600
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10588 5779 10591
rect 6178 10588 6184 10600
rect 5767 10560 6184 10588
rect 5767 10557 5779 10560
rect 5721 10551 5779 10557
rect 6178 10548 6184 10560
rect 6236 10548 6242 10600
rect 6362 10548 6368 10600
rect 6420 10588 6426 10600
rect 6840 10588 6868 10619
rect 6914 10616 6920 10668
rect 6972 10616 6978 10668
rect 7190 10616 7196 10668
rect 7248 10656 7254 10668
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 7248 10628 7389 10656
rect 7248 10616 7254 10628
rect 7377 10625 7389 10628
rect 7423 10625 7435 10659
rect 7377 10619 7435 10625
rect 7484 10588 7512 10696
rect 8496 10696 8769 10724
rect 8496 10668 8524 10696
rect 8757 10693 8769 10696
rect 8803 10693 8815 10727
rect 8864 10724 8892 10764
rect 8938 10752 8944 10804
rect 8996 10752 9002 10804
rect 9585 10795 9643 10801
rect 9585 10761 9597 10795
rect 9631 10792 9643 10795
rect 9858 10792 9864 10804
rect 9631 10764 9864 10792
rect 9631 10761 9643 10764
rect 9585 10755 9643 10761
rect 9858 10752 9864 10764
rect 9916 10752 9922 10804
rect 9968 10764 10732 10792
rect 9968 10724 9996 10764
rect 8864 10696 9996 10724
rect 8757 10687 8815 10693
rect 10134 10684 10140 10736
rect 10192 10724 10198 10736
rect 10704 10724 10732 10764
rect 10962 10752 10968 10804
rect 11020 10792 11026 10804
rect 11057 10795 11115 10801
rect 11057 10792 11069 10795
rect 11020 10764 11069 10792
rect 11020 10752 11026 10764
rect 11057 10761 11069 10764
rect 11103 10761 11115 10795
rect 11057 10755 11115 10761
rect 16669 10795 16727 10801
rect 16669 10761 16681 10795
rect 16715 10761 16727 10795
rect 16669 10755 16727 10761
rect 17037 10795 17095 10801
rect 17037 10761 17049 10795
rect 17083 10792 17095 10795
rect 17310 10792 17316 10804
rect 17083 10764 17316 10792
rect 17083 10761 17095 10764
rect 17037 10755 17095 10761
rect 10192 10696 10640 10724
rect 10704 10696 16252 10724
rect 10192 10684 10198 10696
rect 7558 10616 7564 10668
rect 7616 10616 7622 10668
rect 8478 10616 8484 10668
rect 8536 10616 8542 10668
rect 8573 10659 8631 10665
rect 8573 10625 8585 10659
rect 8619 10656 8631 10659
rect 8662 10656 8668 10668
rect 8619 10628 8668 10656
rect 8619 10625 8631 10628
rect 8573 10619 8631 10625
rect 8662 10616 8668 10628
rect 8720 10616 8726 10668
rect 8846 10616 8852 10668
rect 8904 10616 8910 10668
rect 9030 10616 9036 10668
rect 9088 10656 9094 10668
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 9088 10628 9137 10656
rect 9088 10616 9094 10628
rect 9125 10625 9137 10628
rect 9171 10656 9183 10659
rect 9306 10656 9312 10668
rect 9171 10628 9312 10656
rect 9171 10625 9183 10628
rect 9125 10619 9183 10625
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 9950 10616 9956 10668
rect 10008 10616 10014 10668
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10656 10103 10659
rect 10226 10656 10232 10668
rect 10091 10628 10232 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 10226 10616 10232 10628
rect 10284 10616 10290 10668
rect 10410 10616 10416 10668
rect 10468 10616 10474 10668
rect 10612 10665 10640 10696
rect 10597 10659 10655 10665
rect 10597 10625 10609 10659
rect 10643 10625 10655 10659
rect 10597 10619 10655 10625
rect 10686 10616 10692 10668
rect 10744 10616 10750 10668
rect 10778 10616 10784 10668
rect 10836 10616 10842 10668
rect 8754 10588 8760 10600
rect 6420 10560 7328 10588
rect 7484 10560 8760 10588
rect 6420 10548 6426 10560
rect 6638 10480 6644 10532
rect 6696 10480 6702 10532
rect 3050 10412 3056 10464
rect 3108 10452 3114 10464
rect 3694 10452 3700 10464
rect 3108 10424 3700 10452
rect 3108 10412 3114 10424
rect 3694 10412 3700 10424
rect 3752 10412 3758 10464
rect 5442 10412 5448 10464
rect 5500 10412 5506 10464
rect 6656 10452 6684 10480
rect 6917 10455 6975 10461
rect 6917 10452 6929 10455
rect 6656 10424 6929 10452
rect 6917 10421 6929 10424
rect 6963 10421 6975 10455
rect 6917 10415 6975 10421
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 7101 10455 7159 10461
rect 7101 10452 7113 10455
rect 7064 10424 7113 10452
rect 7064 10412 7070 10424
rect 7101 10421 7113 10424
rect 7147 10452 7159 10455
rect 7190 10452 7196 10464
rect 7147 10424 7196 10452
rect 7147 10421 7159 10424
rect 7101 10415 7159 10421
rect 7190 10412 7196 10424
rect 7248 10412 7254 10464
rect 7300 10452 7328 10560
rect 8754 10548 8760 10560
rect 8812 10588 8818 10600
rect 10137 10591 10195 10597
rect 10137 10588 10149 10591
rect 8812 10560 10149 10588
rect 8812 10548 8818 10560
rect 10137 10557 10149 10560
rect 10183 10557 10195 10591
rect 10137 10551 10195 10557
rect 9122 10480 9128 10532
rect 9180 10480 9186 10532
rect 7561 10455 7619 10461
rect 7561 10452 7573 10455
rect 7300 10424 7573 10452
rect 7561 10421 7573 10424
rect 7607 10421 7619 10455
rect 7561 10415 7619 10421
rect 7742 10412 7748 10464
rect 7800 10452 7806 10464
rect 8389 10455 8447 10461
rect 8389 10452 8401 10455
rect 7800 10424 8401 10452
rect 7800 10412 7806 10424
rect 8389 10421 8401 10424
rect 8435 10452 8447 10455
rect 9674 10452 9680 10464
rect 8435 10424 9680 10452
rect 8435 10421 8447 10424
rect 8389 10415 8447 10421
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 9950 10412 9956 10464
rect 10008 10452 10014 10464
rect 10778 10452 10784 10464
rect 10008 10424 10784 10452
rect 10008 10412 10014 10424
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 15654 10412 15660 10464
rect 15712 10452 15718 10464
rect 16022 10452 16028 10464
rect 15712 10424 16028 10452
rect 15712 10412 15718 10424
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 16114 10412 16120 10464
rect 16172 10412 16178 10464
rect 16224 10452 16252 10696
rect 16301 10659 16359 10665
rect 16301 10625 16313 10659
rect 16347 10656 16359 10659
rect 16684 10656 16712 10755
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 17494 10752 17500 10804
rect 17552 10752 17558 10804
rect 18874 10792 18880 10804
rect 17880 10764 18880 10792
rect 17129 10727 17187 10733
rect 17129 10693 17141 10727
rect 17175 10724 17187 10727
rect 17880 10724 17908 10764
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 19242 10752 19248 10804
rect 19300 10752 19306 10804
rect 19337 10795 19395 10801
rect 19337 10761 19349 10795
rect 19383 10792 19395 10795
rect 19518 10792 19524 10804
rect 19383 10764 19524 10792
rect 19383 10761 19395 10764
rect 19337 10755 19395 10761
rect 19518 10752 19524 10764
rect 19576 10752 19582 10804
rect 20165 10795 20223 10801
rect 20165 10761 20177 10795
rect 20211 10792 20223 10795
rect 20622 10792 20628 10804
rect 20211 10764 20628 10792
rect 20211 10761 20223 10764
rect 20165 10755 20223 10761
rect 20622 10752 20628 10764
rect 20680 10752 20686 10804
rect 22462 10752 22468 10804
rect 22520 10752 22526 10804
rect 17175 10696 17908 10724
rect 17957 10727 18015 10733
rect 17175 10693 17187 10696
rect 17129 10687 17187 10693
rect 17957 10693 17969 10727
rect 18003 10724 18015 10727
rect 19150 10724 19156 10736
rect 18003 10696 19156 10724
rect 18003 10693 18015 10696
rect 17957 10687 18015 10693
rect 19150 10684 19156 10696
rect 19208 10684 19214 10736
rect 19260 10724 19288 10752
rect 19705 10727 19763 10733
rect 19260 10696 19656 10724
rect 16347 10628 16712 10656
rect 16347 10625 16359 10628
rect 16301 10619 16359 10625
rect 17770 10616 17776 10668
rect 17828 10656 17834 10668
rect 17865 10659 17923 10665
rect 17865 10656 17877 10659
rect 17828 10628 17877 10656
rect 17828 10616 17834 10628
rect 17865 10625 17877 10628
rect 17911 10625 17923 10659
rect 17865 10619 17923 10625
rect 19061 10659 19119 10665
rect 19061 10625 19073 10659
rect 19107 10625 19119 10659
rect 19061 10619 19119 10625
rect 19245 10659 19303 10665
rect 19245 10625 19257 10659
rect 19291 10656 19303 10659
rect 19426 10656 19432 10668
rect 19291 10628 19432 10656
rect 19291 10625 19303 10628
rect 19245 10619 19303 10625
rect 17313 10591 17371 10597
rect 17313 10557 17325 10591
rect 17359 10557 17371 10591
rect 17313 10551 17371 10557
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 17328 10520 17356 10551
rect 17678 10520 17684 10532
rect 17328 10492 17684 10520
rect 17678 10480 17684 10492
rect 17736 10520 17742 10532
rect 18064 10520 18092 10551
rect 17736 10492 18092 10520
rect 19076 10520 19104 10619
rect 19426 10616 19432 10628
rect 19484 10616 19490 10668
rect 19518 10616 19524 10668
rect 19576 10616 19582 10668
rect 19628 10656 19656 10696
rect 19705 10693 19717 10727
rect 19751 10724 19763 10727
rect 20809 10727 20867 10733
rect 20809 10724 20821 10727
rect 19751 10696 20821 10724
rect 19751 10693 19763 10696
rect 19705 10687 19763 10693
rect 20809 10693 20821 10696
rect 20855 10693 20867 10727
rect 20809 10687 20867 10693
rect 20990 10684 20996 10736
rect 21048 10724 21054 10736
rect 22480 10724 22508 10752
rect 23842 10724 23848 10736
rect 21048 10696 22048 10724
rect 21048 10684 21054 10696
rect 19797 10659 19855 10665
rect 19797 10656 19809 10659
rect 19628 10628 19809 10656
rect 19797 10625 19809 10628
rect 19843 10625 19855 10659
rect 19797 10619 19855 10625
rect 20346 10616 20352 10668
rect 20404 10616 20410 10668
rect 20717 10659 20775 10665
rect 20717 10625 20729 10659
rect 20763 10656 20775 10659
rect 21542 10656 21548 10668
rect 20763 10628 21548 10656
rect 20763 10625 20775 10628
rect 20717 10619 20775 10625
rect 21542 10616 21548 10628
rect 21600 10616 21606 10668
rect 22020 10665 22048 10696
rect 22204 10696 22508 10724
rect 23690 10696 23848 10724
rect 22204 10665 22232 10696
rect 23842 10684 23848 10696
rect 23900 10724 23906 10736
rect 24118 10724 24124 10736
rect 23900 10696 24124 10724
rect 23900 10684 23906 10696
rect 24118 10684 24124 10696
rect 24176 10684 24182 10736
rect 22005 10659 22063 10665
rect 22005 10625 22017 10659
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 22189 10659 22247 10665
rect 22189 10625 22201 10659
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 19153 10591 19211 10597
rect 19153 10557 19165 10591
rect 19199 10588 19211 10591
rect 19889 10591 19947 10597
rect 19889 10588 19901 10591
rect 19199 10560 19901 10588
rect 19199 10557 19211 10560
rect 19153 10551 19211 10557
rect 19889 10557 19901 10560
rect 19935 10557 19947 10591
rect 19889 10551 19947 10557
rect 20073 10591 20131 10597
rect 20073 10557 20085 10591
rect 20119 10588 20131 10591
rect 20806 10588 20812 10600
rect 20119 10560 20812 10588
rect 20119 10557 20131 10560
rect 20073 10551 20131 10557
rect 20806 10548 20812 10560
rect 20864 10548 20870 10600
rect 21361 10591 21419 10597
rect 21361 10588 21373 10591
rect 20916 10560 21373 10588
rect 20916 10532 20944 10560
rect 21361 10557 21373 10560
rect 21407 10557 21419 10591
rect 21361 10551 21419 10557
rect 22465 10591 22523 10597
rect 22465 10557 22477 10591
rect 22511 10588 22523 10591
rect 22554 10588 22560 10600
rect 22511 10560 22560 10588
rect 22511 10557 22523 10560
rect 22465 10551 22523 10557
rect 22554 10548 22560 10560
rect 22612 10548 22618 10600
rect 24210 10588 24216 10600
rect 23952 10560 24216 10588
rect 20898 10520 20904 10532
rect 19076 10492 20904 10520
rect 17736 10480 17742 10492
rect 20898 10480 20904 10492
rect 20956 10480 20962 10532
rect 21008 10492 22094 10520
rect 21008 10452 21036 10492
rect 16224 10424 21036 10452
rect 21818 10412 21824 10464
rect 21876 10412 21882 10464
rect 22066 10452 22094 10492
rect 23952 10452 23980 10560
rect 24210 10548 24216 10560
rect 24268 10548 24274 10600
rect 24394 10548 24400 10600
rect 24452 10588 24458 10600
rect 24489 10591 24547 10597
rect 24489 10588 24501 10591
rect 24452 10560 24501 10588
rect 24452 10548 24458 10560
rect 24489 10557 24501 10560
rect 24535 10557 24547 10591
rect 24489 10551 24547 10557
rect 24946 10548 24952 10600
rect 25004 10588 25010 10600
rect 25225 10591 25283 10597
rect 25225 10588 25237 10591
rect 25004 10560 25237 10588
rect 25004 10548 25010 10560
rect 25225 10557 25237 10560
rect 25271 10557 25283 10591
rect 25225 10551 25283 10557
rect 25774 10548 25780 10600
rect 25832 10548 25838 10600
rect 22066 10424 23980 10452
rect 25133 10455 25191 10461
rect 25133 10421 25145 10455
rect 25179 10452 25191 10455
rect 25498 10452 25504 10464
rect 25179 10424 25504 10452
rect 25179 10421 25191 10424
rect 25133 10415 25191 10421
rect 25498 10412 25504 10424
rect 25556 10412 25562 10464
rect 1104 10362 26312 10384
rect 1104 10310 4101 10362
rect 4153 10310 4165 10362
rect 4217 10310 4229 10362
rect 4281 10310 4293 10362
rect 4345 10310 4357 10362
rect 4409 10310 10403 10362
rect 10455 10310 10467 10362
rect 10519 10310 10531 10362
rect 10583 10310 10595 10362
rect 10647 10310 10659 10362
rect 10711 10310 16705 10362
rect 16757 10310 16769 10362
rect 16821 10310 16833 10362
rect 16885 10310 16897 10362
rect 16949 10310 16961 10362
rect 17013 10310 23007 10362
rect 23059 10310 23071 10362
rect 23123 10310 23135 10362
rect 23187 10310 23199 10362
rect 23251 10310 23263 10362
rect 23315 10310 26312 10362
rect 1104 10288 26312 10310
rect 5442 10248 5448 10260
rect 2608 10220 5448 10248
rect 2608 10053 2636 10220
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 5626 10208 5632 10260
rect 5684 10248 5690 10260
rect 5905 10251 5963 10257
rect 5905 10248 5917 10251
rect 5684 10220 5917 10248
rect 5684 10208 5690 10220
rect 5905 10217 5917 10220
rect 5951 10217 5963 10251
rect 5905 10211 5963 10217
rect 6086 10208 6092 10260
rect 6144 10208 6150 10260
rect 6178 10208 6184 10260
rect 6236 10248 6242 10260
rect 6641 10251 6699 10257
rect 6641 10248 6653 10251
rect 6236 10220 6653 10248
rect 6236 10208 6242 10220
rect 6641 10217 6653 10220
rect 6687 10217 6699 10251
rect 6641 10211 6699 10217
rect 7558 10208 7564 10260
rect 7616 10248 7622 10260
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 7616 10220 7941 10248
rect 7616 10208 7622 10220
rect 7929 10217 7941 10220
rect 7975 10217 7987 10251
rect 7929 10211 7987 10217
rect 8389 10251 8447 10257
rect 8389 10217 8401 10251
rect 8435 10248 8447 10251
rect 8478 10248 8484 10260
rect 8435 10220 8484 10248
rect 8435 10217 8447 10220
rect 8389 10211 8447 10217
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 9030 10208 9036 10260
rect 9088 10208 9094 10260
rect 9858 10208 9864 10260
rect 9916 10208 9922 10260
rect 10226 10208 10232 10260
rect 10284 10248 10290 10260
rect 10597 10251 10655 10257
rect 10597 10248 10609 10251
rect 10284 10220 10609 10248
rect 10284 10208 10290 10220
rect 10597 10217 10609 10220
rect 10643 10217 10655 10251
rect 10597 10211 10655 10217
rect 15920 10251 15978 10257
rect 15920 10217 15932 10251
rect 15966 10248 15978 10251
rect 16114 10248 16120 10260
rect 15966 10220 16120 10248
rect 15966 10217 15978 10220
rect 15920 10211 15978 10217
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 19426 10208 19432 10260
rect 19484 10248 19490 10260
rect 20152 10251 20210 10257
rect 20152 10248 20164 10251
rect 19484 10220 20164 10248
rect 19484 10208 19490 10220
rect 20152 10217 20164 10220
rect 20198 10248 20210 10251
rect 21818 10248 21824 10260
rect 20198 10220 21824 10248
rect 20198 10217 20210 10220
rect 20152 10211 20210 10217
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 22094 10208 22100 10260
rect 22152 10248 22158 10260
rect 22189 10251 22247 10257
rect 22189 10248 22201 10251
rect 22152 10220 22201 10248
rect 22152 10208 22158 10220
rect 22189 10217 22201 10220
rect 22235 10217 22247 10251
rect 22189 10211 22247 10217
rect 22465 10251 22523 10257
rect 22465 10217 22477 10251
rect 22511 10248 22523 10251
rect 23382 10248 23388 10260
rect 22511 10220 23388 10248
rect 22511 10217 22523 10220
rect 22465 10211 22523 10217
rect 23382 10208 23388 10220
rect 23440 10208 23446 10260
rect 24210 10208 24216 10260
rect 24268 10208 24274 10260
rect 25409 10251 25467 10257
rect 25409 10217 25421 10251
rect 25455 10248 25467 10251
rect 25774 10248 25780 10260
rect 25455 10220 25780 10248
rect 25455 10217 25467 10220
rect 25409 10211 25467 10217
rect 25774 10208 25780 10220
rect 25832 10208 25838 10260
rect 4908 10152 12434 10180
rect 2866 10072 2872 10124
rect 2924 10112 2930 10124
rect 4908 10121 4936 10152
rect 4893 10115 4951 10121
rect 2924 10084 4292 10112
rect 2924 10072 2930 10084
rect 2593 10047 2651 10053
rect 2593 10013 2605 10047
rect 2639 10013 2651 10047
rect 2593 10007 2651 10013
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10044 2835 10047
rect 3050 10044 3056 10056
rect 2823 10016 3056 10044
rect 2823 10013 2835 10016
rect 2777 10007 2835 10013
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 3234 9936 3240 9988
rect 3292 9976 3298 9988
rect 3804 9976 3832 10007
rect 3970 10004 3976 10056
rect 4028 10004 4034 10056
rect 4062 10004 4068 10056
rect 4120 10004 4126 10056
rect 4264 10053 4292 10084
rect 4893 10081 4905 10115
rect 4939 10081 4951 10115
rect 4893 10075 4951 10081
rect 5534 10072 5540 10124
rect 5592 10072 5598 10124
rect 5721 10115 5779 10121
rect 5721 10081 5733 10115
rect 5767 10112 5779 10115
rect 6730 10112 6736 10124
rect 5767 10084 6736 10112
rect 5767 10081 5779 10084
rect 5721 10075 5779 10081
rect 6730 10072 6736 10084
rect 6788 10072 6794 10124
rect 7484 10084 7788 10112
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10044 5503 10047
rect 5491 10016 5580 10044
rect 5491 10013 5503 10016
rect 5445 10007 5503 10013
rect 4080 9976 4108 10004
rect 3292 9948 4108 9976
rect 4433 9979 4491 9985
rect 3292 9936 3298 9948
rect 4433 9945 4445 9979
rect 4479 9976 4491 9979
rect 4525 9979 4583 9985
rect 4525 9976 4537 9979
rect 4479 9948 4537 9976
rect 4479 9945 4491 9948
rect 4433 9939 4491 9945
rect 4525 9945 4537 9948
rect 4571 9945 4583 9979
rect 4525 9939 4583 9945
rect 4614 9936 4620 9988
rect 4672 9976 4678 9988
rect 4709 9979 4767 9985
rect 4709 9976 4721 9979
rect 4672 9948 4721 9976
rect 4672 9936 4678 9948
rect 4709 9945 4721 9948
rect 4755 9945 4767 9979
rect 4709 9939 4767 9945
rect 5552 9976 5580 10016
rect 5626 10004 5632 10056
rect 5684 10004 5690 10056
rect 6362 10004 6368 10056
rect 6420 10004 6426 10056
rect 6457 10047 6515 10053
rect 6457 10013 6469 10047
rect 6503 10044 6515 10047
rect 6822 10044 6828 10056
rect 6503 10016 6828 10044
rect 6503 10013 6515 10016
rect 6457 10007 6515 10013
rect 6822 10004 6828 10016
rect 6880 10044 6886 10056
rect 7484 10044 7512 10084
rect 7760 10056 7788 10084
rect 8956 10084 9628 10112
rect 6880 10016 7512 10044
rect 6880 10004 6886 10016
rect 7558 10004 7564 10056
rect 7616 10004 7622 10056
rect 7742 10004 7748 10056
rect 7800 10004 7806 10056
rect 7926 10004 7932 10056
rect 7984 10004 7990 10056
rect 8113 10047 8171 10053
rect 8113 10013 8125 10047
rect 8159 10013 8171 10047
rect 8113 10007 8171 10013
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10044 8447 10047
rect 8662 10044 8668 10056
rect 8435 10016 8668 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 5997 9979 6055 9985
rect 5997 9976 6009 9979
rect 5552 9948 6009 9976
rect 5552 9920 5580 9948
rect 5997 9945 6009 9948
rect 6043 9945 6055 9979
rect 5997 9939 6055 9945
rect 6917 9979 6975 9985
rect 6917 9945 6929 9979
rect 6963 9976 6975 9979
rect 7006 9976 7012 9988
rect 6963 9948 7012 9976
rect 6963 9945 6975 9948
rect 6917 9939 6975 9945
rect 7006 9936 7012 9948
rect 7064 9936 7070 9988
rect 7101 9979 7159 9985
rect 7101 9945 7113 9979
rect 7147 9976 7159 9979
rect 7576 9976 7604 10004
rect 7147 9948 7604 9976
rect 8128 9976 8156 10007
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 8956 10053 8984 10084
rect 8757 10047 8815 10053
rect 8757 10013 8769 10047
rect 8803 10013 8815 10047
rect 8757 10007 8815 10013
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 8772 9976 8800 10007
rect 9140 9976 9168 10007
rect 9398 10004 9404 10056
rect 9456 10004 9462 10056
rect 9493 10047 9551 10053
rect 9493 10013 9505 10047
rect 9539 10013 9551 10047
rect 9600 10044 9628 10084
rect 9674 10072 9680 10124
rect 9732 10112 9738 10124
rect 9732 10084 10548 10112
rect 9732 10072 9738 10084
rect 9769 10047 9827 10053
rect 9600 10016 9674 10044
rect 9493 10007 9551 10013
rect 9508 9976 9536 10007
rect 8128 9948 8984 9976
rect 9140 9948 9536 9976
rect 9646 9976 9674 10016
rect 9769 10013 9781 10047
rect 9815 10044 9827 10047
rect 9950 10044 9956 10056
rect 9815 10016 9956 10044
rect 9815 10013 9827 10016
rect 9769 10007 9827 10013
rect 9950 10004 9956 10016
rect 10008 10044 10014 10056
rect 10045 10047 10103 10053
rect 10045 10044 10057 10047
rect 10008 10016 10057 10044
rect 10008 10004 10014 10016
rect 10045 10013 10057 10016
rect 10091 10013 10103 10047
rect 10045 10007 10103 10013
rect 10137 10047 10195 10053
rect 10137 10013 10149 10047
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 9858 9976 9864 9988
rect 9646 9948 9864 9976
rect 7147 9945 7159 9948
rect 7101 9939 7159 9945
rect 2406 9868 2412 9920
rect 2464 9868 2470 9920
rect 5534 9868 5540 9920
rect 5592 9868 5598 9920
rect 8570 9868 8576 9920
rect 8628 9868 8634 9920
rect 8956 9908 8984 9948
rect 9217 9911 9275 9917
rect 9217 9908 9229 9911
rect 8956 9880 9229 9908
rect 9217 9877 9229 9880
rect 9263 9877 9275 9911
rect 9508 9908 9536 9948
rect 9858 9936 9864 9948
rect 9916 9976 9922 9988
rect 10152 9976 10180 10007
rect 10318 10004 10324 10056
rect 10376 10004 10382 10056
rect 10410 10004 10416 10056
rect 10468 10004 10474 10056
rect 10520 10053 10548 10084
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10013 10563 10047
rect 10505 10007 10563 10013
rect 10686 10004 10692 10056
rect 10744 10004 10750 10056
rect 10781 10047 10839 10053
rect 10781 10013 10793 10047
rect 10827 10013 10839 10047
rect 10781 10007 10839 10013
rect 10594 9976 10600 9988
rect 9916 9948 10600 9976
rect 9916 9936 9922 9948
rect 10594 9936 10600 9948
rect 10652 9936 10658 9988
rect 10796 9976 10824 10007
rect 10704 9948 10824 9976
rect 12406 9976 12434 10152
rect 14752 10152 15792 10180
rect 14366 10072 14372 10124
rect 14424 10112 14430 10124
rect 14752 10121 14780 10152
rect 14553 10115 14611 10121
rect 14553 10112 14565 10115
rect 14424 10084 14565 10112
rect 14424 10072 14430 10084
rect 14553 10081 14565 10084
rect 14599 10081 14611 10115
rect 14553 10075 14611 10081
rect 14737 10115 14795 10121
rect 14737 10081 14749 10115
rect 14783 10081 14795 10115
rect 14737 10075 14795 10081
rect 15654 10072 15660 10124
rect 15712 10072 15718 10124
rect 15764 10112 15792 10152
rect 18414 10112 18420 10124
rect 15764 10084 18420 10112
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 19889 10115 19947 10121
rect 19889 10081 19901 10115
rect 19935 10112 19947 10115
rect 20254 10112 20260 10124
rect 19935 10084 20260 10112
rect 19935 10081 19947 10084
rect 19889 10075 19947 10081
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 23842 10112 23848 10124
rect 21468 10084 23848 10112
rect 14918 10004 14924 10056
rect 14976 10004 14982 10056
rect 17218 10044 17224 10056
rect 17066 10016 17224 10044
rect 17218 10004 17224 10016
rect 17276 10004 17282 10056
rect 21468 9988 21496 10084
rect 23842 10072 23848 10084
rect 23900 10072 23906 10124
rect 24228 10112 24256 10208
rect 24228 10084 25636 10112
rect 21818 10004 21824 10056
rect 21876 10004 21882 10056
rect 22005 10047 22063 10053
rect 22005 10013 22017 10047
rect 22051 10044 22063 10047
rect 22370 10044 22376 10056
rect 22051 10016 22376 10044
rect 22051 10013 22063 10016
rect 22005 10007 22063 10013
rect 22370 10004 22376 10016
rect 22428 10004 22434 10056
rect 24210 10004 24216 10056
rect 24268 10044 24274 10056
rect 25130 10044 25136 10056
rect 24268 10016 25136 10044
rect 24268 10004 24274 10016
rect 25130 10004 25136 10016
rect 25188 10004 25194 10056
rect 25608 10053 25636 10084
rect 25593 10047 25651 10053
rect 25593 10013 25605 10047
rect 25639 10013 25651 10047
rect 25593 10007 25651 10013
rect 25866 10004 25872 10056
rect 25924 10004 25930 10056
rect 21450 9976 21456 9988
rect 12406 9948 16344 9976
rect 21390 9948 21456 9976
rect 10704 9920 10732 9948
rect 10686 9908 10692 9920
rect 9508 9880 10692 9908
rect 9217 9871 9275 9877
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 13998 9868 14004 9920
rect 14056 9908 14062 9920
rect 14093 9911 14151 9917
rect 14093 9908 14105 9911
rect 14056 9880 14105 9908
rect 14056 9868 14062 9880
rect 14093 9877 14105 9880
rect 14139 9877 14151 9911
rect 14093 9871 14151 9877
rect 14461 9911 14519 9917
rect 14461 9877 14473 9911
rect 14507 9908 14519 9911
rect 14642 9908 14648 9920
rect 14507 9880 14648 9908
rect 14507 9877 14519 9880
rect 14461 9871 14519 9877
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 15105 9911 15163 9917
rect 15105 9877 15117 9911
rect 15151 9908 15163 9911
rect 15286 9908 15292 9920
rect 15151 9880 15292 9908
rect 15151 9877 15163 9880
rect 15105 9871 15163 9877
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 16316 9908 16344 9948
rect 21450 9936 21456 9948
rect 21508 9936 21514 9988
rect 23842 9976 23848 9988
rect 23506 9948 23848 9976
rect 23842 9936 23848 9948
rect 23900 9936 23906 9988
rect 23934 9936 23940 9988
rect 23992 9936 23998 9988
rect 24397 9979 24455 9985
rect 24397 9945 24409 9979
rect 24443 9945 24455 9979
rect 24397 9939 24455 9945
rect 17218 9908 17224 9920
rect 16316 9880 17224 9908
rect 17218 9868 17224 9880
rect 17276 9868 17282 9920
rect 17310 9868 17316 9920
rect 17368 9908 17374 9920
rect 17405 9911 17463 9917
rect 17405 9908 17417 9911
rect 17368 9880 17417 9908
rect 17368 9868 17374 9880
rect 17405 9877 17417 9880
rect 17451 9877 17463 9911
rect 17405 9871 17463 9877
rect 21174 9868 21180 9920
rect 21232 9908 21238 9920
rect 21637 9911 21695 9917
rect 21637 9908 21649 9911
rect 21232 9880 21649 9908
rect 21232 9868 21238 9880
rect 21637 9877 21649 9880
rect 21683 9877 21695 9911
rect 21637 9871 21695 9877
rect 22646 9868 22652 9920
rect 22704 9908 22710 9920
rect 24412 9908 24440 9939
rect 25498 9936 25504 9988
rect 25556 9976 25562 9988
rect 25777 9979 25835 9985
rect 25777 9976 25789 9979
rect 25556 9948 25789 9976
rect 25556 9936 25562 9948
rect 25777 9945 25789 9948
rect 25823 9945 25835 9979
rect 25777 9939 25835 9945
rect 22704 9880 24440 9908
rect 22704 9868 22710 9880
rect 1104 9818 26472 9840
rect 1104 9766 7252 9818
rect 7304 9766 7316 9818
rect 7368 9766 7380 9818
rect 7432 9766 7444 9818
rect 7496 9766 7508 9818
rect 7560 9766 13554 9818
rect 13606 9766 13618 9818
rect 13670 9766 13682 9818
rect 13734 9766 13746 9818
rect 13798 9766 13810 9818
rect 13862 9766 19856 9818
rect 19908 9766 19920 9818
rect 19972 9766 19984 9818
rect 20036 9766 20048 9818
rect 20100 9766 20112 9818
rect 20164 9766 26158 9818
rect 26210 9766 26222 9818
rect 26274 9766 26286 9818
rect 26338 9766 26350 9818
rect 26402 9766 26414 9818
rect 26466 9766 26472 9818
rect 1104 9744 26472 9766
rect 3970 9664 3976 9716
rect 4028 9704 4034 9716
rect 4706 9704 4712 9716
rect 4028 9676 4712 9704
rect 4028 9664 4034 9676
rect 2222 9596 2228 9648
rect 2280 9636 2286 9648
rect 2317 9639 2375 9645
rect 2317 9636 2329 9639
rect 2280 9608 2329 9636
rect 2280 9596 2286 9608
rect 2317 9605 2329 9608
rect 2363 9605 2375 9639
rect 2317 9599 2375 9605
rect 2590 9596 2596 9648
rect 2648 9636 2654 9648
rect 3237 9639 3295 9645
rect 3237 9636 3249 9639
rect 2648 9608 3249 9636
rect 2648 9596 2654 9608
rect 3237 9605 3249 9608
rect 3283 9605 3295 9639
rect 3237 9599 3295 9605
rect 2041 9571 2099 9577
rect 2041 9537 2053 9571
rect 2087 9568 2099 9571
rect 2866 9568 2872 9580
rect 2087 9540 2872 9568
rect 2087 9537 2099 9540
rect 2041 9531 2099 9537
rect 2866 9528 2872 9540
rect 2924 9568 2930 9580
rect 2961 9571 3019 9577
rect 2961 9568 2973 9571
rect 2924 9540 2973 9568
rect 2924 9528 2930 9540
rect 2961 9537 2973 9540
rect 3007 9537 3019 9571
rect 2961 9531 3019 9537
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9500 2375 9503
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2363 9472 2697 9500
rect 2363 9469 2375 9472
rect 2317 9463 2375 9469
rect 2685 9469 2697 9472
rect 2731 9500 2743 9503
rect 3142 9500 3148 9512
rect 2731 9472 3148 9500
rect 2731 9469 2743 9472
rect 2685 9463 2743 9469
rect 3142 9460 3148 9472
rect 3200 9460 3206 9512
rect 1762 9392 1768 9444
rect 1820 9432 1826 9444
rect 2777 9435 2835 9441
rect 2777 9432 2789 9435
rect 1820 9404 2789 9432
rect 1820 9392 1826 9404
rect 2777 9401 2789 9404
rect 2823 9401 2835 9435
rect 3252 9432 3280 9599
rect 3878 9596 3884 9648
rect 3936 9596 3942 9648
rect 4341 9639 4399 9645
rect 4341 9614 4353 9639
rect 4387 9614 4399 9639
rect 3970 9528 3976 9580
rect 4028 9568 4034 9580
rect 4065 9571 4123 9577
rect 4065 9568 4077 9571
rect 4028 9540 4077 9568
rect 4028 9528 4034 9540
rect 4065 9537 4077 9540
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 4154 9528 4160 9580
rect 4212 9568 4218 9580
rect 4212 9540 4292 9568
rect 4338 9562 4344 9614
rect 4396 9562 4402 9614
rect 4448 9577 4476 9676
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 6730 9664 6736 9716
rect 6788 9664 6794 9716
rect 6914 9664 6920 9716
rect 6972 9704 6978 9716
rect 7650 9704 7656 9716
rect 6972 9676 7656 9704
rect 6972 9664 6978 9676
rect 7650 9664 7656 9676
rect 7708 9664 7714 9716
rect 8665 9707 8723 9713
rect 8665 9673 8677 9707
rect 8711 9704 8723 9707
rect 8754 9704 8760 9716
rect 8711 9676 8760 9704
rect 8711 9673 8723 9676
rect 8665 9667 8723 9673
rect 8754 9664 8760 9676
rect 8812 9664 8818 9716
rect 8846 9664 8852 9716
rect 8904 9704 8910 9716
rect 9125 9707 9183 9713
rect 9125 9704 9137 9707
rect 8904 9676 9137 9704
rect 8904 9664 8910 9676
rect 9125 9673 9137 9676
rect 9171 9673 9183 9707
rect 9125 9667 9183 9673
rect 9582 9664 9588 9716
rect 9640 9664 9646 9716
rect 9674 9664 9680 9716
rect 9732 9704 9738 9716
rect 10137 9707 10195 9713
rect 10137 9704 10149 9707
rect 9732 9676 10149 9704
rect 9732 9664 9738 9676
rect 10137 9673 10149 9676
rect 10183 9673 10195 9707
rect 10137 9667 10195 9673
rect 10686 9664 10692 9716
rect 10744 9664 10750 9716
rect 10778 9664 10784 9716
rect 10836 9704 10842 9716
rect 10873 9707 10931 9713
rect 10873 9704 10885 9707
rect 10836 9676 10885 9704
rect 10836 9664 10842 9676
rect 10873 9673 10885 9676
rect 10919 9673 10931 9707
rect 10873 9667 10931 9673
rect 14366 9664 14372 9716
rect 14424 9664 14430 9716
rect 14829 9707 14887 9713
rect 14829 9673 14841 9707
rect 14875 9704 14887 9707
rect 14918 9704 14924 9716
rect 14875 9676 14924 9704
rect 14875 9673 14887 9676
rect 14829 9667 14887 9673
rect 14918 9664 14924 9676
rect 14976 9664 14982 9716
rect 17126 9664 17132 9716
rect 17184 9664 17190 9716
rect 17218 9664 17224 9716
rect 17276 9704 17282 9716
rect 22830 9704 22836 9716
rect 17276 9676 22836 9704
rect 17276 9664 17282 9676
rect 22830 9664 22836 9676
rect 22888 9664 22894 9716
rect 23431 9707 23489 9713
rect 23431 9673 23443 9707
rect 23477 9704 23489 9707
rect 24394 9704 24400 9716
rect 23477 9676 24400 9704
rect 23477 9673 23489 9676
rect 23431 9667 23489 9673
rect 24394 9664 24400 9676
rect 24452 9664 24458 9716
rect 25866 9664 25872 9716
rect 25924 9664 25930 9716
rect 4433 9571 4491 9577
rect 4212 9528 4218 9540
rect 3326 9460 3332 9512
rect 3384 9500 3390 9512
rect 3384 9472 4200 9500
rect 3384 9460 3390 9472
rect 4172 9441 4200 9472
rect 3605 9435 3663 9441
rect 3252 9404 3372 9432
rect 2777 9395 2835 9401
rect 2130 9324 2136 9376
rect 2188 9324 2194 9376
rect 2869 9367 2927 9373
rect 2869 9333 2881 9367
rect 2915 9364 2927 9367
rect 2958 9364 2964 9376
rect 2915 9336 2964 9364
rect 2915 9333 2927 9336
rect 2869 9327 2927 9333
rect 2958 9324 2964 9336
rect 3016 9364 3022 9376
rect 3053 9367 3111 9373
rect 3053 9364 3065 9367
rect 3016 9336 3065 9364
rect 3016 9324 3022 9336
rect 3053 9333 3065 9336
rect 3099 9333 3111 9367
rect 3053 9327 3111 9333
rect 3234 9324 3240 9376
rect 3292 9324 3298 9376
rect 3344 9364 3372 9404
rect 3605 9401 3617 9435
rect 3651 9432 3663 9435
rect 4157 9435 4215 9441
rect 3651 9404 4016 9432
rect 3651 9401 3663 9404
rect 3605 9395 3663 9401
rect 3988 9376 4016 9404
rect 4157 9401 4169 9435
rect 4203 9401 4215 9435
rect 4157 9395 4215 9401
rect 3694 9364 3700 9376
rect 3344 9336 3700 9364
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 3970 9324 3976 9376
rect 4028 9324 4034 9376
rect 4264 9364 4292 9540
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 4522 9528 4528 9580
rect 4580 9528 4586 9580
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 4798 9568 4804 9580
rect 4755 9540 4804 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 6748 9577 6776 9664
rect 9600 9636 9628 9664
rect 9953 9639 10011 9645
rect 9600 9608 9720 9636
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9537 6791 9571
rect 6733 9531 6791 9537
rect 6822 9528 6828 9580
rect 6880 9528 6886 9580
rect 8478 9528 8484 9580
rect 8536 9528 8542 9580
rect 8662 9528 8668 9580
rect 8720 9568 8726 9580
rect 9692 9577 9720 9608
rect 9953 9605 9965 9639
rect 9999 9605 10011 9639
rect 9953 9599 10011 9605
rect 8849 9571 8907 9577
rect 8849 9568 8861 9571
rect 8720 9540 8861 9568
rect 8720 9528 8726 9540
rect 8849 9537 8861 9540
rect 8895 9537 8907 9571
rect 8849 9531 8907 9537
rect 9677 9571 9735 9577
rect 9677 9537 9689 9571
rect 9723 9537 9735 9571
rect 9677 9531 9735 9537
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9568 9827 9571
rect 9858 9568 9864 9580
rect 9815 9540 9864 9568
rect 9815 9537 9827 9540
rect 9769 9531 9827 9537
rect 9858 9528 9864 9540
rect 9916 9528 9922 9580
rect 9968 9568 9996 9599
rect 10042 9596 10048 9648
rect 10100 9636 10106 9648
rect 10962 9636 10968 9648
rect 10100 9608 10968 9636
rect 10100 9596 10106 9608
rect 10962 9596 10968 9608
rect 11020 9636 11026 9648
rect 14384 9636 14412 9664
rect 15289 9639 15347 9645
rect 15289 9636 15301 9639
rect 11020 9608 12434 9636
rect 14384 9608 15301 9636
rect 11020 9596 11026 9608
rect 10134 9568 10140 9580
rect 9968 9540 10140 9568
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 10318 9528 10324 9580
rect 10376 9528 10382 9580
rect 10410 9528 10416 9580
rect 10468 9568 10474 9580
rect 11146 9577 11152 9580
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 10468 9540 10793 9568
rect 10468 9528 10474 9540
rect 10781 9537 10793 9540
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 10873 9571 10931 9577
rect 10873 9537 10885 9571
rect 10919 9537 10931 9571
rect 11050 9571 11108 9577
rect 11050 9566 11062 9571
rect 10873 9531 10931 9537
rect 10980 9538 11062 9566
rect 6641 9503 6699 9509
rect 6641 9469 6653 9503
rect 6687 9500 6699 9503
rect 6840 9500 6868 9528
rect 6687 9472 6868 9500
rect 8496 9500 8524 9528
rect 8941 9503 8999 9509
rect 8941 9500 8953 9503
rect 8496 9472 8953 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 8941 9469 8953 9472
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 9953 9503 10011 9509
rect 9953 9469 9965 9503
rect 9999 9500 10011 9503
rect 10333 9500 10361 9528
rect 9999 9472 10361 9500
rect 10505 9503 10563 9509
rect 9999 9469 10011 9472
rect 9953 9463 10011 9469
rect 10505 9469 10517 9503
rect 10551 9500 10563 9503
rect 10594 9500 10600 9512
rect 10551 9472 10600 9500
rect 10551 9469 10563 9472
rect 10505 9463 10563 9469
rect 5810 9392 5816 9444
rect 5868 9432 5874 9444
rect 6365 9435 6423 9441
rect 6365 9432 6377 9435
rect 5868 9404 6377 9432
rect 5868 9392 5874 9404
rect 6365 9401 6377 9404
rect 6411 9401 6423 9435
rect 9140 9432 9168 9463
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 10888 9444 10916 9531
rect 10870 9432 10876 9444
rect 9140 9404 10876 9432
rect 6365 9395 6423 9401
rect 10870 9392 10876 9404
rect 10928 9392 10934 9444
rect 10980 9432 11008 9538
rect 11050 9537 11062 9538
rect 11096 9537 11108 9571
rect 11050 9531 11108 9537
rect 11137 9571 11152 9577
rect 11137 9537 11149 9571
rect 11137 9531 11152 9537
rect 11146 9528 11152 9531
rect 11204 9528 11210 9580
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9537 11391 9571
rect 12406 9568 12434 9608
rect 15289 9605 15301 9608
rect 15335 9605 15347 9639
rect 15289 9599 15347 9605
rect 16945 9639 17003 9645
rect 16945 9605 16957 9639
rect 16991 9636 17003 9639
rect 17034 9636 17040 9648
rect 16991 9608 17040 9636
rect 16991 9605 17003 9608
rect 16945 9599 17003 9605
rect 17034 9596 17040 9608
rect 17092 9596 17098 9648
rect 17144 9636 17172 9664
rect 17144 9608 17434 9636
rect 19702 9596 19708 9648
rect 19760 9636 19766 9648
rect 20809 9639 20867 9645
rect 20809 9636 20821 9639
rect 19760 9608 20821 9636
rect 19760 9596 19766 9608
rect 20809 9605 20821 9608
rect 20855 9605 20867 9639
rect 20809 9599 20867 9605
rect 23842 9596 23848 9648
rect 23900 9596 23906 9648
rect 25314 9596 25320 9648
rect 25372 9596 25378 9648
rect 12713 9571 12771 9577
rect 12713 9568 12725 9571
rect 12406 9540 12725 9568
rect 11333 9531 11391 9537
rect 12713 9537 12725 9540
rect 12759 9537 12771 9571
rect 12713 9531 12771 9537
rect 11054 9432 11060 9444
rect 10980 9404 11060 9432
rect 11054 9392 11060 9404
rect 11112 9392 11118 9444
rect 11149 9435 11207 9441
rect 11149 9401 11161 9435
rect 11195 9401 11207 9435
rect 11149 9395 11207 9401
rect 4522 9364 4528 9376
rect 4264 9336 4528 9364
rect 4522 9324 4528 9336
rect 4580 9324 4586 9376
rect 4614 9324 4620 9376
rect 4672 9364 4678 9376
rect 4709 9367 4767 9373
rect 4709 9364 4721 9367
rect 4672 9336 4721 9364
rect 4672 9324 4678 9336
rect 4709 9333 4721 9336
rect 4755 9333 4767 9367
rect 4709 9327 4767 9333
rect 5626 9324 5632 9376
rect 5684 9364 5690 9376
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 5684 9336 6561 9364
rect 5684 9324 5690 9336
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 6549 9327 6607 9333
rect 10410 9324 10416 9376
rect 10468 9364 10474 9376
rect 11164 9364 11192 9395
rect 11348 9376 11376 9531
rect 14090 9528 14096 9580
rect 14148 9568 14154 9580
rect 15102 9568 15108 9580
rect 14148 9540 15108 9568
rect 14148 9528 14154 9540
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 15194 9528 15200 9580
rect 15252 9528 15258 9580
rect 16022 9528 16028 9580
rect 16080 9568 16086 9580
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 16080 9540 16681 9568
rect 16080 9528 16086 9540
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 22646 9568 22652 9580
rect 16669 9531 16727 9537
rect 18524 9540 22652 9568
rect 12986 9460 12992 9512
rect 13044 9460 13050 9512
rect 14642 9460 14648 9512
rect 14700 9500 14706 9512
rect 14737 9503 14795 9509
rect 14737 9500 14749 9503
rect 14700 9472 14749 9500
rect 14700 9460 14706 9472
rect 14737 9469 14749 9472
rect 14783 9469 14795 9503
rect 14737 9463 14795 9469
rect 15473 9503 15531 9509
rect 15473 9469 15485 9503
rect 15519 9500 15531 9503
rect 15519 9472 16436 9500
rect 15519 9469 15531 9472
rect 15473 9463 15531 9469
rect 16408 9376 16436 9472
rect 17586 9460 17592 9512
rect 17644 9500 17650 9512
rect 18524 9500 18552 9540
rect 22646 9528 22652 9540
rect 22704 9528 22710 9580
rect 24857 9571 24915 9577
rect 24857 9537 24869 9571
rect 24903 9568 24915 9571
rect 24946 9568 24952 9580
rect 24903 9540 24952 9568
rect 24903 9537 24915 9540
rect 24857 9531 24915 9537
rect 24946 9528 24952 9540
rect 25004 9528 25010 9580
rect 25130 9528 25136 9580
rect 25188 9568 25194 9580
rect 25225 9571 25283 9577
rect 25225 9568 25237 9571
rect 25188 9540 25237 9568
rect 25188 9528 25194 9540
rect 25225 9537 25237 9540
rect 25271 9537 25283 9571
rect 25332 9568 25360 9596
rect 25409 9571 25467 9577
rect 25409 9568 25421 9571
rect 25332 9540 25421 9568
rect 25225 9531 25283 9537
rect 25409 9537 25421 9540
rect 25455 9537 25467 9571
rect 25409 9531 25467 9537
rect 17644 9472 18552 9500
rect 18601 9503 18659 9509
rect 17644 9460 17650 9472
rect 18601 9469 18613 9503
rect 18647 9469 18659 9503
rect 18601 9463 18659 9469
rect 18616 9432 18644 9463
rect 19610 9460 19616 9512
rect 19668 9500 19674 9512
rect 19889 9503 19947 9509
rect 19889 9500 19901 9503
rect 19668 9472 19901 9500
rect 19668 9460 19674 9472
rect 19889 9469 19901 9472
rect 19935 9500 19947 9503
rect 20625 9503 20683 9509
rect 20625 9500 20637 9503
rect 19935 9472 20637 9500
rect 19935 9469 19947 9472
rect 19889 9463 19947 9469
rect 20625 9469 20637 9472
rect 20671 9469 20683 9503
rect 20625 9463 20683 9469
rect 21082 9460 21088 9512
rect 21140 9500 21146 9512
rect 21361 9503 21419 9509
rect 21361 9500 21373 9503
rect 21140 9472 21373 9500
rect 21140 9460 21146 9472
rect 21361 9469 21373 9472
rect 21407 9469 21419 9503
rect 22373 9503 22431 9509
rect 22373 9500 22385 9503
rect 21361 9463 21419 9469
rect 22066 9472 22385 9500
rect 18432 9404 18644 9432
rect 10468 9336 11192 9364
rect 10468 9324 10474 9336
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 13722 9364 13728 9376
rect 11388 9336 13728 9364
rect 11388 9324 11394 9336
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 16390 9324 16396 9376
rect 16448 9324 16454 9376
rect 17678 9324 17684 9376
rect 17736 9364 17742 9376
rect 18432 9373 18460 9404
rect 18966 9392 18972 9444
rect 19024 9432 19030 9444
rect 19337 9435 19395 9441
rect 19337 9432 19349 9435
rect 19024 9404 19349 9432
rect 19024 9392 19030 9404
rect 19337 9401 19349 9404
rect 19383 9401 19395 9435
rect 19337 9395 19395 9401
rect 21174 9392 21180 9444
rect 21232 9432 21238 9444
rect 22066 9432 22094 9472
rect 22373 9469 22385 9472
rect 22419 9469 22431 9503
rect 22373 9463 22431 9469
rect 21232 9404 22094 9432
rect 21232 9392 21238 9404
rect 18417 9367 18475 9373
rect 18417 9364 18429 9367
rect 17736 9336 18429 9364
rect 17736 9324 17742 9336
rect 18417 9333 18429 9336
rect 18463 9333 18475 9367
rect 18417 9327 18475 9333
rect 19242 9324 19248 9376
rect 19300 9324 19306 9376
rect 19610 9324 19616 9376
rect 19668 9364 19674 9376
rect 20073 9367 20131 9373
rect 20073 9364 20085 9367
rect 19668 9336 20085 9364
rect 19668 9324 19674 9336
rect 20073 9333 20085 9336
rect 20119 9333 20131 9367
rect 20073 9327 20131 9333
rect 21634 9324 21640 9376
rect 21692 9364 21698 9376
rect 21821 9367 21879 9373
rect 21821 9364 21833 9367
rect 21692 9336 21833 9364
rect 21692 9324 21698 9336
rect 21821 9333 21833 9336
rect 21867 9333 21879 9367
rect 21821 9327 21879 9333
rect 25682 9324 25688 9376
rect 25740 9324 25746 9376
rect 1104 9274 26312 9296
rect 1104 9222 4101 9274
rect 4153 9222 4165 9274
rect 4217 9222 4229 9274
rect 4281 9222 4293 9274
rect 4345 9222 4357 9274
rect 4409 9222 10403 9274
rect 10455 9222 10467 9274
rect 10519 9222 10531 9274
rect 10583 9222 10595 9274
rect 10647 9222 10659 9274
rect 10711 9222 16705 9274
rect 16757 9222 16769 9274
rect 16821 9222 16833 9274
rect 16885 9222 16897 9274
rect 16949 9222 16961 9274
rect 17013 9222 23007 9274
rect 23059 9222 23071 9274
rect 23123 9222 23135 9274
rect 23187 9222 23199 9274
rect 23251 9222 23263 9274
rect 23315 9222 26312 9274
rect 1104 9200 26312 9222
rect 2682 9120 2688 9172
rect 2740 9160 2746 9172
rect 3234 9160 3240 9172
rect 2740 9132 3240 9160
rect 2740 9120 2746 9132
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 3878 9120 3884 9172
rect 3936 9160 3942 9172
rect 4430 9160 4436 9172
rect 3936 9132 4436 9160
rect 3936 9120 3942 9132
rect 4430 9120 4436 9132
rect 4488 9160 4494 9172
rect 5629 9163 5687 9169
rect 5629 9160 5641 9163
rect 4488 9132 5641 9160
rect 4488 9120 4494 9132
rect 5629 9129 5641 9132
rect 5675 9129 5687 9163
rect 5629 9123 5687 9129
rect 6546 9120 6552 9172
rect 6604 9160 6610 9172
rect 6733 9163 6791 9169
rect 6733 9160 6745 9163
rect 6604 9132 6745 9160
rect 6604 9120 6610 9132
rect 6733 9129 6745 9132
rect 6779 9129 6791 9163
rect 8478 9160 8484 9172
rect 6733 9123 6791 9129
rect 7484 9132 8484 9160
rect 4246 9092 4252 9104
rect 3988 9064 4252 9092
rect 1673 9027 1731 9033
rect 1673 8993 1685 9027
rect 1719 9024 1731 9027
rect 2406 9024 2412 9036
rect 1719 8996 2412 9024
rect 1719 8993 1731 8996
rect 1673 8987 1731 8993
rect 2406 8984 2412 8996
rect 2464 8984 2470 9036
rect 2866 8984 2872 9036
rect 2924 9024 2930 9036
rect 3421 9027 3479 9033
rect 3421 9024 3433 9027
rect 2924 8996 3433 9024
rect 2924 8984 2930 8996
rect 3421 8993 3433 8996
rect 3467 9024 3479 9027
rect 3988 9024 4016 9064
rect 4246 9052 4252 9064
rect 4304 9092 4310 9104
rect 5258 9092 5264 9104
rect 4304 9064 5264 9092
rect 4304 9052 4310 9064
rect 5258 9052 5264 9064
rect 5316 9052 5322 9104
rect 7484 9101 7512 9132
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 9398 9120 9404 9172
rect 9456 9160 9462 9172
rect 10137 9163 10195 9169
rect 10137 9160 10149 9163
rect 9456 9132 10149 9160
rect 9456 9120 9462 9132
rect 10137 9129 10149 9132
rect 10183 9129 10195 9163
rect 10137 9123 10195 9129
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 11330 9160 11336 9172
rect 10928 9132 11336 9160
rect 10928 9120 10934 9132
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 13265 9163 13323 9169
rect 13265 9160 13277 9163
rect 13044 9132 13277 9160
rect 13044 9120 13050 9132
rect 13265 9129 13277 9132
rect 13311 9129 13323 9163
rect 13265 9123 13323 9129
rect 13924 9132 14688 9160
rect 7469 9095 7527 9101
rect 7469 9061 7481 9095
rect 7515 9061 7527 9095
rect 7742 9092 7748 9104
rect 7469 9055 7527 9061
rect 7576 9064 7748 9092
rect 3467 8996 4016 9024
rect 3467 8993 3479 8996
rect 3421 8987 3479 8993
rect 1394 8916 1400 8968
rect 1452 8916 1458 8968
rect 2774 8916 2780 8968
rect 2832 8916 2838 8968
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8956 3847 8959
rect 3878 8956 3884 8968
rect 3835 8928 3884 8956
rect 3835 8925 3847 8928
rect 3789 8919 3847 8925
rect 3878 8916 3884 8928
rect 3936 8916 3942 8968
rect 3988 8965 4016 8996
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 4890 9024 4896 9036
rect 4479 8996 4896 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 7576 9024 7604 9064
rect 7742 9052 7748 9064
rect 7800 9052 7806 9104
rect 8205 9095 8263 9101
rect 8205 9061 8217 9095
rect 8251 9092 8263 9095
rect 8662 9092 8668 9104
rect 8251 9064 8668 9092
rect 8251 9061 8263 9064
rect 8205 9055 8263 9061
rect 8662 9052 8668 9064
rect 8720 9052 8726 9104
rect 8754 9052 8760 9104
rect 8812 9092 8818 9104
rect 13924 9092 13952 9132
rect 14660 9104 14688 9132
rect 15102 9120 15108 9172
rect 15160 9160 15166 9172
rect 17954 9160 17960 9172
rect 15160 9132 17960 9160
rect 15160 9120 15166 9132
rect 17954 9120 17960 9132
rect 18012 9120 18018 9172
rect 19242 9120 19248 9172
rect 19300 9120 19306 9172
rect 8812 9064 13952 9092
rect 8812 9052 8818 9064
rect 13998 9052 14004 9104
rect 14056 9052 14062 9104
rect 14642 9052 14648 9104
rect 14700 9052 14706 9104
rect 16390 9052 16396 9104
rect 16448 9092 16454 9104
rect 19260 9092 19288 9120
rect 16448 9064 18552 9092
rect 16448 9052 16454 9064
rect 5000 8996 5212 9024
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 4249 8959 4307 8965
rect 4249 8956 4261 8959
rect 4212 8928 4261 8956
rect 4212 8916 4218 8928
rect 4249 8925 4261 8928
rect 4295 8956 4307 8959
rect 4614 8956 4620 8968
rect 4295 8928 4620 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 4706 8916 4712 8968
rect 4764 8916 4770 8968
rect 4798 8916 4804 8968
rect 4856 8956 4862 8968
rect 5000 8956 5028 8996
rect 4856 8928 5028 8956
rect 5077 8959 5135 8965
rect 4856 8916 4862 8928
rect 5077 8925 5089 8959
rect 5123 8925 5135 8959
rect 5077 8919 5135 8925
rect 4062 8848 4068 8900
rect 4120 8888 4126 8900
rect 4525 8891 4583 8897
rect 4525 8888 4537 8891
rect 4120 8860 4537 8888
rect 4120 8848 4126 8860
rect 4525 8857 4537 8860
rect 4571 8857 4583 8891
rect 4632 8888 4660 8916
rect 5092 8888 5120 8919
rect 4632 8860 5120 8888
rect 5184 8888 5212 8996
rect 6840 8996 7604 9024
rect 7653 9027 7711 9033
rect 5258 8916 5264 8968
rect 5316 8916 5322 8968
rect 6840 8965 6868 8996
rect 7653 8993 7665 9027
rect 7699 9024 7711 9027
rect 8772 9024 8800 9052
rect 11885 9027 11943 9033
rect 7699 8996 8800 9024
rect 9646 8996 10364 9024
rect 7699 8993 7711 8996
rect 7653 8987 7711 8993
rect 7944 8965 7972 8996
rect 5537 8959 5595 8965
rect 5537 8956 5549 8959
rect 5368 8928 5549 8956
rect 5368 8888 5396 8928
rect 5537 8925 5549 8928
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 6825 8959 6883 8965
rect 6825 8925 6837 8959
rect 6871 8925 6883 8959
rect 6825 8919 6883 8925
rect 7469 8959 7527 8965
rect 7469 8925 7481 8959
rect 7515 8956 7527 8959
rect 7745 8959 7803 8965
rect 7745 8956 7757 8959
rect 7515 8928 7757 8956
rect 7515 8925 7527 8928
rect 7469 8919 7527 8925
rect 7745 8925 7757 8928
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8925 7987 8959
rect 7929 8919 7987 8925
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8956 8355 8959
rect 8386 8956 8392 8968
rect 8343 8928 8392 8956
rect 8343 8925 8355 8928
rect 8297 8919 8355 8925
rect 5184 8860 5396 8888
rect 5445 8891 5503 8897
rect 4525 8851 4583 8857
rect 5445 8857 5457 8891
rect 5491 8857 5503 8891
rect 6656 8888 6684 8919
rect 7098 8888 7104 8900
rect 6656 8860 7104 8888
rect 5445 8851 5503 8857
rect 3786 8780 3792 8832
rect 3844 8820 3850 8832
rect 5460 8820 5488 8851
rect 7098 8848 7104 8860
rect 7156 8848 7162 8900
rect 3844 8792 5488 8820
rect 3844 8780 3850 8792
rect 6730 8780 6736 8832
rect 6788 8820 6794 8832
rect 7484 8820 7512 8919
rect 8386 8916 8392 8928
rect 8444 8956 8450 8968
rect 9646 8956 9674 8996
rect 8444 8928 9674 8956
rect 8444 8916 8450 8928
rect 9950 8916 9956 8968
rect 10008 8956 10014 8968
rect 10045 8959 10103 8965
rect 10045 8956 10057 8959
rect 10008 8928 10057 8956
rect 10008 8916 10014 8928
rect 10045 8925 10057 8928
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10336 8956 10364 8996
rect 11885 8993 11897 9027
rect 11931 9024 11943 9027
rect 12066 9024 12072 9036
rect 11931 8996 12072 9024
rect 11931 8993 11943 8996
rect 11885 8987 11943 8993
rect 12066 8984 12072 8996
rect 12124 8984 12130 9036
rect 13449 8959 13507 8965
rect 10336 8928 13400 8956
rect 10229 8919 10287 8925
rect 6788 8792 7512 8820
rect 10060 8820 10088 8919
rect 10244 8888 10272 8919
rect 10318 8888 10324 8900
rect 10244 8860 10324 8888
rect 10318 8848 10324 8860
rect 10376 8888 10382 8900
rect 10870 8888 10876 8900
rect 10376 8860 10876 8888
rect 10376 8848 10382 8860
rect 10870 8848 10876 8860
rect 10928 8848 10934 8900
rect 11241 8823 11299 8829
rect 11241 8820 11253 8823
rect 10060 8792 11253 8820
rect 6788 8780 6794 8792
rect 11241 8789 11253 8792
rect 11287 8789 11299 8823
rect 11241 8783 11299 8789
rect 11606 8780 11612 8832
rect 11664 8780 11670 8832
rect 11701 8823 11759 8829
rect 11701 8789 11713 8823
rect 11747 8820 11759 8823
rect 11790 8820 11796 8832
rect 11747 8792 11796 8820
rect 11747 8789 11759 8792
rect 11701 8783 11759 8789
rect 11790 8780 11796 8792
rect 11848 8820 11854 8832
rect 12342 8820 12348 8832
rect 11848 8792 12348 8820
rect 11848 8780 11854 8792
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 13372 8820 13400 8928
rect 13449 8925 13461 8959
rect 13495 8956 13507 8959
rect 14016 8956 14044 9052
rect 14185 9027 14243 9033
rect 14185 8993 14197 9027
rect 14231 9024 14243 9027
rect 15194 9024 15200 9036
rect 14231 8996 15200 9024
rect 14231 8993 14243 8996
rect 14185 8987 14243 8993
rect 15194 8984 15200 8996
rect 15252 8984 15258 9036
rect 15286 8984 15292 9036
rect 15344 9024 15350 9036
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 15344 8996 15669 9024
rect 15344 8984 15350 8996
rect 15657 8993 15669 8996
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 9024 15991 9027
rect 16022 9024 16028 9036
rect 15979 8996 16028 9024
rect 15979 8993 15991 8996
rect 15933 8987 15991 8993
rect 16022 8984 16028 8996
rect 16080 8984 16086 9036
rect 16684 9033 16712 9064
rect 18524 9036 18552 9064
rect 18616 9064 19288 9092
rect 16669 9027 16727 9033
rect 16669 8993 16681 9027
rect 16715 8993 16727 9027
rect 16669 8987 16727 8993
rect 16761 9027 16819 9033
rect 16761 8993 16773 9027
rect 16807 9024 16819 9027
rect 17678 9024 17684 9036
rect 16807 8996 17684 9024
rect 16807 8993 16819 8996
rect 16761 8987 16819 8993
rect 17678 8984 17684 8996
rect 17736 8984 17742 9036
rect 18414 8984 18420 9036
rect 18472 8984 18478 9036
rect 18506 8984 18512 9036
rect 18564 8984 18570 9036
rect 18616 9033 18644 9064
rect 18601 9027 18659 9033
rect 18601 8993 18613 9027
rect 18647 8993 18659 9027
rect 20165 9027 20223 9033
rect 20165 9024 20177 9027
rect 18601 8987 18659 8993
rect 19260 8996 20177 9024
rect 13495 8928 14044 8956
rect 16040 8956 16068 8984
rect 17034 8956 17040 8968
rect 16040 8928 17040 8956
rect 13495 8925 13507 8928
rect 13449 8919 13507 8925
rect 17034 8916 17040 8928
rect 17092 8956 17098 8968
rect 18049 8959 18107 8965
rect 18049 8956 18061 8959
rect 17092 8928 18061 8956
rect 17092 8916 17098 8928
rect 18049 8925 18061 8928
rect 18095 8925 18107 8959
rect 18432 8956 18460 8984
rect 19260 8968 19288 8996
rect 20165 8993 20177 8996
rect 20211 8993 20223 9027
rect 20165 8987 20223 8993
rect 22281 9027 22339 9033
rect 22281 8993 22293 9027
rect 22327 9024 22339 9027
rect 22327 8996 24256 9024
rect 22327 8993 22339 8996
rect 22281 8987 22339 8993
rect 24228 8968 24256 8996
rect 18432 8928 18644 8956
rect 18049 8919 18107 8925
rect 17126 8888 17132 8900
rect 15226 8860 17132 8888
rect 17126 8848 17132 8860
rect 17184 8848 17190 8900
rect 17313 8891 17371 8897
rect 17313 8857 17325 8891
rect 17359 8888 17371 8891
rect 17586 8888 17592 8900
rect 17359 8860 17592 8888
rect 17359 8857 17371 8860
rect 17313 8851 17371 8857
rect 17586 8848 17592 8860
rect 17644 8848 17650 8900
rect 18616 8832 18644 8928
rect 19242 8916 19248 8968
rect 19300 8916 19306 8968
rect 23842 8956 23848 8968
rect 23690 8928 23848 8956
rect 23842 8916 23848 8928
rect 23900 8916 23906 8968
rect 24210 8916 24216 8968
rect 24268 8916 24274 8968
rect 20441 8891 20499 8897
rect 20441 8857 20453 8891
rect 20487 8888 20499 8891
rect 20714 8888 20720 8900
rect 20487 8860 20720 8888
rect 20487 8857 20499 8860
rect 20441 8851 20499 8857
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 21450 8848 21456 8900
rect 21508 8848 21514 8900
rect 22557 8891 22615 8897
rect 22557 8857 22569 8891
rect 22603 8857 22615 8891
rect 25314 8888 25320 8900
rect 22557 8851 22615 8857
rect 23860 8860 25320 8888
rect 15010 8820 15016 8832
rect 13372 8792 15016 8820
rect 15010 8780 15016 8792
rect 15068 8780 15074 8832
rect 16574 8780 16580 8832
rect 16632 8820 16638 8832
rect 16853 8823 16911 8829
rect 16853 8820 16865 8823
rect 16632 8792 16865 8820
rect 16632 8780 16638 8792
rect 16853 8789 16865 8792
rect 16899 8789 16911 8823
rect 16853 8783 16911 8789
rect 17218 8780 17224 8832
rect 17276 8780 17282 8832
rect 18598 8780 18604 8832
rect 18656 8780 18662 8832
rect 18690 8780 18696 8832
rect 18748 8780 18754 8832
rect 19061 8823 19119 8829
rect 19061 8789 19073 8823
rect 19107 8820 19119 8823
rect 19334 8820 19340 8832
rect 19107 8792 19340 8820
rect 19107 8789 19119 8792
rect 19061 8783 19119 8789
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 21910 8780 21916 8832
rect 21968 8780 21974 8832
rect 22572 8820 22600 8851
rect 23566 8820 23572 8832
rect 22572 8792 23572 8820
rect 23566 8780 23572 8792
rect 23624 8820 23630 8832
rect 23860 8820 23888 8860
rect 25314 8848 25320 8860
rect 25372 8848 25378 8900
rect 23624 8792 23888 8820
rect 24029 8823 24087 8829
rect 23624 8780 23630 8792
rect 24029 8789 24041 8823
rect 24075 8820 24087 8823
rect 24946 8820 24952 8832
rect 24075 8792 24952 8820
rect 24075 8789 24087 8792
rect 24029 8783 24087 8789
rect 24946 8780 24952 8792
rect 25004 8780 25010 8832
rect 1104 8730 26472 8752
rect 1104 8678 7252 8730
rect 7304 8678 7316 8730
rect 7368 8678 7380 8730
rect 7432 8678 7444 8730
rect 7496 8678 7508 8730
rect 7560 8678 13554 8730
rect 13606 8678 13618 8730
rect 13670 8678 13682 8730
rect 13734 8678 13746 8730
rect 13798 8678 13810 8730
rect 13862 8678 19856 8730
rect 19908 8678 19920 8730
rect 19972 8678 19984 8730
rect 20036 8678 20048 8730
rect 20100 8678 20112 8730
rect 20164 8678 26158 8730
rect 26210 8678 26222 8730
rect 26274 8678 26286 8730
rect 26338 8678 26350 8730
rect 26402 8678 26414 8730
rect 26466 8678 26472 8730
rect 1104 8656 26472 8678
rect 1578 8576 1584 8628
rect 1636 8576 1642 8628
rect 2593 8619 2651 8625
rect 2056 8588 2452 8616
rect 1302 8440 1308 8492
rect 1360 8480 1366 8492
rect 2056 8489 2084 8588
rect 2314 8548 2320 8560
rect 2148 8520 2320 8548
rect 2148 8489 2176 8520
rect 2314 8508 2320 8520
rect 2372 8508 2378 8560
rect 2424 8548 2452 8588
rect 2593 8585 2605 8619
rect 2639 8616 2651 8619
rect 2682 8616 2688 8628
rect 2639 8588 2688 8616
rect 2639 8585 2651 8588
rect 2593 8579 2651 8585
rect 2682 8576 2688 8588
rect 2740 8576 2746 8628
rect 3326 8616 3332 8628
rect 3068 8588 3332 8616
rect 2424 8520 2820 8548
rect 2682 8489 2688 8492
rect 1397 8483 1455 8489
rect 1397 8480 1409 8483
rect 1360 8452 1409 8480
rect 1360 8440 1366 8452
rect 1397 8449 1409 8452
rect 1443 8449 1455 8483
rect 1397 8443 1455 8449
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8449 2191 8483
rect 2133 8443 2191 8449
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8449 2467 8483
rect 2681 8480 2688 8489
rect 2643 8452 2688 8480
rect 2409 8443 2467 8449
rect 2681 8443 2688 8452
rect 2317 8415 2375 8421
rect 2317 8381 2329 8415
rect 2363 8381 2375 8415
rect 2424 8412 2452 8443
rect 2682 8440 2688 8443
rect 2740 8440 2746 8492
rect 2792 8480 2820 8520
rect 2866 8480 2872 8492
rect 2792 8452 2872 8480
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3068 8412 3096 8588
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 4062 8576 4068 8628
rect 4120 8576 4126 8628
rect 4246 8576 4252 8628
rect 4304 8576 4310 8628
rect 7561 8619 7619 8625
rect 5920 8588 6776 8616
rect 4080 8548 4108 8576
rect 3160 8520 4108 8548
rect 3160 8489 3188 8520
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 3329 8483 3387 8489
rect 3329 8449 3341 8483
rect 3375 8449 3387 8483
rect 3329 8443 3387 8449
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 3786 8480 3792 8492
rect 3651 8452 3792 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 2424 8384 3096 8412
rect 2317 8375 2375 8381
rect 2130 8304 2136 8356
rect 2188 8304 2194 8356
rect 2222 8304 2228 8356
rect 2280 8304 2286 8356
rect 2332 8344 2360 8375
rect 3142 8344 3148 8356
rect 2332 8316 3148 8344
rect 3142 8304 3148 8316
rect 3200 8304 3206 8356
rect 3344 8344 3372 8443
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 3896 8489 3924 8520
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8449 3939 8483
rect 3881 8443 3939 8449
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8480 4031 8483
rect 4062 8480 4068 8492
rect 4019 8452 4068 8480
rect 4019 8449 4031 8452
rect 3973 8443 4031 8449
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 4154 8440 4160 8492
rect 4212 8440 4218 8492
rect 4264 8489 4292 8576
rect 5920 8557 5948 8588
rect 5905 8551 5963 8557
rect 4724 8520 5120 8548
rect 4724 8492 4752 8520
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8449 4307 8483
rect 4249 8443 4307 8449
rect 4706 8440 4712 8492
rect 4764 8440 4770 8492
rect 4890 8440 4896 8492
rect 4948 8440 4954 8492
rect 5092 8489 5120 8520
rect 5905 8517 5917 8551
rect 5951 8517 5963 8551
rect 5905 8511 5963 8517
rect 5997 8551 6055 8557
rect 5997 8517 6009 8551
rect 6043 8517 6055 8551
rect 6748 8548 6776 8588
rect 7561 8585 7573 8619
rect 7607 8616 7619 8619
rect 7650 8616 7656 8628
rect 7607 8588 7656 8616
rect 7607 8585 7619 8588
rect 7561 8579 7619 8585
rect 7650 8576 7656 8588
rect 7708 8576 7714 8628
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 8205 8619 8263 8625
rect 8205 8616 8217 8619
rect 7800 8588 8217 8616
rect 7800 8576 7806 8588
rect 8205 8585 8217 8588
rect 8251 8585 8263 8619
rect 8205 8579 8263 8585
rect 8386 8576 8392 8628
rect 8444 8616 8450 8628
rect 10873 8619 10931 8625
rect 8444 8588 8610 8616
rect 8444 8576 8450 8588
rect 7837 8551 7895 8557
rect 7837 8548 7849 8551
rect 6748 8520 7512 8548
rect 5997 8511 6055 8517
rect 5810 8489 5816 8492
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8449 5135 8483
rect 5808 8480 5816 8489
rect 5771 8452 5816 8480
rect 5077 8443 5135 8449
rect 5808 8443 5816 8452
rect 5810 8440 5816 8443
rect 5868 8440 5874 8492
rect 3510 8372 3516 8424
rect 3568 8372 3574 8424
rect 3694 8372 3700 8424
rect 3752 8412 3758 8424
rect 4801 8415 4859 8421
rect 3752 8384 4476 8412
rect 3752 8372 3758 8384
rect 4448 8353 4476 8384
rect 4801 8381 4813 8415
rect 4847 8381 4859 8415
rect 4801 8375 4859 8381
rect 4341 8347 4399 8353
rect 4341 8344 4353 8347
rect 3344 8316 4353 8344
rect 4341 8313 4353 8316
rect 4387 8313 4399 8347
rect 4341 8307 4399 8313
rect 4433 8347 4491 8353
rect 4433 8313 4445 8347
rect 4479 8313 4491 8347
rect 4433 8307 4491 8313
rect 2148 8276 2176 8304
rect 2409 8279 2467 8285
rect 2409 8276 2421 8279
rect 2148 8248 2421 8276
rect 2409 8245 2421 8248
rect 2455 8245 2467 8279
rect 2409 8239 2467 8245
rect 2498 8236 2504 8288
rect 2556 8276 2562 8288
rect 2866 8276 2872 8288
rect 2556 8248 2872 8276
rect 2556 8236 2562 8248
rect 2866 8236 2872 8248
rect 2924 8236 2930 8288
rect 3694 8236 3700 8288
rect 3752 8236 3758 8288
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 4522 8276 4528 8288
rect 4120 8248 4528 8276
rect 4120 8236 4126 8248
rect 4522 8236 4528 8248
rect 4580 8276 4586 8288
rect 4816 8276 4844 8375
rect 5626 8372 5632 8424
rect 5684 8412 5690 8424
rect 5905 8415 5963 8421
rect 5905 8412 5917 8415
rect 5684 8384 5917 8412
rect 5684 8372 5690 8384
rect 5905 8381 5917 8384
rect 5951 8381 5963 8415
rect 5905 8375 5963 8381
rect 4890 8304 4896 8356
rect 4948 8304 4954 8356
rect 6012 8344 6040 8511
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8480 6239 8483
rect 6270 8480 6276 8492
rect 6227 8452 6276 8480
rect 6227 8449 6239 8452
rect 6181 8443 6239 8449
rect 6270 8440 6276 8452
rect 6328 8440 6334 8492
rect 6822 8440 6828 8492
rect 6880 8440 6886 8492
rect 6638 8372 6644 8424
rect 6696 8372 6702 8424
rect 7006 8372 7012 8424
rect 7064 8412 7070 8424
rect 7377 8415 7435 8421
rect 7377 8412 7389 8415
rect 7064 8384 7389 8412
rect 7064 8372 7070 8384
rect 7377 8381 7389 8384
rect 7423 8381 7435 8415
rect 7484 8412 7512 8520
rect 7668 8520 7849 8548
rect 7668 8424 7696 8520
rect 7837 8517 7849 8520
rect 7883 8517 7895 8551
rect 7837 8511 7895 8517
rect 7742 8440 7748 8492
rect 7800 8440 7806 8492
rect 7929 8483 7987 8489
rect 7929 8480 7941 8483
rect 7852 8452 7941 8480
rect 7650 8412 7656 8424
rect 7484 8384 7656 8412
rect 7377 8375 7435 8381
rect 7650 8372 7656 8384
rect 7708 8372 7714 8424
rect 6914 8344 6920 8356
rect 6012 8316 6920 8344
rect 6914 8304 6920 8316
rect 6972 8344 6978 8356
rect 7852 8344 7880 8452
rect 7929 8449 7941 8452
rect 7975 8449 7987 8483
rect 7929 8443 7987 8449
rect 8018 8440 8024 8492
rect 8076 8480 8082 8492
rect 8582 8489 8610 8588
rect 10873 8585 10885 8619
rect 10919 8616 10931 8619
rect 11054 8616 11060 8628
rect 10919 8588 11060 8616
rect 10919 8585 10931 8588
rect 10873 8579 10931 8585
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11609 8619 11667 8625
rect 11609 8616 11621 8619
rect 11151 8588 11621 8616
rect 11151 8548 11179 8588
rect 11609 8585 11621 8588
rect 11655 8585 11667 8619
rect 11609 8579 11667 8585
rect 13906 8576 13912 8628
rect 13964 8616 13970 8628
rect 14734 8616 14740 8628
rect 13964 8588 14740 8616
rect 13964 8576 13970 8588
rect 14734 8576 14740 8588
rect 14792 8576 14798 8628
rect 15194 8576 15200 8628
rect 15252 8576 15258 8628
rect 16482 8576 16488 8628
rect 16540 8576 16546 8628
rect 17218 8576 17224 8628
rect 17276 8576 17282 8628
rect 19058 8616 19064 8628
rect 17328 8588 18276 8616
rect 13081 8551 13139 8557
rect 13081 8548 13093 8551
rect 10428 8520 11179 8548
rect 11348 8520 13093 8548
rect 8113 8483 8171 8489
rect 8113 8480 8125 8483
rect 8076 8452 8125 8480
rect 8076 8440 8082 8452
rect 8113 8449 8125 8452
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 8573 8483 8631 8489
rect 8573 8449 8585 8483
rect 8619 8449 8631 8483
rect 8573 8443 8631 8449
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 8481 8415 8539 8421
rect 8481 8381 8493 8415
rect 8527 8412 8539 8415
rect 8772 8412 8800 8440
rect 8527 8384 8800 8412
rect 8527 8381 8539 8384
rect 8481 8375 8539 8381
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 10428 8421 10456 8520
rect 10505 8483 10563 8489
rect 10505 8449 10517 8483
rect 10551 8480 10563 8483
rect 11057 8483 11115 8489
rect 11057 8480 11069 8483
rect 10551 8452 11069 8480
rect 10551 8449 10563 8452
rect 10505 8443 10563 8449
rect 11057 8449 11069 8452
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 10413 8415 10471 8421
rect 10413 8412 10425 8415
rect 9732 8384 10425 8412
rect 9732 8372 9738 8384
rect 10413 8381 10425 8384
rect 10459 8381 10471 8415
rect 10413 8375 10471 8381
rect 6972 8316 7880 8344
rect 6972 8304 6978 8316
rect 4580 8248 4844 8276
rect 4580 8236 4586 8248
rect 6822 8236 6828 8288
rect 6880 8276 6886 8288
rect 8389 8279 8447 8285
rect 8389 8276 8401 8279
rect 6880 8248 8401 8276
rect 6880 8236 6886 8248
rect 8389 8245 8401 8248
rect 8435 8245 8447 8279
rect 10428 8276 10456 8375
rect 11072 8344 11100 8443
rect 11348 8421 11376 8520
rect 13081 8517 13093 8520
rect 13127 8548 13139 8551
rect 15010 8548 15016 8560
rect 13127 8520 13860 8548
rect 14582 8520 15016 8548
rect 13127 8517 13139 8520
rect 13081 8511 13139 8517
rect 13832 8492 13860 8520
rect 15010 8508 15016 8520
rect 15068 8508 15074 8560
rect 11698 8440 11704 8492
rect 11756 8440 11762 8492
rect 12066 8440 12072 8492
rect 12124 8440 12130 8492
rect 12342 8480 12348 8492
rect 12303 8452 12348 8480
rect 12342 8440 12348 8452
rect 12400 8480 12406 8492
rect 12713 8483 12771 8489
rect 12713 8480 12725 8483
rect 12400 8452 12725 8480
rect 12400 8440 12406 8452
rect 12713 8449 12725 8452
rect 12759 8449 12771 8483
rect 12713 8443 12771 8449
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 11333 8415 11391 8421
rect 11333 8381 11345 8415
rect 11379 8381 11391 8415
rect 11333 8375 11391 8381
rect 11440 8384 11744 8412
rect 11440 8344 11468 8384
rect 11072 8316 11468 8344
rect 11716 8344 11744 8384
rect 12912 8344 12940 8443
rect 12986 8440 12992 8492
rect 13044 8440 13050 8492
rect 13170 8440 13176 8492
rect 13228 8440 13234 8492
rect 13814 8440 13820 8492
rect 13872 8440 13878 8492
rect 14185 8483 14243 8489
rect 14185 8480 14197 8483
rect 14016 8452 14197 8480
rect 13004 8412 13032 8440
rect 14016 8412 14044 8452
rect 14185 8449 14197 8452
rect 14231 8449 14243 8483
rect 14185 8443 14243 8449
rect 14921 8483 14979 8489
rect 14921 8449 14933 8483
rect 14967 8480 14979 8483
rect 15212 8480 15240 8576
rect 16301 8551 16359 8557
rect 16301 8517 16313 8551
rect 16347 8548 16359 8551
rect 16500 8548 16528 8576
rect 16347 8520 16528 8548
rect 16347 8517 16359 8520
rect 16301 8511 16359 8517
rect 14967 8452 15240 8480
rect 15841 8483 15899 8489
rect 14967 8449 14979 8452
rect 14921 8443 14979 8449
rect 15841 8449 15853 8483
rect 15887 8480 15899 8483
rect 16117 8483 16175 8489
rect 16117 8480 16129 8483
rect 15887 8452 16129 8480
rect 15887 8449 15899 8452
rect 15841 8443 15899 8449
rect 16117 8449 16129 8452
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 16485 8483 16543 8489
rect 16485 8449 16497 8483
rect 16531 8480 16543 8483
rect 16574 8480 16580 8492
rect 16531 8452 16580 8480
rect 16531 8449 16543 8452
rect 16485 8443 16543 8449
rect 16574 8440 16580 8452
rect 16632 8440 16638 8492
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8480 17003 8483
rect 17236 8480 17264 8576
rect 16991 8452 17264 8480
rect 16991 8449 17003 8452
rect 16945 8443 17003 8449
rect 13004 8384 14044 8412
rect 16022 8372 16028 8424
rect 16080 8372 16086 8424
rect 17126 8372 17132 8424
rect 17184 8412 17190 8424
rect 17328 8412 17356 8588
rect 17586 8508 17592 8560
rect 17644 8548 17650 8560
rect 18141 8551 18199 8557
rect 18141 8548 18153 8551
rect 17644 8520 18153 8548
rect 17644 8508 17650 8520
rect 18141 8517 18153 8520
rect 18187 8517 18199 8551
rect 18248 8548 18276 8588
rect 18708 8588 19064 8616
rect 18708 8548 18736 8588
rect 19058 8576 19064 8588
rect 19116 8616 19122 8628
rect 20717 8619 20775 8625
rect 19116 8588 20392 8616
rect 19116 8576 19122 8588
rect 18248 8520 18814 8548
rect 18141 8511 18199 8517
rect 19702 8508 19708 8560
rect 19760 8548 19766 8560
rect 19981 8551 20039 8557
rect 19981 8548 19993 8551
rect 19760 8520 19993 8548
rect 19760 8508 19766 8520
rect 19981 8517 19993 8520
rect 20027 8517 20039 8551
rect 19981 8511 20039 8517
rect 17405 8483 17463 8489
rect 17405 8449 17417 8483
rect 17451 8480 17463 8483
rect 17451 8452 18368 8480
rect 17451 8449 17463 8452
rect 17405 8443 17463 8449
rect 18340 8424 18368 8452
rect 17184 8384 17356 8412
rect 18233 8415 18291 8421
rect 17184 8372 17190 8384
rect 18233 8381 18245 8415
rect 18279 8381 18291 8415
rect 18233 8375 18291 8381
rect 11716 8316 14596 8344
rect 14568 8288 14596 8316
rect 14734 8304 14740 8356
rect 14792 8344 14798 8356
rect 15657 8347 15715 8353
rect 15657 8344 15669 8347
rect 14792 8316 15669 8344
rect 14792 8304 14798 8316
rect 15657 8313 15669 8316
rect 15703 8313 15715 8347
rect 18248 8344 18276 8375
rect 18322 8372 18328 8424
rect 18380 8412 18386 8424
rect 19242 8412 19248 8424
rect 18380 8384 19248 8412
rect 18380 8372 18386 8384
rect 19242 8372 19248 8384
rect 19300 8412 19306 8424
rect 20257 8415 20315 8421
rect 20257 8412 20269 8415
rect 19300 8384 20269 8412
rect 19300 8372 19306 8384
rect 20257 8381 20269 8384
rect 20303 8381 20315 8415
rect 20257 8375 20315 8381
rect 18598 8344 18604 8356
rect 18248 8316 18604 8344
rect 15657 8307 15715 8313
rect 18598 8304 18604 8316
rect 18656 8304 18662 8356
rect 20364 8344 20392 8588
rect 20717 8585 20729 8619
rect 20763 8616 20775 8619
rect 20806 8616 20812 8628
rect 20763 8588 20812 8616
rect 20763 8585 20775 8588
rect 20717 8579 20775 8585
rect 20806 8576 20812 8588
rect 20864 8576 20870 8628
rect 21082 8576 21088 8628
rect 21140 8576 21146 8628
rect 21818 8576 21824 8628
rect 21876 8576 21882 8628
rect 21910 8576 21916 8628
rect 21968 8616 21974 8628
rect 23753 8619 23811 8625
rect 21968 8588 22094 8616
rect 21968 8576 21974 8588
rect 20901 8483 20959 8489
rect 20901 8449 20913 8483
rect 20947 8480 20959 8483
rect 21100 8480 21128 8576
rect 21177 8551 21235 8557
rect 21177 8517 21189 8551
rect 21223 8548 21235 8551
rect 21266 8548 21272 8560
rect 21223 8520 21272 8548
rect 21223 8517 21235 8520
rect 21177 8511 21235 8517
rect 21266 8508 21272 8520
rect 21324 8508 21330 8560
rect 20947 8452 21128 8480
rect 20947 8449 20959 8452
rect 20901 8443 20959 8449
rect 21085 8415 21143 8421
rect 21085 8381 21097 8415
rect 21131 8412 21143 8415
rect 22066 8412 22094 8588
rect 23753 8585 23765 8619
rect 23799 8616 23811 8619
rect 23934 8616 23940 8628
rect 23799 8588 23940 8616
rect 23799 8585 23811 8588
rect 23753 8579 23811 8585
rect 23934 8576 23940 8588
rect 23992 8576 23998 8628
rect 25593 8619 25651 8625
rect 25593 8585 25605 8619
rect 25639 8616 25651 8619
rect 25682 8616 25688 8628
rect 25639 8588 25688 8616
rect 25639 8585 25651 8588
rect 25593 8579 25651 8585
rect 25682 8576 25688 8588
rect 25740 8576 25746 8628
rect 24210 8548 24216 8560
rect 23860 8520 24216 8548
rect 23658 8440 23664 8492
rect 23716 8480 23722 8492
rect 23860 8489 23888 8520
rect 24210 8508 24216 8520
rect 24268 8508 24274 8560
rect 23845 8483 23903 8489
rect 23845 8480 23857 8483
rect 23716 8452 23857 8480
rect 23716 8440 23722 8452
rect 23845 8449 23857 8452
rect 23891 8449 23903 8483
rect 23845 8443 23903 8449
rect 22373 8415 22431 8421
rect 22373 8412 22385 8415
rect 21131 8384 22385 8412
rect 21131 8381 21143 8384
rect 21085 8375 21143 8381
rect 22373 8381 22385 8384
rect 22419 8381 22431 8415
rect 22373 8375 22431 8381
rect 23201 8415 23259 8421
rect 23201 8381 23213 8415
rect 23247 8412 23259 8415
rect 23382 8412 23388 8424
rect 23247 8384 23388 8412
rect 23247 8381 23259 8384
rect 23201 8375 23259 8381
rect 23382 8372 23388 8384
rect 23440 8372 23446 8424
rect 24121 8415 24179 8421
rect 24121 8381 24133 8415
rect 24167 8412 24179 8415
rect 25130 8412 25136 8424
rect 24167 8384 25136 8412
rect 24167 8381 24179 8384
rect 24121 8375 24179 8381
rect 25130 8372 25136 8384
rect 25188 8372 25194 8424
rect 20364 8316 23980 8344
rect 11149 8279 11207 8285
rect 11149 8276 11161 8279
rect 10428 8248 11161 8276
rect 8389 8239 8447 8245
rect 11149 8245 11161 8248
rect 11195 8245 11207 8279
rect 11149 8239 11207 8245
rect 11238 8236 11244 8288
rect 11296 8236 11302 8288
rect 13262 8236 13268 8288
rect 13320 8236 13326 8288
rect 14550 8236 14556 8288
rect 14608 8236 14614 8288
rect 17129 8279 17187 8285
rect 17129 8245 17141 8279
rect 17175 8276 17187 8279
rect 17218 8276 17224 8288
rect 17175 8248 17224 8276
rect 17175 8245 17187 8248
rect 17129 8239 17187 8245
rect 17218 8236 17224 8248
rect 17276 8236 17282 8288
rect 21174 8236 21180 8288
rect 21232 8236 21238 8288
rect 23952 8276 23980 8316
rect 25240 8288 25268 8466
rect 25222 8276 25228 8288
rect 23952 8248 25228 8276
rect 25222 8236 25228 8248
rect 25280 8236 25286 8288
rect 1104 8186 26312 8208
rect 1104 8134 4101 8186
rect 4153 8134 4165 8186
rect 4217 8134 4229 8186
rect 4281 8134 4293 8186
rect 4345 8134 4357 8186
rect 4409 8134 10403 8186
rect 10455 8134 10467 8186
rect 10519 8134 10531 8186
rect 10583 8134 10595 8186
rect 10647 8134 10659 8186
rect 10711 8134 16705 8186
rect 16757 8134 16769 8186
rect 16821 8134 16833 8186
rect 16885 8134 16897 8186
rect 16949 8134 16961 8186
rect 17013 8134 23007 8186
rect 23059 8134 23071 8186
rect 23123 8134 23135 8186
rect 23187 8134 23199 8186
rect 23251 8134 23263 8186
rect 23315 8134 26312 8186
rect 1104 8112 26312 8134
rect 2866 8032 2872 8084
rect 2924 8032 2930 8084
rect 3142 8032 3148 8084
rect 3200 8072 3206 8084
rect 3786 8072 3792 8084
rect 3200 8044 3792 8072
rect 3200 8032 3206 8044
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 5534 8032 5540 8084
rect 5592 8032 5598 8084
rect 7098 8032 7104 8084
rect 7156 8072 7162 8084
rect 7469 8075 7527 8081
rect 7469 8072 7481 8075
rect 7156 8044 7481 8072
rect 7156 8032 7162 8044
rect 7469 8041 7481 8044
rect 7515 8041 7527 8075
rect 7469 8035 7527 8041
rect 10870 8032 10876 8084
rect 10928 8032 10934 8084
rect 11238 8032 11244 8084
rect 11296 8032 11302 8084
rect 22465 8075 22523 8081
rect 22465 8041 22477 8075
rect 22511 8072 22523 8075
rect 22554 8072 22560 8084
rect 22511 8044 22560 8072
rect 22511 8041 22523 8044
rect 22465 8035 22523 8041
rect 22554 8032 22560 8044
rect 22612 8032 22618 8084
rect 3804 7936 3832 8032
rect 7650 7964 7656 8016
rect 7708 7964 7714 8016
rect 7742 7964 7748 8016
rect 7800 8004 7806 8016
rect 7929 8007 7987 8013
rect 7929 8004 7941 8007
rect 7800 7976 7941 8004
rect 7800 7964 7806 7976
rect 7929 7973 7941 7976
rect 7975 7973 7987 8007
rect 7929 7967 7987 7973
rect 4985 7939 5043 7945
rect 3804 7908 4016 7936
rect 2869 7871 2927 7877
rect 2869 7837 2881 7871
rect 2915 7868 2927 7871
rect 2958 7868 2964 7880
rect 2915 7840 2964 7868
rect 2915 7837 2927 7840
rect 2869 7831 2927 7837
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3326 7868 3332 7880
rect 3099 7840 3332 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3326 7828 3332 7840
rect 3384 7828 3390 7880
rect 3694 7828 3700 7880
rect 3752 7868 3758 7880
rect 3988 7877 4016 7908
rect 4985 7905 4997 7939
rect 5031 7936 5043 7939
rect 11256 7936 11284 8032
rect 13262 8004 13268 8016
rect 12406 7976 13268 8004
rect 5031 7908 6132 7936
rect 5031 7905 5043 7908
rect 4985 7899 5043 7905
rect 6104 7880 6132 7908
rect 7392 7908 8800 7936
rect 3789 7871 3847 7877
rect 3789 7868 3801 7871
rect 3752 7840 3801 7868
rect 3752 7828 3758 7840
rect 3789 7837 3801 7840
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7868 5227 7871
rect 5810 7868 5816 7880
rect 5215 7840 5816 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 5810 7828 5816 7840
rect 5868 7868 5874 7880
rect 5868 7840 6040 7868
rect 5868 7828 5874 7840
rect 5077 7803 5135 7809
rect 5077 7769 5089 7803
rect 5123 7800 5135 7803
rect 5902 7800 5908 7812
rect 5123 7772 5908 7800
rect 5123 7769 5135 7772
rect 5077 7763 5135 7769
rect 5902 7760 5908 7772
rect 5960 7760 5966 7812
rect 6012 7800 6040 7840
rect 6086 7828 6092 7880
rect 6144 7828 6150 7880
rect 6362 7828 6368 7880
rect 6420 7828 6426 7880
rect 6454 7828 6460 7880
rect 6512 7828 6518 7880
rect 6546 7828 6552 7880
rect 6604 7868 6610 7880
rect 7392 7877 7420 7908
rect 8772 7880 8800 7908
rect 11072 7908 11284 7936
rect 11333 7939 11391 7945
rect 6825 7871 6883 7877
rect 6825 7868 6837 7871
rect 6604 7840 6837 7868
rect 6604 7828 6610 7840
rect 6825 7837 6837 7840
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7837 7435 7871
rect 7377 7831 7435 7837
rect 7561 7871 7619 7877
rect 7561 7837 7573 7871
rect 7607 7837 7619 7871
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 7561 7831 7619 7837
rect 7668 7840 7941 7868
rect 6380 7800 6408 7828
rect 6012 7772 6408 7800
rect 6840 7800 6868 7831
rect 7576 7800 7604 7831
rect 6840 7772 7604 7800
rect 3970 7692 3976 7744
rect 4028 7692 4034 7744
rect 6270 7692 6276 7744
rect 6328 7732 6334 7744
rect 7668 7732 7696 7840
rect 7929 7837 7941 7840
rect 7975 7868 7987 7871
rect 8018 7868 8024 7880
rect 7975 7840 8024 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 8128 7800 8156 7831
rect 8754 7828 8760 7880
rect 8812 7828 8818 7880
rect 11072 7877 11100 7908
rect 11333 7905 11345 7939
rect 11379 7936 11391 7939
rect 12406 7936 12434 7976
rect 13262 7964 13268 7976
rect 13320 7964 13326 8016
rect 13814 7964 13820 8016
rect 13872 8004 13878 8016
rect 14093 8007 14151 8013
rect 14093 8004 14105 8007
rect 13872 7976 14105 8004
rect 13872 7964 13878 7976
rect 14093 7973 14105 7976
rect 14139 7973 14151 8007
rect 14093 7967 14151 7973
rect 11379 7908 12434 7936
rect 11379 7905 11391 7908
rect 11333 7899 11391 7905
rect 12526 7896 12532 7948
rect 12584 7936 12590 7948
rect 12621 7939 12679 7945
rect 12621 7936 12633 7939
rect 12584 7908 12633 7936
rect 12584 7896 12590 7908
rect 12621 7905 12633 7908
rect 12667 7905 12679 7939
rect 12621 7899 12679 7905
rect 12894 7896 12900 7948
rect 12952 7896 12958 7948
rect 13906 7896 13912 7948
rect 13964 7936 13970 7948
rect 14369 7939 14427 7945
rect 14369 7936 14381 7939
rect 13964 7908 14381 7936
rect 13964 7896 13970 7908
rect 14369 7905 14381 7908
rect 14415 7905 14427 7939
rect 14369 7899 14427 7905
rect 14550 7896 14556 7948
rect 14608 7936 14614 7948
rect 15289 7939 15347 7945
rect 15289 7936 15301 7939
rect 14608 7908 15301 7936
rect 14608 7896 14614 7908
rect 15289 7905 15301 7908
rect 15335 7905 15347 7939
rect 16577 7939 16635 7945
rect 16577 7936 16589 7939
rect 15289 7899 15347 7905
rect 16040 7908 16589 7936
rect 16040 7880 16068 7908
rect 16577 7905 16589 7908
rect 16623 7905 16635 7939
rect 16577 7899 16635 7905
rect 17034 7896 17040 7948
rect 17092 7896 17098 7948
rect 18506 7896 18512 7948
rect 18564 7936 18570 7948
rect 19889 7939 19947 7945
rect 19889 7936 19901 7939
rect 18564 7908 19901 7936
rect 18564 7896 18570 7908
rect 19889 7905 19901 7908
rect 19935 7905 19947 7939
rect 19889 7899 19947 7905
rect 21634 7896 21640 7948
rect 21692 7896 21698 7948
rect 21913 7939 21971 7945
rect 21913 7905 21925 7939
rect 21959 7936 21971 7939
rect 23658 7936 23664 7948
rect 21959 7908 23664 7936
rect 21959 7905 21971 7908
rect 21913 7899 21971 7905
rect 23658 7896 23664 7908
rect 23716 7896 23722 7948
rect 24946 7896 24952 7948
rect 25004 7896 25010 7948
rect 25314 7896 25320 7948
rect 25372 7936 25378 7948
rect 25685 7939 25743 7945
rect 25685 7936 25697 7939
rect 25372 7908 25697 7936
rect 25372 7896 25378 7908
rect 25685 7905 25697 7908
rect 25731 7905 25743 7939
rect 25685 7899 25743 7905
rect 25958 7896 25964 7948
rect 26016 7896 26022 7948
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7837 11115 7871
rect 11057 7831 11115 7837
rect 11241 7871 11299 7877
rect 11241 7837 11253 7871
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7868 11483 7871
rect 12066 7868 12072 7880
rect 11471 7840 12072 7868
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 8036 7772 8156 7800
rect 11256 7800 11284 7831
rect 12066 7828 12072 7840
rect 12124 7828 12130 7880
rect 12253 7871 12311 7877
rect 12253 7837 12265 7871
rect 12299 7837 12311 7871
rect 12253 7831 12311 7837
rect 12437 7871 12495 7877
rect 12437 7837 12449 7871
rect 12483 7868 12495 7871
rect 12710 7868 12716 7880
rect 12483 7840 12716 7868
rect 12483 7837 12495 7840
rect 12437 7831 12495 7837
rect 11790 7800 11796 7812
rect 11256 7772 11796 7800
rect 8036 7744 8064 7772
rect 11790 7760 11796 7772
rect 11848 7760 11854 7812
rect 12268 7800 12296 7831
rect 12710 7828 12716 7840
rect 12768 7828 12774 7880
rect 12986 7828 12992 7880
rect 13044 7868 13050 7880
rect 13262 7868 13268 7880
rect 13044 7840 13268 7868
rect 13044 7828 13050 7840
rect 13262 7828 13268 7840
rect 13320 7828 13326 7880
rect 14458 7828 14464 7880
rect 14516 7828 14522 7880
rect 15654 7828 15660 7880
rect 15712 7828 15718 7880
rect 16022 7828 16028 7880
rect 16080 7828 16086 7880
rect 16482 7828 16488 7880
rect 16540 7828 16546 7880
rect 16669 7871 16727 7877
rect 16669 7837 16681 7871
rect 16715 7837 16727 7871
rect 16669 7831 16727 7837
rect 12268 7772 12434 7800
rect 6328 7704 7696 7732
rect 6328 7692 6334 7704
rect 8018 7692 8024 7744
rect 8076 7692 8082 7744
rect 12406 7732 12434 7772
rect 16574 7760 16580 7812
rect 16632 7800 16638 7812
rect 16684 7800 16712 7831
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 19429 7871 19487 7877
rect 19429 7868 19441 7871
rect 19392 7840 19441 7868
rect 19392 7828 19398 7840
rect 19429 7837 19441 7840
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 22186 7828 22192 7880
rect 22244 7868 22250 7880
rect 22281 7871 22339 7877
rect 22281 7868 22293 7871
rect 22244 7840 22293 7868
rect 22244 7828 22250 7840
rect 22281 7837 22293 7840
rect 22327 7837 22339 7871
rect 22281 7831 22339 7837
rect 22373 7871 22431 7877
rect 22373 7837 22385 7871
rect 22419 7837 22431 7871
rect 22373 7831 22431 7837
rect 16632 7772 16712 7800
rect 16632 7760 16638 7772
rect 13998 7732 14004 7744
rect 12406 7704 14004 7732
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 16684 7732 16712 7772
rect 17218 7760 17224 7812
rect 17276 7800 17282 7812
rect 17313 7803 17371 7809
rect 17313 7800 17325 7803
rect 17276 7772 17325 7800
rect 17276 7760 17282 7772
rect 17313 7769 17325 7772
rect 17359 7769 17371 7803
rect 17313 7763 17371 7769
rect 17586 7760 17592 7812
rect 17644 7800 17650 7812
rect 19061 7803 19119 7809
rect 17644 7772 17802 7800
rect 17644 7760 17650 7772
rect 19061 7769 19073 7803
rect 19107 7769 19119 7803
rect 22005 7803 22063 7809
rect 22005 7800 22017 7803
rect 21206 7772 21312 7800
rect 19061 7763 19119 7769
rect 18046 7732 18052 7744
rect 16684 7704 18052 7732
rect 18046 7692 18052 7704
rect 18104 7732 18110 7744
rect 19076 7732 19104 7763
rect 21284 7744 21312 7772
rect 21928 7772 22017 7800
rect 21928 7744 21956 7772
rect 22005 7769 22017 7772
rect 22051 7769 22063 7803
rect 22388 7800 22416 7831
rect 22005 7763 22063 7769
rect 22296 7772 22416 7800
rect 22296 7744 22324 7772
rect 18104 7704 19104 7732
rect 18104 7692 18110 7704
rect 19242 7692 19248 7744
rect 19300 7692 19306 7744
rect 21266 7692 21272 7744
rect 21324 7732 21330 7744
rect 21450 7732 21456 7744
rect 21324 7704 21456 7732
rect 21324 7692 21330 7704
rect 21450 7692 21456 7704
rect 21508 7692 21514 7744
rect 21910 7692 21916 7744
rect 21968 7692 21974 7744
rect 22094 7692 22100 7744
rect 22152 7692 22158 7744
rect 22278 7692 22284 7744
rect 22336 7692 22342 7744
rect 24118 7692 24124 7744
rect 24176 7732 24182 7744
rect 24397 7735 24455 7741
rect 24397 7732 24409 7735
rect 24176 7704 24409 7732
rect 24176 7692 24182 7704
rect 24397 7701 24409 7704
rect 24443 7701 24455 7735
rect 24397 7695 24455 7701
rect 1104 7642 26472 7664
rect 1104 7590 7252 7642
rect 7304 7590 7316 7642
rect 7368 7590 7380 7642
rect 7432 7590 7444 7642
rect 7496 7590 7508 7642
rect 7560 7590 13554 7642
rect 13606 7590 13618 7642
rect 13670 7590 13682 7642
rect 13734 7590 13746 7642
rect 13798 7590 13810 7642
rect 13862 7590 19856 7642
rect 19908 7590 19920 7642
rect 19972 7590 19984 7642
rect 20036 7590 20048 7642
rect 20100 7590 20112 7642
rect 20164 7590 26158 7642
rect 26210 7590 26222 7642
rect 26274 7590 26286 7642
rect 26338 7590 26350 7642
rect 26402 7590 26414 7642
rect 26466 7590 26472 7642
rect 1104 7568 26472 7590
rect 6914 7488 6920 7540
rect 6972 7528 6978 7540
rect 7009 7531 7067 7537
rect 7009 7528 7021 7531
rect 6972 7500 7021 7528
rect 6972 7488 6978 7500
rect 7009 7497 7021 7500
rect 7055 7497 7067 7531
rect 7009 7491 7067 7497
rect 7926 7488 7932 7540
rect 7984 7528 7990 7540
rect 8757 7531 8815 7537
rect 8757 7528 8769 7531
rect 7984 7500 8769 7528
rect 7984 7488 7990 7500
rect 8757 7497 8769 7500
rect 8803 7497 8815 7531
rect 8757 7491 8815 7497
rect 11606 7488 11612 7540
rect 11664 7528 11670 7540
rect 11701 7531 11759 7537
rect 11701 7528 11713 7531
rect 11664 7500 11713 7528
rect 11664 7488 11670 7500
rect 11701 7497 11713 7500
rect 11747 7497 11759 7531
rect 11701 7491 11759 7497
rect 14458 7488 14464 7540
rect 14516 7528 14522 7540
rect 15102 7528 15108 7540
rect 14516 7500 15108 7528
rect 14516 7488 14522 7500
rect 15102 7488 15108 7500
rect 15160 7528 15166 7540
rect 15473 7531 15531 7537
rect 15473 7528 15485 7531
rect 15160 7500 15485 7528
rect 15160 7488 15166 7500
rect 15473 7497 15485 7500
rect 15519 7497 15531 7531
rect 15473 7491 15531 7497
rect 16482 7488 16488 7540
rect 16540 7528 16546 7540
rect 17497 7531 17555 7537
rect 17497 7528 17509 7531
rect 16540 7500 17509 7528
rect 16540 7488 16546 7500
rect 17497 7497 17509 7500
rect 17543 7528 17555 7531
rect 18690 7528 18696 7540
rect 17543 7500 18696 7528
rect 17543 7497 17555 7500
rect 17497 7491 17555 7497
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 19242 7528 19248 7540
rect 18984 7500 19248 7528
rect 6638 7420 6644 7472
rect 6696 7460 6702 7472
rect 7193 7463 7251 7469
rect 7193 7460 7205 7463
rect 6696 7432 7205 7460
rect 6696 7420 6702 7432
rect 7193 7429 7205 7432
rect 7239 7460 7251 7463
rect 8018 7460 8024 7472
rect 7239 7432 8024 7460
rect 7239 7429 7251 7432
rect 7193 7423 7251 7429
rect 8018 7420 8024 7432
rect 8076 7420 8082 7472
rect 9401 7463 9459 7469
rect 9401 7460 9413 7463
rect 8864 7432 9413 7460
rect 6086 7352 6092 7404
rect 6144 7352 6150 7404
rect 6362 7352 6368 7404
rect 6420 7392 6426 7404
rect 6420 7364 6776 7392
rect 6420 7352 6426 7364
rect 6104 7324 6132 7352
rect 6457 7327 6515 7333
rect 6457 7324 6469 7327
rect 6104 7296 6469 7324
rect 6457 7293 6469 7296
rect 6503 7293 6515 7327
rect 6457 7287 6515 7293
rect 6546 7284 6552 7336
rect 6604 7324 6610 7336
rect 6641 7327 6699 7333
rect 6641 7324 6653 7327
rect 6604 7296 6653 7324
rect 6604 7284 6610 7296
rect 6641 7293 6653 7296
rect 6687 7293 6699 7327
rect 6748 7324 6776 7364
rect 6822 7352 6828 7404
rect 6880 7392 6886 7404
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 6880 7364 7389 7392
rect 6880 7352 6886 7364
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 7742 7352 7748 7404
rect 7800 7352 7806 7404
rect 8662 7352 8668 7404
rect 8720 7352 8726 7404
rect 8864 7401 8892 7432
rect 9401 7429 9413 7432
rect 9447 7429 9459 7463
rect 13081 7463 13139 7469
rect 13081 7460 13093 7463
rect 9401 7423 9459 7429
rect 11716 7432 13093 7460
rect 11716 7404 11744 7432
rect 13081 7429 13093 7432
rect 13127 7460 13139 7463
rect 13170 7460 13176 7472
rect 13127 7432 13176 7460
rect 13127 7429 13139 7432
rect 13081 7423 13139 7429
rect 13170 7420 13176 7432
rect 13228 7420 13234 7472
rect 14752 7432 15884 7460
rect 8849 7395 8907 7401
rect 8849 7361 8861 7395
rect 8895 7361 8907 7395
rect 8849 7355 8907 7361
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7361 9367 7395
rect 9309 7355 9367 7361
rect 9493 7395 9551 7401
rect 9493 7361 9505 7395
rect 9539 7392 9551 7395
rect 9582 7392 9588 7404
rect 9539 7364 9588 7392
rect 9539 7361 9551 7364
rect 9493 7355 9551 7361
rect 7760 7324 7788 7352
rect 6748 7296 7788 7324
rect 9324 7324 9352 7355
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 11698 7352 11704 7404
rect 11756 7352 11762 7404
rect 11790 7352 11796 7404
rect 11848 7392 11854 7404
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11848 7364 11897 7392
rect 11848 7352 11854 7364
rect 11885 7361 11897 7364
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 12161 7395 12219 7401
rect 12161 7361 12173 7395
rect 12207 7392 12219 7395
rect 12434 7392 12440 7404
rect 12207 7364 12440 7392
rect 12207 7361 12219 7364
rect 12161 7355 12219 7361
rect 12434 7352 12440 7364
rect 12492 7352 12498 7404
rect 12621 7395 12679 7401
rect 12621 7361 12633 7395
rect 12667 7392 12679 7395
rect 12986 7392 12992 7404
rect 12667 7364 12992 7392
rect 12667 7361 12679 7364
rect 12621 7355 12679 7361
rect 12986 7352 12992 7364
rect 13044 7352 13050 7404
rect 13449 7395 13507 7401
rect 13449 7361 13461 7395
rect 13495 7392 13507 7395
rect 13998 7392 14004 7404
rect 13495 7364 14004 7392
rect 13495 7361 13507 7364
rect 13449 7355 13507 7361
rect 13998 7352 14004 7364
rect 14056 7392 14062 7404
rect 14366 7392 14372 7404
rect 14056 7364 14372 7392
rect 14056 7352 14062 7364
rect 14366 7352 14372 7364
rect 14424 7352 14430 7404
rect 14752 7401 14780 7432
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7361 14795 7395
rect 14737 7355 14795 7361
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7361 15163 7395
rect 15105 7355 15163 7361
rect 9398 7324 9404 7336
rect 9324 7296 9404 7324
rect 6641 7287 6699 7293
rect 9398 7284 9404 7296
rect 9456 7324 9462 7336
rect 12526 7324 12532 7336
rect 9456 7296 12532 7324
rect 9456 7284 9462 7296
rect 12526 7284 12532 7296
rect 12584 7324 12590 7336
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 12584 7296 14657 7324
rect 12584 7284 12590 7296
rect 14645 7293 14657 7296
rect 14691 7293 14703 7327
rect 15120 7324 15148 7355
rect 15654 7352 15660 7404
rect 15712 7352 15718 7404
rect 15856 7401 15884 7432
rect 15841 7395 15899 7401
rect 15841 7361 15853 7395
rect 15887 7392 15899 7395
rect 16500 7392 16528 7488
rect 17586 7460 17592 7472
rect 17236 7432 17592 7460
rect 17236 7404 17264 7432
rect 17586 7420 17592 7432
rect 17644 7460 17650 7472
rect 18984 7469 19012 7500
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 20714 7488 20720 7540
rect 20772 7488 20778 7540
rect 21085 7531 21143 7537
rect 21085 7497 21097 7531
rect 21131 7528 21143 7531
rect 21818 7528 21824 7540
rect 21131 7500 21824 7528
rect 21131 7497 21143 7500
rect 21085 7491 21143 7497
rect 21818 7488 21824 7500
rect 21876 7488 21882 7540
rect 24118 7528 24124 7540
rect 23952 7500 24124 7528
rect 18969 7463 19027 7469
rect 17644 7432 17802 7460
rect 17644 7420 17650 7432
rect 18969 7429 18981 7463
rect 19015 7429 19027 7463
rect 18969 7423 19027 7429
rect 21358 7420 21364 7472
rect 21416 7460 21422 7472
rect 21726 7460 21732 7472
rect 21416 7432 21732 7460
rect 21416 7420 21422 7432
rect 21726 7420 21732 7432
rect 21784 7420 21790 7472
rect 23014 7420 23020 7472
rect 23072 7460 23078 7472
rect 23952 7469 23980 7500
rect 24118 7488 24124 7500
rect 24176 7488 24182 7540
rect 25406 7488 25412 7540
rect 25464 7488 25470 7540
rect 23293 7463 23351 7469
rect 23293 7460 23305 7463
rect 23072 7432 23305 7460
rect 23072 7420 23078 7432
rect 23293 7429 23305 7432
rect 23339 7429 23351 7463
rect 23293 7423 23351 7429
rect 23937 7463 23995 7469
rect 23937 7429 23949 7463
rect 23983 7429 23995 7463
rect 25222 7460 25228 7472
rect 25162 7432 25228 7460
rect 23937 7423 23995 7429
rect 25222 7420 25228 7432
rect 25280 7420 25286 7472
rect 15887 7364 16528 7392
rect 15887 7361 15899 7364
rect 15841 7355 15899 7361
rect 17218 7352 17224 7404
rect 17276 7352 17282 7404
rect 17310 7352 17316 7404
rect 17368 7352 17374 7404
rect 20901 7395 20959 7401
rect 20901 7361 20913 7395
rect 20947 7361 20959 7395
rect 20901 7355 20959 7361
rect 21177 7395 21235 7401
rect 21177 7361 21189 7395
rect 21223 7392 21235 7395
rect 21376 7392 21404 7420
rect 21223 7364 21404 7392
rect 21223 7361 21235 7364
rect 21177 7355 21235 7361
rect 15749 7327 15807 7333
rect 15749 7324 15761 7327
rect 15120 7296 15761 7324
rect 14645 7287 14703 7293
rect 15749 7293 15761 7296
rect 15795 7293 15807 7327
rect 15749 7287 15807 7293
rect 15933 7327 15991 7333
rect 15933 7293 15945 7327
rect 15979 7324 15991 7327
rect 16574 7324 16580 7336
rect 15979 7296 16580 7324
rect 15979 7293 15991 7296
rect 15933 7287 15991 7293
rect 15764 7256 15792 7287
rect 16574 7284 16580 7296
rect 16632 7284 16638 7336
rect 19245 7327 19303 7333
rect 19245 7293 19257 7327
rect 19291 7293 19303 7327
rect 20916 7324 20944 7355
rect 21634 7352 21640 7404
rect 21692 7352 21698 7404
rect 21652 7324 21680 7352
rect 20916 7296 21680 7324
rect 19245 7287 19303 7293
rect 16482 7256 16488 7268
rect 15764 7228 16488 7256
rect 16482 7216 16488 7228
rect 16540 7216 16546 7268
rect 11882 7148 11888 7200
rect 11940 7188 11946 7200
rect 11977 7191 12035 7197
rect 11977 7188 11989 7191
rect 11940 7160 11989 7188
rect 11940 7148 11946 7160
rect 11977 7157 11989 7160
rect 12023 7157 12035 7191
rect 11977 7151 12035 7157
rect 13909 7191 13967 7197
rect 13909 7157 13921 7191
rect 13955 7188 13967 7191
rect 13998 7188 14004 7200
rect 13955 7160 14004 7188
rect 13955 7157 13967 7160
rect 13909 7151 13967 7157
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 15010 7148 15016 7200
rect 15068 7148 15074 7200
rect 15286 7148 15292 7200
rect 15344 7148 15350 7200
rect 16669 7191 16727 7197
rect 16669 7157 16681 7191
rect 16715 7188 16727 7191
rect 17126 7188 17132 7200
rect 16715 7160 17132 7188
rect 16715 7157 16727 7160
rect 16669 7151 16727 7157
rect 17126 7148 17132 7160
rect 17184 7148 17190 7200
rect 18322 7148 18328 7200
rect 18380 7188 18386 7200
rect 19260 7188 19288 7287
rect 22002 7284 22008 7336
rect 22060 7324 22066 7336
rect 22204 7324 22232 7378
rect 22060 7296 22232 7324
rect 23569 7327 23627 7333
rect 22060 7284 22066 7296
rect 23569 7293 23581 7327
rect 23615 7324 23627 7327
rect 23658 7324 23664 7336
rect 23615 7296 23664 7324
rect 23615 7293 23627 7296
rect 23569 7287 23627 7293
rect 23658 7284 23664 7296
rect 23716 7284 23722 7336
rect 18380 7160 19288 7188
rect 21821 7191 21879 7197
rect 18380 7148 18386 7160
rect 21821 7157 21833 7191
rect 21867 7188 21879 7191
rect 22278 7188 22284 7200
rect 21867 7160 22284 7188
rect 21867 7157 21879 7160
rect 21821 7151 21879 7157
rect 22278 7148 22284 7160
rect 22336 7148 22342 7200
rect 1104 7098 26312 7120
rect 1104 7046 4101 7098
rect 4153 7046 4165 7098
rect 4217 7046 4229 7098
rect 4281 7046 4293 7098
rect 4345 7046 4357 7098
rect 4409 7046 10403 7098
rect 10455 7046 10467 7098
rect 10519 7046 10531 7098
rect 10583 7046 10595 7098
rect 10647 7046 10659 7098
rect 10711 7046 16705 7098
rect 16757 7046 16769 7098
rect 16821 7046 16833 7098
rect 16885 7046 16897 7098
rect 16949 7046 16961 7098
rect 17013 7046 23007 7098
rect 23059 7046 23071 7098
rect 23123 7046 23135 7098
rect 23187 7046 23199 7098
rect 23251 7046 23263 7098
rect 23315 7046 26312 7098
rect 1104 7024 26312 7046
rect 5902 6944 5908 6996
rect 5960 6944 5966 6996
rect 6638 6944 6644 6996
rect 6696 6984 6702 6996
rect 7009 6987 7067 6993
rect 7009 6984 7021 6987
rect 6696 6956 7021 6984
rect 6696 6944 6702 6956
rect 7009 6953 7021 6956
rect 7055 6953 7067 6987
rect 7009 6947 7067 6953
rect 11136 6987 11194 6993
rect 11136 6953 11148 6987
rect 11182 6984 11194 6987
rect 11882 6984 11888 6996
rect 11182 6956 11888 6984
rect 11182 6953 11194 6956
rect 11136 6947 11194 6953
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 12710 6944 12716 6996
rect 12768 6984 12774 6996
rect 13081 6987 13139 6993
rect 13081 6984 13093 6987
rect 12768 6956 13093 6984
rect 12768 6944 12774 6956
rect 13081 6953 13093 6956
rect 13127 6953 13139 6987
rect 13081 6947 13139 6953
rect 13817 6987 13875 6993
rect 13817 6953 13829 6987
rect 13863 6984 13875 6987
rect 13906 6984 13912 6996
rect 13863 6956 13912 6984
rect 13863 6953 13875 6956
rect 13817 6947 13875 6953
rect 13906 6944 13912 6956
rect 13964 6944 13970 6996
rect 21545 6987 21603 6993
rect 21545 6953 21557 6987
rect 21591 6953 21603 6987
rect 21545 6947 21603 6953
rect 2593 6851 2651 6857
rect 2593 6817 2605 6851
rect 2639 6848 2651 6851
rect 3050 6848 3056 6860
rect 2639 6820 3056 6848
rect 2639 6817 2651 6820
rect 2593 6811 2651 6817
rect 3050 6808 3056 6820
rect 3108 6808 3114 6860
rect 6365 6851 6423 6857
rect 6365 6817 6377 6851
rect 6411 6848 6423 6851
rect 6656 6848 6684 6944
rect 12621 6919 12679 6925
rect 12621 6885 12633 6919
rect 12667 6916 12679 6919
rect 12894 6916 12900 6928
rect 12667 6888 12900 6916
rect 12667 6885 12679 6888
rect 12621 6879 12679 6885
rect 12894 6876 12900 6888
rect 12952 6876 12958 6928
rect 13832 6888 14228 6916
rect 6411 6820 6684 6848
rect 6411 6817 6423 6820
rect 6365 6811 6423 6817
rect 10870 6808 10876 6860
rect 10928 6808 10934 6860
rect 13832 6848 13860 6888
rect 12820 6820 13860 6848
rect 13924 6820 14136 6848
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6749 2467 6783
rect 2409 6743 2467 6749
rect 2685 6783 2743 6789
rect 2685 6749 2697 6783
rect 2731 6780 2743 6783
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2731 6752 2973 6780
rect 2731 6749 2743 6752
rect 2685 6743 2743 6749
rect 2961 6749 2973 6752
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 2424 6712 2452 6743
rect 3142 6740 3148 6792
rect 3200 6780 3206 6792
rect 3513 6783 3571 6789
rect 3513 6780 3525 6783
rect 3200 6752 3525 6780
rect 3200 6740 3206 6752
rect 3513 6749 3525 6752
rect 3559 6749 3571 6783
rect 3513 6743 3571 6749
rect 5810 6740 5816 6792
rect 5868 6780 5874 6792
rect 6089 6783 6147 6789
rect 6089 6780 6101 6783
rect 5868 6752 6101 6780
rect 5868 6740 5874 6752
rect 6089 6749 6101 6752
rect 6135 6749 6147 6783
rect 6089 6743 6147 6749
rect 6270 6740 6276 6792
rect 6328 6780 6334 6792
rect 6454 6780 6460 6792
rect 6328 6752 6460 6780
rect 6328 6740 6334 6752
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 8294 6740 8300 6792
rect 8352 6782 8358 6792
rect 8352 6754 8432 6782
rect 8352 6740 8358 6754
rect 5718 6712 5724 6724
rect 2424 6684 5724 6712
rect 5718 6672 5724 6684
rect 5776 6672 5782 6724
rect 7006 6672 7012 6724
rect 7064 6712 7070 6724
rect 7834 6712 7840 6724
rect 7064 6684 7840 6712
rect 7064 6672 7070 6684
rect 7834 6672 7840 6684
rect 7892 6672 7898 6724
rect 8404 6712 8432 6754
rect 8478 6740 8484 6792
rect 8536 6740 8542 6792
rect 9398 6740 9404 6792
rect 9456 6740 9462 6792
rect 9582 6740 9588 6792
rect 9640 6740 9646 6792
rect 9861 6783 9919 6789
rect 9861 6749 9873 6783
rect 9907 6780 9919 6783
rect 10134 6780 10140 6792
rect 9907 6752 10140 6780
rect 9907 6749 9919 6752
rect 9861 6743 9919 6749
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 8662 6712 8668 6724
rect 8404 6684 8668 6712
rect 8662 6672 8668 6684
rect 8720 6712 8726 6724
rect 9217 6715 9275 6721
rect 9217 6712 9229 6715
rect 8720 6684 9229 6712
rect 8720 6672 8726 6684
rect 9217 6681 9229 6684
rect 9263 6681 9275 6715
rect 9217 6675 9275 6681
rect 9324 6684 11560 6712
rect 1946 6604 1952 6656
rect 2004 6644 2010 6656
rect 2225 6647 2283 6653
rect 2225 6644 2237 6647
rect 2004 6616 2237 6644
rect 2004 6604 2010 6616
rect 2225 6613 2237 6616
rect 2271 6613 2283 6647
rect 2225 6607 2283 6613
rect 6638 6604 6644 6656
rect 6696 6644 6702 6656
rect 9324 6644 9352 6684
rect 6696 6616 9352 6644
rect 6696 6604 6702 6616
rect 9398 6604 9404 6656
rect 9456 6644 9462 6656
rect 9677 6647 9735 6653
rect 9677 6644 9689 6647
rect 9456 6616 9689 6644
rect 9456 6604 9462 6616
rect 9677 6613 9689 6616
rect 9723 6613 9735 6647
rect 11532 6644 11560 6684
rect 12158 6672 12164 6724
rect 12216 6672 12222 6724
rect 12820 6656 12848 6820
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6780 12955 6783
rect 12986 6780 12992 6792
rect 12943 6752 12992 6780
rect 12943 6749 12955 6752
rect 12897 6743 12955 6749
rect 12986 6740 12992 6752
rect 13044 6740 13050 6792
rect 13740 6789 13768 6820
rect 13924 6789 13952 6820
rect 13081 6783 13139 6789
rect 13081 6749 13093 6783
rect 13127 6749 13139 6783
rect 13081 6743 13139 6749
rect 13725 6783 13783 6789
rect 13725 6749 13737 6783
rect 13771 6749 13783 6783
rect 13725 6743 13783 6749
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6749 13967 6783
rect 13909 6743 13967 6749
rect 13096 6712 13124 6743
rect 13998 6740 14004 6792
rect 14056 6740 14062 6792
rect 14108 6789 14136 6820
rect 14093 6783 14151 6789
rect 14093 6749 14105 6783
rect 14139 6749 14151 6783
rect 14200 6780 14228 6888
rect 14366 6876 14372 6928
rect 14424 6876 14430 6928
rect 21560 6916 21588 6947
rect 21726 6944 21732 6996
rect 21784 6944 21790 6996
rect 22738 6984 22744 6996
rect 22066 6956 22744 6984
rect 22066 6916 22094 6956
rect 22738 6944 22744 6956
rect 22796 6944 22802 6996
rect 23842 6984 23848 6996
rect 23032 6956 23848 6984
rect 21560 6888 22094 6916
rect 22370 6876 22376 6928
rect 22428 6876 22434 6928
rect 22922 6876 22928 6928
rect 22980 6876 22986 6928
rect 15102 6808 15108 6860
rect 15160 6808 15166 6860
rect 15565 6851 15623 6857
rect 15565 6817 15577 6851
rect 15611 6848 15623 6851
rect 15654 6848 15660 6860
rect 15611 6820 15660 6848
rect 15611 6817 15623 6820
rect 15565 6811 15623 6817
rect 15654 6808 15660 6820
rect 15712 6808 15718 6860
rect 16301 6851 16359 6857
rect 16301 6848 16313 6851
rect 15764 6820 16313 6848
rect 14829 6783 14887 6789
rect 14829 6780 14841 6783
rect 14200 6752 14841 6780
rect 14093 6743 14151 6749
rect 14829 6749 14841 6752
rect 14875 6749 14887 6783
rect 14829 6743 14887 6749
rect 14016 6712 14044 6740
rect 13096 6684 14044 6712
rect 12526 6644 12532 6656
rect 11532 6616 12532 6644
rect 9677 6607 9735 6613
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 12802 6604 12808 6656
rect 12860 6604 12866 6656
rect 14108 6644 14136 6743
rect 14642 6672 14648 6724
rect 14700 6712 14706 6724
rect 15764 6712 15792 6820
rect 16301 6817 16313 6820
rect 16347 6848 16359 6851
rect 16347 6820 16528 6848
rect 16347 6817 16359 6820
rect 16301 6811 16359 6817
rect 16500 6780 16528 6820
rect 16574 6808 16580 6860
rect 16632 6848 16638 6860
rect 16669 6851 16727 6857
rect 16669 6848 16681 6851
rect 16632 6820 16681 6848
rect 16632 6808 16638 6820
rect 16669 6817 16681 6820
rect 16715 6817 16727 6851
rect 17037 6851 17095 6857
rect 17037 6848 17049 6851
rect 16669 6811 16727 6817
rect 16776 6820 17049 6848
rect 16776 6780 16804 6820
rect 17037 6817 17049 6820
rect 17083 6848 17095 6851
rect 17494 6848 17500 6860
rect 17083 6820 17500 6848
rect 17083 6817 17095 6820
rect 17037 6811 17095 6817
rect 17494 6808 17500 6820
rect 17552 6808 17558 6860
rect 22940 6848 22968 6876
rect 23032 6857 23060 6956
rect 23842 6944 23848 6956
rect 23900 6944 23906 6996
rect 24121 6987 24179 6993
rect 24121 6953 24133 6987
rect 24167 6984 24179 6987
rect 24397 6987 24455 6993
rect 24397 6984 24409 6987
rect 24167 6956 24409 6984
rect 24167 6953 24179 6956
rect 24121 6947 24179 6953
rect 24397 6953 24409 6956
rect 24443 6953 24455 6987
rect 24397 6947 24455 6953
rect 25130 6944 25136 6996
rect 25188 6944 25194 6996
rect 23106 6876 23112 6928
rect 23164 6916 23170 6928
rect 23164 6888 24532 6916
rect 23164 6876 23170 6888
rect 24504 6857 24532 6888
rect 22204 6820 22968 6848
rect 23017 6851 23075 6857
rect 22204 6792 22232 6820
rect 23017 6817 23029 6851
rect 23063 6817 23075 6851
rect 23017 6811 23075 6817
rect 24489 6851 24547 6857
rect 24489 6817 24501 6851
rect 24535 6817 24547 6851
rect 24489 6811 24547 6817
rect 25406 6808 25412 6860
rect 25464 6848 25470 6860
rect 25685 6851 25743 6857
rect 25685 6848 25697 6851
rect 25464 6820 25697 6848
rect 25464 6808 25470 6820
rect 25685 6817 25697 6820
rect 25731 6817 25743 6851
rect 25685 6811 25743 6817
rect 14700 6684 15792 6712
rect 16408 6712 16436 6766
rect 16500 6752 16804 6780
rect 16853 6783 16911 6789
rect 16853 6749 16865 6783
rect 16899 6780 16911 6783
rect 17405 6783 17463 6789
rect 17405 6780 17417 6783
rect 16899 6752 16988 6780
rect 16899 6749 16911 6752
rect 16853 6743 16911 6749
rect 16960 6712 16988 6752
rect 16408 6684 16988 6712
rect 14700 6672 14706 6684
rect 16960 6656 16988 6684
rect 17052 6752 17417 6780
rect 17052 6656 17080 6752
rect 17405 6749 17417 6752
rect 17451 6749 17463 6783
rect 17405 6743 17463 6749
rect 17589 6783 17647 6789
rect 17589 6749 17601 6783
rect 17635 6780 17647 6783
rect 17635 6752 18000 6780
rect 17635 6749 17647 6752
rect 17589 6743 17647 6749
rect 17972 6656 18000 6752
rect 18782 6740 18788 6792
rect 18840 6740 18846 6792
rect 21637 6783 21695 6789
rect 21637 6749 21649 6783
rect 21683 6749 21695 6783
rect 21637 6743 21695 6749
rect 21652 6712 21680 6743
rect 21910 6740 21916 6792
rect 21968 6740 21974 6792
rect 22094 6789 22100 6792
rect 22078 6783 22100 6789
rect 22078 6749 22090 6783
rect 22078 6743 22100 6749
rect 22094 6740 22100 6743
rect 22152 6740 22158 6792
rect 22186 6740 22192 6792
rect 22244 6740 22250 6792
rect 22278 6740 22284 6792
rect 22336 6780 22342 6792
rect 22336 6774 22876 6780
rect 22922 6774 22928 6792
rect 22336 6752 22928 6774
rect 22336 6740 22342 6752
rect 22848 6746 22928 6752
rect 22922 6740 22928 6746
rect 22980 6740 22986 6792
rect 23106 6740 23112 6792
rect 23164 6780 23170 6792
rect 23477 6783 23535 6789
rect 23477 6780 23489 6783
rect 23164 6752 23489 6780
rect 23164 6740 23170 6752
rect 23477 6749 23489 6752
rect 23523 6749 23535 6783
rect 23477 6743 23535 6749
rect 24397 6783 24455 6789
rect 24397 6749 24409 6783
rect 24443 6749 24455 6783
rect 24397 6743 24455 6749
rect 22554 6712 22560 6724
rect 21652 6684 22560 6712
rect 22554 6672 22560 6684
rect 22612 6672 22618 6724
rect 24412 6712 24440 6743
rect 23216 6684 24440 6712
rect 15930 6644 15936 6656
rect 14108 6616 15936 6644
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 16942 6604 16948 6656
rect 17000 6604 17006 6656
rect 17034 6604 17040 6656
rect 17092 6604 17098 6656
rect 17402 6604 17408 6656
rect 17460 6604 17466 6656
rect 17954 6604 17960 6656
rect 18012 6604 18018 6656
rect 18598 6604 18604 6656
rect 18656 6604 18662 6656
rect 21177 6647 21235 6653
rect 21177 6613 21189 6647
rect 21223 6644 21235 6647
rect 21910 6644 21916 6656
rect 21223 6616 21916 6644
rect 21223 6613 21235 6616
rect 21177 6607 21235 6613
rect 21910 6604 21916 6616
rect 21968 6644 21974 6656
rect 23216 6644 23244 6684
rect 21968 6616 23244 6644
rect 21968 6604 21974 6616
rect 23842 6604 23848 6656
rect 23900 6644 23906 6656
rect 24765 6647 24823 6653
rect 24765 6644 24777 6647
rect 23900 6616 24777 6644
rect 23900 6604 23906 6616
rect 24765 6613 24777 6616
rect 24811 6613 24823 6647
rect 24765 6607 24823 6613
rect 1104 6554 26472 6576
rect 1104 6502 7252 6554
rect 7304 6502 7316 6554
rect 7368 6502 7380 6554
rect 7432 6502 7444 6554
rect 7496 6502 7508 6554
rect 7560 6502 13554 6554
rect 13606 6502 13618 6554
rect 13670 6502 13682 6554
rect 13734 6502 13746 6554
rect 13798 6502 13810 6554
rect 13862 6502 19856 6554
rect 19908 6502 19920 6554
rect 19972 6502 19984 6554
rect 20036 6502 20048 6554
rect 20100 6502 20112 6554
rect 20164 6502 26158 6554
rect 26210 6502 26222 6554
rect 26274 6502 26286 6554
rect 26338 6502 26350 6554
rect 26402 6502 26414 6554
rect 26466 6502 26472 6554
rect 1104 6480 26472 6502
rect 1946 6440 1952 6452
rect 1688 6412 1952 6440
rect 1688 6381 1716 6412
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 6086 6400 6092 6452
rect 6144 6440 6150 6452
rect 6181 6443 6239 6449
rect 6181 6440 6193 6443
rect 6144 6412 6193 6440
rect 6144 6400 6150 6412
rect 6181 6409 6193 6412
rect 6227 6409 6239 6443
rect 6181 6403 6239 6409
rect 6546 6400 6552 6452
rect 6604 6400 6610 6452
rect 7929 6443 7987 6449
rect 7929 6409 7941 6443
rect 7975 6440 7987 6443
rect 8294 6440 8300 6452
rect 7975 6412 8300 6440
rect 7975 6409 7987 6412
rect 7929 6403 7987 6409
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 8478 6400 8484 6452
rect 8536 6440 8542 6452
rect 8573 6443 8631 6449
rect 8573 6440 8585 6443
rect 8536 6412 8585 6440
rect 8536 6400 8542 6412
rect 8573 6409 8585 6412
rect 8619 6409 8631 6443
rect 8573 6403 8631 6409
rect 11330 6400 11336 6452
rect 11388 6440 11394 6452
rect 11882 6440 11888 6452
rect 11388 6412 11888 6440
rect 11388 6400 11394 6412
rect 11882 6400 11888 6412
rect 11940 6440 11946 6452
rect 11977 6443 12035 6449
rect 11977 6440 11989 6443
rect 11940 6412 11989 6440
rect 11940 6400 11946 6412
rect 11977 6409 11989 6412
rect 12023 6409 12035 6443
rect 11977 6403 12035 6409
rect 12434 6400 12440 6452
rect 12492 6400 12498 6452
rect 12986 6400 12992 6452
rect 13044 6440 13050 6452
rect 13173 6443 13231 6449
rect 13173 6440 13185 6443
rect 13044 6412 13185 6440
rect 13044 6400 13050 6412
rect 13173 6409 13185 6412
rect 13219 6409 13231 6443
rect 13173 6403 13231 6409
rect 13725 6443 13783 6449
rect 13725 6409 13737 6443
rect 13771 6440 13783 6443
rect 13998 6440 14004 6452
rect 13771 6412 14004 6440
rect 13771 6409 13783 6412
rect 13725 6403 13783 6409
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 16942 6400 16948 6452
rect 17000 6400 17006 6452
rect 17402 6400 17408 6452
rect 17460 6400 17466 6452
rect 17494 6400 17500 6452
rect 17552 6440 17558 6452
rect 19518 6440 19524 6452
rect 17552 6412 19524 6440
rect 17552 6400 17558 6412
rect 19518 6400 19524 6412
rect 19576 6440 19582 6452
rect 20073 6443 20131 6449
rect 20073 6440 20085 6443
rect 19576 6412 20085 6440
rect 19576 6400 19582 6412
rect 20073 6409 20085 6412
rect 20119 6409 20131 6443
rect 22370 6440 22376 6452
rect 20073 6403 20131 6409
rect 21652 6412 22376 6440
rect 1673 6375 1731 6381
rect 1673 6341 1685 6375
rect 1719 6341 1731 6375
rect 9309 6375 9367 6381
rect 1673 6335 1731 6341
rect 7760 6344 8432 6372
rect 1394 6264 1400 6316
rect 1452 6264 1458 6316
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3418 6304 3424 6316
rect 2832 6276 3424 6304
rect 2832 6264 2838 6276
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6304 5595 6307
rect 5626 6304 5632 6316
rect 5583 6276 5632 6304
rect 5583 6273 5595 6276
rect 5537 6267 5595 6273
rect 5626 6264 5632 6276
rect 5684 6304 5690 6316
rect 7760 6313 7788 6344
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 5684 6276 6377 6304
rect 5684 6264 5690 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 7745 6307 7803 6313
rect 7745 6273 7757 6307
rect 7791 6273 7803 6307
rect 7745 6267 7803 6273
rect 8021 6307 8079 6313
rect 8021 6273 8033 6307
rect 8067 6304 8079 6307
rect 8113 6307 8171 6313
rect 8113 6304 8125 6307
rect 8067 6276 8125 6304
rect 8067 6273 8079 6276
rect 8021 6267 8079 6273
rect 8113 6273 8125 6276
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 5258 6196 5264 6248
rect 5316 6196 5322 6248
rect 6564 6236 6592 6267
rect 5828 6208 6592 6236
rect 5828 6180 5856 6208
rect 6914 6196 6920 6248
rect 6972 6196 6978 6248
rect 5810 6128 5816 6180
rect 5868 6128 5874 6180
rect 8128 6112 8156 6267
rect 3142 6060 3148 6112
rect 3200 6060 3206 6112
rect 6178 6060 6184 6112
rect 6236 6100 6242 6112
rect 7561 6103 7619 6109
rect 7561 6100 7573 6103
rect 6236 6072 7573 6100
rect 6236 6060 6242 6072
rect 7561 6069 7573 6072
rect 7607 6069 7619 6103
rect 7561 6063 7619 6069
rect 8110 6060 8116 6112
rect 8168 6060 8174 6112
rect 8404 6109 8432 6344
rect 9309 6341 9321 6375
rect 9355 6372 9367 6375
rect 9398 6372 9404 6384
rect 9355 6344 9404 6372
rect 9355 6341 9367 6344
rect 9309 6335 9367 6341
rect 9398 6332 9404 6344
rect 9456 6332 9462 6384
rect 12069 6375 12127 6381
rect 12069 6341 12081 6375
rect 12115 6372 12127 6375
rect 12894 6372 12900 6384
rect 12115 6344 12900 6372
rect 12115 6341 12127 6344
rect 12069 6335 12127 6341
rect 12894 6332 12900 6344
rect 12952 6332 12958 6384
rect 16114 6372 16120 6384
rect 13369 6344 13860 6372
rect 9033 6307 9091 6313
rect 9033 6273 9045 6307
rect 9079 6273 9091 6307
rect 9033 6267 9091 6273
rect 9048 6236 9076 6267
rect 10318 6264 10324 6316
rect 10376 6304 10382 6316
rect 13369 6313 13397 6344
rect 13832 6313 13860 6344
rect 14200 6344 16120 6372
rect 13357 6307 13415 6313
rect 10376 6276 12434 6304
rect 10376 6264 10382 6276
rect 10870 6236 10876 6248
rect 9048 6208 10876 6236
rect 10870 6196 10876 6208
rect 10928 6196 10934 6248
rect 11882 6196 11888 6248
rect 11940 6196 11946 6248
rect 12406 6236 12434 6276
rect 13357 6273 13369 6307
rect 13403 6273 13415 6307
rect 13357 6267 13415 6273
rect 13541 6307 13599 6313
rect 13541 6273 13553 6307
rect 13587 6304 13599 6307
rect 13633 6307 13691 6313
rect 13633 6304 13645 6307
rect 13587 6276 13645 6304
rect 13587 6273 13599 6276
rect 13541 6267 13599 6273
rect 13633 6273 13645 6276
rect 13679 6273 13691 6307
rect 13633 6267 13691 6273
rect 13817 6307 13875 6313
rect 13817 6273 13829 6307
rect 13863 6304 13875 6307
rect 13998 6304 14004 6316
rect 13863 6276 14004 6304
rect 13863 6273 13875 6276
rect 13817 6267 13875 6273
rect 13648 6236 13676 6267
rect 13998 6264 14004 6276
rect 14056 6264 14062 6316
rect 14200 6313 14228 6344
rect 16114 6332 16120 6344
rect 16172 6332 16178 6384
rect 14185 6307 14243 6313
rect 14185 6273 14197 6307
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 14200 6236 14228 6267
rect 14642 6264 14648 6316
rect 14700 6264 14706 6316
rect 14921 6307 14979 6313
rect 14921 6273 14933 6307
rect 14967 6273 14979 6307
rect 14921 6267 14979 6273
rect 12406 6208 13216 6236
rect 13648 6208 14228 6236
rect 8846 6128 8852 6180
rect 8904 6168 8910 6180
rect 8904 6140 9168 6168
rect 8904 6128 8910 6140
rect 8389 6103 8447 6109
rect 8389 6069 8401 6103
rect 8435 6100 8447 6103
rect 8938 6100 8944 6112
rect 8435 6072 8944 6100
rect 8435 6069 8447 6072
rect 8389 6063 8447 6069
rect 8938 6060 8944 6072
rect 8996 6060 9002 6112
rect 9140 6100 9168 6140
rect 10318 6100 10324 6112
rect 9140 6072 10324 6100
rect 10318 6060 10324 6072
rect 10376 6100 10382 6112
rect 10781 6103 10839 6109
rect 10781 6100 10793 6103
rect 10376 6072 10793 6100
rect 10376 6060 10382 6072
rect 10781 6069 10793 6072
rect 10827 6069 10839 6103
rect 13188 6100 13216 6208
rect 14458 6196 14464 6248
rect 14516 6196 14522 6248
rect 13906 6128 13912 6180
rect 13964 6168 13970 6180
rect 14936 6168 14964 6267
rect 15286 6264 15292 6316
rect 15344 6264 15350 6316
rect 15381 6307 15439 6313
rect 15381 6273 15393 6307
rect 15427 6304 15439 6307
rect 16960 6304 16988 6400
rect 17052 6344 17264 6372
rect 17052 6316 17080 6344
rect 15427 6276 16988 6304
rect 15427 6273 15439 6276
rect 15381 6267 15439 6273
rect 17034 6264 17040 6316
rect 17092 6264 17098 6316
rect 17236 6313 17264 6344
rect 17129 6307 17187 6313
rect 17129 6273 17141 6307
rect 17175 6273 17187 6307
rect 17129 6267 17187 6273
rect 17221 6307 17279 6313
rect 17221 6273 17233 6307
rect 17267 6273 17279 6307
rect 17221 6267 17279 6273
rect 17144 6236 17172 6267
rect 17420 6245 17448 6400
rect 18046 6332 18052 6384
rect 18104 6332 18110 6384
rect 19058 6332 19064 6384
rect 19116 6332 19122 6384
rect 17497 6307 17555 6313
rect 17497 6273 17509 6307
rect 17543 6304 17555 6307
rect 18064 6304 18092 6332
rect 17543 6276 18092 6304
rect 17543 6273 17555 6276
rect 17497 6267 17555 6273
rect 18322 6264 18328 6316
rect 18380 6264 18386 6316
rect 21652 6313 21680 6412
rect 22370 6400 22376 6412
rect 22428 6400 22434 6452
rect 23658 6400 23664 6452
rect 23716 6440 23722 6452
rect 23716 6412 25452 6440
rect 23716 6400 23722 6412
rect 22830 6332 22836 6384
rect 22888 6372 22894 6384
rect 22888 6344 23966 6372
rect 22888 6332 22894 6344
rect 21637 6307 21695 6313
rect 21637 6273 21649 6307
rect 21683 6273 21695 6307
rect 21637 6267 21695 6273
rect 23569 6307 23627 6313
rect 23569 6273 23581 6307
rect 23615 6304 23627 6307
rect 23658 6304 23664 6316
rect 23615 6276 23664 6304
rect 23615 6273 23627 6276
rect 23569 6267 23627 6273
rect 23658 6264 23664 6276
rect 23716 6264 23722 6316
rect 25424 6313 25452 6412
rect 25409 6307 25467 6313
rect 25409 6273 25421 6307
rect 25455 6273 25467 6307
rect 25409 6267 25467 6273
rect 17405 6239 17463 6245
rect 17144 6208 17264 6236
rect 13964 6140 14964 6168
rect 17236 6168 17264 6208
rect 17405 6205 17417 6239
rect 17451 6205 17463 6239
rect 17405 6199 17463 6205
rect 18598 6196 18604 6248
rect 18656 6196 18662 6248
rect 23293 6239 23351 6245
rect 23293 6205 23305 6239
rect 23339 6236 23351 6239
rect 23339 6208 23520 6236
rect 23339 6205 23351 6208
rect 23293 6199 23351 6205
rect 17589 6171 17647 6177
rect 17589 6168 17601 6171
rect 17236 6140 17601 6168
rect 13964 6128 13970 6140
rect 17589 6137 17601 6140
rect 17635 6137 17647 6171
rect 17589 6131 17647 6137
rect 17681 6171 17739 6177
rect 17681 6137 17693 6171
rect 17727 6168 17739 6171
rect 17954 6168 17960 6180
rect 17727 6140 17960 6168
rect 17727 6137 17739 6140
rect 17681 6131 17739 6137
rect 14090 6100 14096 6112
rect 13188 6072 14096 6100
rect 10781 6063 10839 6069
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 14274 6060 14280 6112
rect 14332 6060 14338 6112
rect 14829 6103 14887 6109
rect 14829 6069 14841 6103
rect 14875 6100 14887 6103
rect 15013 6103 15071 6109
rect 15013 6100 15025 6103
rect 14875 6072 15025 6100
rect 14875 6069 14887 6072
rect 14829 6063 14887 6069
rect 15013 6069 15025 6072
rect 15059 6069 15071 6103
rect 15013 6063 15071 6069
rect 15562 6060 15568 6112
rect 15620 6060 15626 6112
rect 16574 6060 16580 6112
rect 16632 6100 16638 6112
rect 17696 6100 17724 6131
rect 17954 6128 17960 6140
rect 18012 6128 18018 6180
rect 22002 6168 22008 6180
rect 21284 6140 22008 6168
rect 21284 6112 21312 6140
rect 22002 6128 22008 6140
rect 22060 6168 22066 6180
rect 22060 6140 22324 6168
rect 22060 6128 22066 6140
rect 16632 6072 17724 6100
rect 16632 6060 16638 6072
rect 21266 6060 21272 6112
rect 21324 6060 21330 6112
rect 21542 6060 21548 6112
rect 21600 6060 21606 6112
rect 21821 6103 21879 6109
rect 21821 6069 21833 6103
rect 21867 6100 21879 6103
rect 22186 6100 22192 6112
rect 21867 6072 22192 6100
rect 21867 6069 21879 6072
rect 21821 6063 21879 6069
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 22296 6100 22324 6140
rect 23492 6112 23520 6208
rect 25130 6196 25136 6248
rect 25188 6196 25194 6248
rect 23566 6128 23572 6180
rect 23624 6168 23630 6180
rect 23661 6171 23719 6177
rect 23661 6168 23673 6171
rect 23624 6140 23673 6168
rect 23624 6128 23630 6140
rect 23661 6137 23673 6140
rect 23707 6137 23719 6171
rect 23661 6131 23719 6137
rect 22830 6100 22836 6112
rect 22296 6072 22836 6100
rect 22830 6060 22836 6072
rect 22888 6060 22894 6112
rect 23474 6060 23480 6112
rect 23532 6060 23538 6112
rect 1104 6010 26312 6032
rect 1104 5958 4101 6010
rect 4153 5958 4165 6010
rect 4217 5958 4229 6010
rect 4281 5958 4293 6010
rect 4345 5958 4357 6010
rect 4409 5958 10403 6010
rect 10455 5958 10467 6010
rect 10519 5958 10531 6010
rect 10583 5958 10595 6010
rect 10647 5958 10659 6010
rect 10711 5958 16705 6010
rect 16757 5958 16769 6010
rect 16821 5958 16833 6010
rect 16885 5958 16897 6010
rect 16949 5958 16961 6010
rect 17013 5958 23007 6010
rect 23059 5958 23071 6010
rect 23123 5958 23135 6010
rect 23187 5958 23199 6010
rect 23251 5958 23263 6010
rect 23315 5958 26312 6010
rect 1104 5936 26312 5958
rect 5258 5856 5264 5908
rect 5316 5856 5322 5908
rect 6733 5899 6791 5905
rect 6733 5865 6745 5899
rect 6779 5896 6791 5899
rect 6914 5896 6920 5908
rect 6779 5868 6920 5896
rect 6779 5865 6791 5868
rect 6733 5859 6791 5865
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 8110 5856 8116 5908
rect 8168 5896 8174 5908
rect 8205 5899 8263 5905
rect 8205 5896 8217 5899
rect 8168 5868 8217 5896
rect 8168 5856 8174 5868
rect 8205 5865 8217 5868
rect 8251 5865 8263 5899
rect 8205 5859 8263 5865
rect 8938 5856 8944 5908
rect 8996 5856 9002 5908
rect 9122 5856 9128 5908
rect 9180 5856 9186 5908
rect 9232 5868 10088 5896
rect 5718 5828 5724 5840
rect 5000 5800 5724 5828
rect 5000 5769 5028 5800
rect 5718 5788 5724 5800
rect 5776 5828 5782 5840
rect 9232 5828 9260 5868
rect 5776 5800 6776 5828
rect 5776 5788 5782 5800
rect 4985 5763 5043 5769
rect 4985 5729 4997 5763
rect 5031 5729 5043 5763
rect 4985 5723 5043 5729
rect 5534 5720 5540 5772
rect 5592 5720 5598 5772
rect 5902 5760 5908 5772
rect 5736 5732 5908 5760
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5692 4951 5695
rect 5736 5692 5764 5732
rect 5902 5720 5908 5732
rect 5960 5760 5966 5772
rect 5960 5732 6316 5760
rect 5960 5720 5966 5732
rect 4939 5664 5764 5692
rect 5813 5695 5871 5701
rect 4939 5661 4951 5664
rect 4893 5655 4951 5661
rect 5813 5661 5825 5695
rect 5859 5692 5871 5695
rect 6178 5692 6184 5704
rect 5859 5664 6184 5692
rect 5859 5661 5871 5664
rect 5813 5655 5871 5661
rect 6178 5652 6184 5664
rect 6236 5652 6242 5704
rect 6288 5692 6316 5732
rect 6454 5720 6460 5772
rect 6512 5720 6518 5772
rect 6748 5704 6776 5800
rect 7576 5800 9260 5828
rect 7576 5769 7604 5800
rect 9674 5788 9680 5840
rect 9732 5788 9738 5840
rect 10060 5828 10088 5868
rect 10134 5856 10140 5908
rect 10192 5856 10198 5908
rect 11606 5856 11612 5908
rect 11664 5856 11670 5908
rect 12802 5896 12808 5908
rect 12406 5868 12808 5896
rect 11425 5831 11483 5837
rect 11425 5828 11437 5831
rect 9876 5800 9996 5828
rect 10060 5800 11437 5828
rect 7561 5763 7619 5769
rect 7561 5729 7573 5763
rect 7607 5729 7619 5763
rect 7561 5723 7619 5729
rect 9490 5720 9496 5772
rect 9548 5760 9554 5772
rect 9692 5760 9720 5788
rect 9876 5760 9904 5800
rect 9968 5769 9996 5800
rect 11425 5797 11437 5800
rect 11471 5797 11483 5831
rect 11425 5791 11483 5797
rect 9548 5732 9904 5760
rect 9953 5763 10011 5769
rect 9548 5720 9554 5732
rect 9953 5729 9965 5763
rect 9999 5729 10011 5763
rect 9953 5723 10011 5729
rect 10042 5720 10048 5772
rect 10100 5760 10106 5772
rect 10597 5763 10655 5769
rect 10597 5760 10609 5763
rect 10100 5732 10609 5760
rect 10100 5720 10106 5732
rect 10597 5729 10609 5732
rect 10643 5729 10655 5763
rect 10597 5723 10655 5729
rect 6549 5695 6607 5701
rect 6549 5692 6561 5695
rect 6288 5664 6561 5692
rect 6549 5661 6561 5664
rect 6595 5692 6607 5695
rect 6638 5692 6644 5704
rect 6595 5664 6644 5692
rect 6595 5661 6607 5664
rect 6549 5655 6607 5661
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 6730 5652 6736 5704
rect 6788 5692 6794 5704
rect 7076 5695 7134 5701
rect 7076 5692 7088 5695
rect 6788 5664 7088 5692
rect 6788 5652 6794 5664
rect 7076 5661 7088 5664
rect 7122 5661 7134 5695
rect 7076 5655 7134 5661
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5661 8447 5695
rect 8389 5655 8447 5661
rect 8665 5695 8723 5701
rect 8665 5661 8677 5695
rect 8711 5692 8723 5695
rect 9214 5692 9220 5704
rect 8711 5664 9220 5692
rect 8711 5661 8723 5664
rect 8665 5655 8723 5661
rect 6270 5584 6276 5636
rect 6328 5624 6334 5636
rect 7193 5627 7251 5633
rect 7193 5624 7205 5627
rect 6328 5596 7205 5624
rect 6328 5584 6334 5596
rect 7193 5593 7205 5596
rect 7239 5593 7251 5627
rect 8404 5624 8432 5655
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 9674 5692 9680 5704
rect 9646 5652 9680 5692
rect 9732 5652 9738 5704
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5692 9919 5695
rect 10612 5692 10640 5723
rect 10686 5720 10692 5772
rect 10744 5720 10750 5772
rect 11701 5763 11759 5769
rect 11701 5729 11713 5763
rect 11747 5760 11759 5763
rect 12406 5760 12434 5868
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 13265 5899 13323 5905
rect 13265 5865 13277 5899
rect 13311 5896 13323 5899
rect 13998 5896 14004 5908
rect 13311 5868 14004 5896
rect 13311 5865 13323 5868
rect 13265 5859 13323 5865
rect 13998 5856 14004 5868
rect 14056 5856 14062 5908
rect 15562 5856 15568 5908
rect 15620 5856 15626 5908
rect 15930 5856 15936 5908
rect 15988 5856 15994 5908
rect 18782 5856 18788 5908
rect 18840 5896 18846 5908
rect 19245 5899 19303 5905
rect 19245 5896 19257 5899
rect 18840 5868 19257 5896
rect 18840 5856 18846 5868
rect 19245 5865 19257 5868
rect 19291 5865 19303 5899
rect 19245 5859 19303 5865
rect 22554 5856 22560 5908
rect 22612 5896 22618 5908
rect 22741 5899 22799 5905
rect 22741 5896 22753 5899
rect 22612 5868 22753 5896
rect 22612 5856 22618 5868
rect 22741 5865 22753 5868
rect 22787 5865 22799 5899
rect 22741 5859 22799 5865
rect 12820 5828 12848 5856
rect 15381 5831 15439 5837
rect 15381 5828 15393 5831
rect 12820 5800 15393 5828
rect 15381 5797 15393 5800
rect 15427 5797 15439 5831
rect 15381 5791 15439 5797
rect 11747 5732 12434 5760
rect 11747 5729 11759 5732
rect 11701 5723 11759 5729
rect 12526 5720 12532 5772
rect 12584 5760 12590 5772
rect 13081 5763 13139 5769
rect 12584 5732 12664 5760
rect 12584 5720 12590 5732
rect 10778 5692 10784 5704
rect 9907 5664 10088 5692
rect 10612 5664 10784 5692
rect 9907 5661 9919 5664
rect 9861 5655 9919 5661
rect 9309 5627 9367 5633
rect 9309 5624 9321 5627
rect 8404 5596 9321 5624
rect 7193 5587 7251 5593
rect 9309 5593 9321 5596
rect 9355 5624 9367 5627
rect 9646 5624 9674 5652
rect 9355 5596 9674 5624
rect 9355 5593 9367 5596
rect 9309 5587 9367 5593
rect 6917 5559 6975 5565
rect 6917 5525 6929 5559
rect 6963 5556 6975 5559
rect 7006 5556 7012 5568
rect 6963 5528 7012 5556
rect 6963 5525 6975 5528
rect 6917 5519 6975 5525
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 7285 5559 7343 5565
rect 7285 5525 7297 5559
rect 7331 5556 7343 5559
rect 8110 5556 8116 5568
rect 7331 5528 8116 5556
rect 7331 5525 7343 5528
rect 7285 5519 7343 5525
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 8573 5559 8631 5565
rect 8573 5525 8585 5559
rect 8619 5556 8631 5559
rect 8938 5556 8944 5568
rect 8619 5528 8944 5556
rect 8619 5525 8631 5528
rect 8573 5519 8631 5525
rect 8938 5516 8944 5528
rect 8996 5516 9002 5568
rect 9109 5559 9167 5565
rect 9109 5525 9121 5559
rect 9155 5556 9167 5559
rect 9214 5556 9220 5568
rect 9155 5528 9220 5556
rect 9155 5525 9167 5528
rect 9109 5519 9167 5525
rect 9214 5516 9220 5528
rect 9272 5516 9278 5568
rect 9493 5559 9551 5565
rect 9493 5525 9505 5559
rect 9539 5556 9551 5559
rect 9582 5556 9588 5568
rect 9539 5528 9588 5556
rect 9539 5525 9551 5528
rect 9493 5519 9551 5525
rect 9582 5516 9588 5528
rect 9640 5556 9646 5568
rect 9674 5556 9680 5568
rect 9640 5528 9680 5556
rect 9640 5516 9646 5528
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 9950 5516 9956 5568
rect 10008 5556 10014 5568
rect 10060 5556 10088 5664
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 11793 5695 11851 5701
rect 11793 5661 11805 5695
rect 11839 5661 11851 5695
rect 12636 5692 12664 5732
rect 13081 5729 13093 5763
rect 13127 5760 13139 5763
rect 15580 5760 15608 5856
rect 19076 5800 19840 5828
rect 13127 5732 15608 5760
rect 13127 5729 13139 5732
rect 13081 5723 13139 5729
rect 17034 5720 17040 5772
rect 17092 5760 17098 5772
rect 17092 5732 18000 5760
rect 17092 5720 17098 5732
rect 13170 5692 13176 5704
rect 12636 5664 13176 5692
rect 11793 5655 11851 5661
rect 10008 5528 10088 5556
rect 10008 5516 10014 5528
rect 10318 5516 10324 5568
rect 10376 5556 10382 5568
rect 10505 5559 10563 5565
rect 10505 5556 10517 5559
rect 10376 5528 10517 5556
rect 10376 5516 10382 5528
rect 10505 5525 10517 5528
rect 10551 5525 10563 5559
rect 11808 5556 11836 5655
rect 13170 5652 13176 5664
rect 13228 5692 13234 5704
rect 13357 5695 13415 5701
rect 13357 5692 13369 5695
rect 13228 5664 13369 5692
rect 13228 5652 13234 5664
rect 13357 5661 13369 5664
rect 13403 5661 13415 5695
rect 13357 5655 13415 5661
rect 15565 5695 15623 5701
rect 15565 5661 15577 5695
rect 15611 5692 15623 5695
rect 15841 5695 15899 5701
rect 15841 5692 15853 5695
rect 15611 5664 15853 5692
rect 15611 5661 15623 5664
rect 15565 5655 15623 5661
rect 15841 5661 15853 5664
rect 15887 5692 15899 5695
rect 15930 5692 15936 5704
rect 15887 5664 15936 5692
rect 15887 5661 15899 5664
rect 15841 5655 15899 5661
rect 15930 5652 15936 5664
rect 15988 5652 15994 5704
rect 16025 5695 16083 5701
rect 16025 5661 16037 5695
rect 16071 5661 16083 5695
rect 16025 5655 16083 5661
rect 17589 5695 17647 5701
rect 17589 5661 17601 5695
rect 17635 5692 17647 5695
rect 17862 5692 17868 5704
rect 17635 5664 17868 5692
rect 17635 5661 17647 5664
rect 17589 5655 17647 5661
rect 15749 5627 15807 5633
rect 15749 5593 15761 5627
rect 15795 5624 15807 5627
rect 16040 5624 16068 5655
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 17972 5701 18000 5732
rect 18046 5720 18052 5772
rect 18104 5769 18110 5772
rect 18104 5763 18132 5769
rect 18120 5729 18132 5763
rect 18104 5723 18132 5729
rect 18104 5720 18110 5723
rect 18506 5720 18512 5772
rect 18564 5720 18570 5772
rect 18601 5763 18659 5769
rect 18601 5729 18613 5763
rect 18647 5760 18659 5763
rect 18966 5760 18972 5772
rect 18647 5732 18972 5760
rect 18647 5729 18659 5732
rect 18601 5723 18659 5729
rect 18966 5720 18972 5732
rect 19024 5720 19030 5772
rect 17957 5695 18015 5701
rect 17957 5661 17969 5695
rect 18003 5692 18015 5695
rect 18690 5692 18696 5704
rect 18003 5664 18696 5692
rect 18003 5661 18015 5664
rect 17957 5655 18015 5661
rect 18690 5652 18696 5664
rect 18748 5652 18754 5704
rect 18782 5652 18788 5704
rect 18840 5692 18846 5704
rect 19076 5692 19104 5800
rect 19518 5720 19524 5772
rect 19576 5720 19582 5772
rect 19610 5720 19616 5772
rect 19668 5760 19674 5772
rect 19812 5769 19840 5800
rect 19705 5763 19763 5769
rect 19705 5760 19717 5763
rect 19668 5732 19717 5760
rect 19668 5720 19674 5732
rect 19705 5729 19717 5732
rect 19751 5729 19763 5763
rect 19705 5723 19763 5729
rect 19797 5763 19855 5769
rect 19797 5729 19809 5763
rect 19843 5729 19855 5763
rect 19797 5723 19855 5729
rect 21542 5720 21548 5772
rect 21600 5760 21606 5772
rect 22189 5763 22247 5769
rect 22189 5760 22201 5763
rect 21600 5732 22201 5760
rect 21600 5720 21606 5732
rect 22189 5729 22201 5732
rect 22235 5729 22247 5763
rect 22189 5723 22247 5729
rect 22465 5763 22523 5769
rect 22465 5729 22477 5763
rect 22511 5760 22523 5763
rect 23658 5760 23664 5772
rect 22511 5732 23664 5760
rect 22511 5729 22523 5732
rect 22465 5723 22523 5729
rect 23658 5720 23664 5732
rect 23716 5720 23722 5772
rect 18840 5664 19104 5692
rect 18840 5652 18846 5664
rect 18414 5624 18420 5636
rect 15795 5596 17632 5624
rect 15795 5593 15807 5596
rect 15749 5587 15807 5593
rect 17604 5568 17632 5596
rect 17972 5596 18420 5624
rect 17972 5568 18000 5596
rect 18414 5584 18420 5596
rect 18472 5624 18478 5636
rect 19536 5624 19564 5720
rect 19613 5627 19671 5633
rect 19613 5624 19625 5627
rect 18472 5596 19472 5624
rect 19536 5596 19625 5624
rect 18472 5584 18478 5596
rect 12805 5559 12863 5565
rect 12805 5556 12817 5559
rect 11808 5528 12817 5556
rect 10505 5519 10563 5525
rect 12805 5525 12817 5528
rect 12851 5525 12863 5559
rect 12805 5519 12863 5525
rect 17586 5516 17592 5568
rect 17644 5516 17650 5568
rect 17865 5559 17923 5565
rect 17865 5525 17877 5559
rect 17911 5556 17923 5559
rect 17954 5556 17960 5568
rect 17911 5528 17960 5556
rect 17911 5525 17923 5528
rect 17865 5519 17923 5525
rect 17954 5516 17960 5528
rect 18012 5516 18018 5568
rect 18230 5516 18236 5568
rect 18288 5516 18294 5568
rect 18690 5516 18696 5568
rect 18748 5516 18754 5568
rect 19058 5516 19064 5568
rect 19116 5516 19122 5568
rect 19444 5556 19472 5596
rect 19613 5593 19625 5596
rect 19659 5593 19671 5627
rect 19613 5587 19671 5593
rect 20441 5627 20499 5633
rect 20441 5593 20453 5627
rect 20487 5593 20499 5627
rect 20441 5587 20499 5593
rect 20456 5556 20484 5587
rect 19444 5528 20484 5556
rect 21100 5556 21128 5678
rect 22738 5652 22744 5704
rect 22796 5692 22802 5704
rect 23017 5695 23075 5701
rect 23017 5692 23029 5695
rect 22796 5664 23029 5692
rect 22796 5652 22802 5664
rect 23017 5661 23029 5664
rect 23063 5661 23075 5695
rect 23017 5655 23075 5661
rect 21266 5556 21272 5568
rect 21100 5528 21272 5556
rect 21266 5516 21272 5528
rect 21324 5516 21330 5568
rect 22094 5516 22100 5568
rect 22152 5556 22158 5568
rect 22557 5559 22615 5565
rect 22557 5556 22569 5559
rect 22152 5528 22569 5556
rect 22152 5516 22158 5528
rect 22557 5525 22569 5528
rect 22603 5525 22615 5559
rect 22557 5519 22615 5525
rect 1104 5466 26472 5488
rect 1104 5414 7252 5466
rect 7304 5414 7316 5466
rect 7368 5414 7380 5466
rect 7432 5414 7444 5466
rect 7496 5414 7508 5466
rect 7560 5414 13554 5466
rect 13606 5414 13618 5466
rect 13670 5414 13682 5466
rect 13734 5414 13746 5466
rect 13798 5414 13810 5466
rect 13862 5414 19856 5466
rect 19908 5414 19920 5466
rect 19972 5414 19984 5466
rect 20036 5414 20048 5466
rect 20100 5414 20112 5466
rect 20164 5414 26158 5466
rect 26210 5414 26222 5466
rect 26274 5414 26286 5466
rect 26338 5414 26350 5466
rect 26402 5414 26414 5466
rect 26466 5414 26472 5466
rect 1104 5392 26472 5414
rect 4801 5355 4859 5361
rect 4801 5321 4813 5355
rect 4847 5352 4859 5355
rect 4847 5324 5488 5352
rect 4847 5321 4859 5324
rect 4801 5315 4859 5321
rect 5460 5284 5488 5324
rect 5534 5312 5540 5364
rect 5592 5312 5598 5364
rect 5626 5312 5632 5364
rect 5684 5312 5690 5364
rect 5997 5355 6055 5361
rect 5997 5321 6009 5355
rect 6043 5352 6055 5355
rect 6178 5352 6184 5364
rect 6043 5324 6184 5352
rect 6043 5321 6055 5324
rect 5997 5315 6055 5321
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 8110 5312 8116 5364
rect 8168 5312 8174 5364
rect 9033 5355 9091 5361
rect 9033 5352 9045 5355
rect 8956 5324 9045 5352
rect 4724 5256 5212 5284
rect 5460 5256 5856 5284
rect 4724 5225 4752 5256
rect 5184 5225 5212 5256
rect 4709 5219 4767 5225
rect 4709 5185 4721 5219
rect 4755 5185 4767 5219
rect 4709 5179 4767 5185
rect 4887 5219 4945 5225
rect 4887 5185 4899 5219
rect 4933 5185 4945 5219
rect 4887 5179 4945 5185
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5216 5227 5219
rect 5626 5216 5632 5228
rect 5215 5188 5632 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 3970 5108 3976 5160
rect 4028 5108 4034 5160
rect 4908 5148 4936 5179
rect 5626 5176 5632 5188
rect 5684 5176 5690 5228
rect 5828 5225 5856 5256
rect 6730 5244 6736 5296
rect 6788 5244 6794 5296
rect 8846 5284 8852 5296
rect 7484 5256 8852 5284
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 6086 5176 6092 5228
rect 6144 5176 6150 5228
rect 7006 5176 7012 5228
rect 7064 5176 7070 5228
rect 7484 5225 7512 5256
rect 8846 5244 8852 5256
rect 8904 5244 8910 5296
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5216 8355 5219
rect 8956 5216 8984 5324
rect 9033 5321 9045 5324
rect 9079 5352 9091 5355
rect 9214 5352 9220 5364
rect 9079 5324 9220 5352
rect 9079 5321 9091 5324
rect 9033 5315 9091 5321
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 9490 5312 9496 5364
rect 9548 5312 9554 5364
rect 9674 5312 9680 5364
rect 9732 5352 9738 5364
rect 11606 5352 11612 5364
rect 9732 5324 11612 5352
rect 9732 5312 9738 5324
rect 11606 5312 11612 5324
rect 11664 5312 11670 5364
rect 13262 5312 13268 5364
rect 13320 5352 13326 5364
rect 16574 5352 16580 5364
rect 13320 5324 16580 5352
rect 13320 5312 13326 5324
rect 9508 5284 9536 5312
rect 9140 5256 9536 5284
rect 8343 5188 8984 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 5261 5151 5319 5157
rect 5261 5148 5273 5151
rect 4908 5120 5273 5148
rect 5261 5117 5273 5120
rect 5307 5148 5319 5151
rect 6270 5148 6276 5160
rect 5307 5120 6276 5148
rect 5307 5117 5319 5120
rect 5261 5111 5319 5117
rect 6270 5108 6276 5120
rect 6328 5108 6334 5160
rect 8128 5148 8156 5179
rect 9030 5176 9036 5228
rect 9088 5176 9094 5228
rect 9140 5225 9168 5256
rect 9766 5244 9772 5296
rect 9824 5284 9830 5296
rect 10686 5284 10692 5296
rect 9824 5256 10692 5284
rect 9824 5244 9830 5256
rect 10686 5244 10692 5256
rect 10744 5244 10750 5296
rect 14274 5284 14280 5296
rect 12912 5256 14280 5284
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 9306 5176 9312 5228
rect 9364 5216 9370 5228
rect 9585 5219 9643 5225
rect 9585 5216 9597 5219
rect 9364 5188 9597 5216
rect 9364 5176 9370 5188
rect 9585 5185 9597 5188
rect 9631 5185 9643 5219
rect 9585 5179 9643 5185
rect 9674 5176 9680 5228
rect 9732 5216 9738 5228
rect 9950 5216 9956 5228
rect 9732 5188 9956 5216
rect 9732 5186 9775 5188
rect 9732 5176 9738 5186
rect 9950 5176 9956 5188
rect 10008 5176 10014 5228
rect 9048 5148 9076 5176
rect 8128 5120 9076 5148
rect 9858 5108 9864 5160
rect 9916 5148 9922 5160
rect 12912 5148 12940 5256
rect 12986 5176 12992 5228
rect 13044 5216 13050 5228
rect 13173 5219 13231 5225
rect 13173 5216 13185 5219
rect 13044 5188 13185 5216
rect 13044 5176 13050 5188
rect 13173 5185 13185 5188
rect 13219 5185 13231 5219
rect 13173 5179 13231 5185
rect 13262 5176 13268 5228
rect 13320 5176 13326 5228
rect 13464 5225 13492 5256
rect 14274 5244 14280 5256
rect 14332 5244 14338 5296
rect 16132 5225 16160 5324
rect 16574 5312 16580 5324
rect 16632 5312 16638 5364
rect 17586 5312 17592 5364
rect 17644 5312 17650 5364
rect 18141 5355 18199 5361
rect 18141 5321 18153 5355
rect 18187 5321 18199 5355
rect 18690 5352 18696 5364
rect 18141 5315 18199 5321
rect 18248 5324 18696 5352
rect 18156 5284 18184 5315
rect 18248 5293 18276 5324
rect 18690 5312 18696 5324
rect 18748 5352 18754 5364
rect 20349 5355 20407 5361
rect 20349 5352 20361 5355
rect 18748 5324 20361 5352
rect 18748 5312 18754 5324
rect 20349 5321 20361 5324
rect 20395 5321 20407 5355
rect 20349 5315 20407 5321
rect 23474 5312 23480 5364
rect 23532 5312 23538 5364
rect 16224 5256 17356 5284
rect 13449 5219 13507 5225
rect 13449 5185 13461 5219
rect 13495 5185 13507 5219
rect 13449 5179 13507 5185
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5185 16175 5219
rect 16117 5179 16175 5185
rect 9916 5120 12940 5148
rect 9916 5108 9922 5120
rect 3988 5080 4016 5108
rect 11422 5080 11428 5092
rect 3988 5052 11428 5080
rect 11422 5040 11428 5052
rect 11480 5040 11486 5092
rect 8846 4972 8852 5024
rect 8904 4972 8910 5024
rect 8938 4972 8944 5024
rect 8996 5012 9002 5024
rect 12618 5012 12624 5024
rect 8996 4984 12624 5012
rect 8996 4972 9002 4984
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 12710 4972 12716 5024
rect 12768 5012 12774 5024
rect 12805 5015 12863 5021
rect 12805 5012 12817 5015
rect 12768 4984 12817 5012
rect 12768 4972 12774 4984
rect 12805 4981 12817 4984
rect 12851 4981 12863 5015
rect 12912 5012 12940 5120
rect 13081 5151 13139 5157
rect 13081 5117 13093 5151
rect 13127 5148 13139 5151
rect 16025 5151 16083 5157
rect 16025 5148 16037 5151
rect 13127 5120 16037 5148
rect 13127 5117 13139 5120
rect 13081 5111 13139 5117
rect 16025 5117 16037 5120
rect 16071 5148 16083 5151
rect 16224 5148 16252 5256
rect 17034 5176 17040 5228
rect 17092 5176 17098 5228
rect 17328 5225 17356 5256
rect 17420 5256 17908 5284
rect 17420 5225 17448 5256
rect 17880 5228 17908 5256
rect 18064 5256 18184 5284
rect 18233 5287 18291 5293
rect 17129 5219 17187 5225
rect 17129 5185 17141 5219
rect 17175 5185 17187 5219
rect 17129 5179 17187 5185
rect 17313 5219 17371 5225
rect 17313 5185 17325 5219
rect 17359 5185 17371 5219
rect 17313 5179 17371 5185
rect 17405 5219 17463 5225
rect 17405 5185 17417 5219
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 17773 5219 17831 5225
rect 17773 5185 17785 5219
rect 17819 5185 17831 5219
rect 17773 5179 17831 5185
rect 17144 5148 17172 5179
rect 16071 5120 16252 5148
rect 17052 5120 17172 5148
rect 17788 5148 17816 5179
rect 17862 5176 17868 5228
rect 17920 5216 17926 5228
rect 18064 5225 18092 5256
rect 18233 5253 18245 5287
rect 18279 5253 18291 5287
rect 18233 5247 18291 5253
rect 18414 5244 18420 5296
rect 18472 5244 18478 5296
rect 21266 5284 21272 5296
rect 20102 5256 21272 5284
rect 21266 5244 21272 5256
rect 21324 5244 21330 5296
rect 17957 5219 18015 5225
rect 17957 5216 17969 5219
rect 17920 5188 17969 5216
rect 17920 5176 17926 5188
rect 17957 5185 17969 5188
rect 18003 5185 18015 5219
rect 17957 5179 18015 5185
rect 18049 5219 18107 5225
rect 18049 5185 18061 5219
rect 18095 5185 18107 5219
rect 18049 5179 18107 5185
rect 18138 5176 18144 5228
rect 18196 5176 18202 5228
rect 17788 5120 18276 5148
rect 16071 5117 16083 5120
rect 16025 5111 16083 5117
rect 17052 5080 17080 5120
rect 18248 5092 18276 5120
rect 18322 5108 18328 5160
rect 18380 5148 18386 5160
rect 18601 5151 18659 5157
rect 18601 5148 18613 5151
rect 18380 5120 18613 5148
rect 18380 5108 18386 5120
rect 18601 5117 18613 5120
rect 18647 5117 18659 5151
rect 18601 5111 18659 5117
rect 18877 5151 18935 5157
rect 18877 5117 18889 5151
rect 18923 5148 18935 5151
rect 18966 5148 18972 5160
rect 18923 5120 18972 5148
rect 18923 5117 18935 5120
rect 18877 5111 18935 5117
rect 18138 5080 18144 5092
rect 17052 5052 18144 5080
rect 18138 5040 18144 5052
rect 18196 5040 18202 5092
rect 18230 5040 18236 5092
rect 18288 5040 18294 5092
rect 12989 5015 13047 5021
rect 12989 5012 13001 5015
rect 12912 4984 13001 5012
rect 12805 4975 12863 4981
rect 12989 4981 13001 4984
rect 13035 5012 13047 5015
rect 13078 5012 13084 5024
rect 13035 4984 13084 5012
rect 13035 4981 13047 4984
rect 12989 4975 13047 4981
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 13354 4972 13360 5024
rect 13412 4972 13418 5024
rect 16853 5015 16911 5021
rect 16853 4981 16865 5015
rect 16899 5012 16911 5015
rect 17034 5012 17040 5024
rect 16899 4984 17040 5012
rect 16899 4981 16911 4984
rect 16853 4975 16911 4981
rect 17034 4972 17040 4984
rect 17092 4972 17098 5024
rect 18616 5012 18644 5111
rect 18966 5108 18972 5120
rect 19024 5108 19030 5160
rect 22554 5108 22560 5160
rect 22612 5148 22618 5160
rect 22833 5151 22891 5157
rect 22833 5148 22845 5151
rect 22612 5120 22845 5148
rect 22612 5108 22618 5120
rect 22833 5117 22845 5120
rect 22879 5117 22891 5151
rect 22833 5111 22891 5117
rect 18874 5012 18880 5024
rect 18616 4984 18880 5012
rect 18874 4972 18880 4984
rect 18932 4972 18938 5024
rect 1104 4922 26312 4944
rect 1104 4870 4101 4922
rect 4153 4870 4165 4922
rect 4217 4870 4229 4922
rect 4281 4870 4293 4922
rect 4345 4870 4357 4922
rect 4409 4870 10403 4922
rect 10455 4870 10467 4922
rect 10519 4870 10531 4922
rect 10583 4870 10595 4922
rect 10647 4870 10659 4922
rect 10711 4870 16705 4922
rect 16757 4870 16769 4922
rect 16821 4870 16833 4922
rect 16885 4870 16897 4922
rect 16949 4870 16961 4922
rect 17013 4870 23007 4922
rect 23059 4870 23071 4922
rect 23123 4870 23135 4922
rect 23187 4870 23199 4922
rect 23251 4870 23263 4922
rect 23315 4870 26312 4922
rect 1104 4848 26312 4870
rect 5810 4768 5816 4820
rect 5868 4768 5874 4820
rect 6086 4768 6092 4820
rect 6144 4768 6150 4820
rect 7006 4768 7012 4820
rect 7064 4768 7070 4820
rect 8938 4768 8944 4820
rect 8996 4768 9002 4820
rect 9033 4811 9091 4817
rect 9033 4777 9045 4811
rect 9079 4808 9091 4811
rect 9122 4808 9128 4820
rect 9079 4780 9128 4808
rect 9079 4777 9091 4780
rect 9033 4771 9091 4777
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 9306 4768 9312 4820
rect 9364 4768 9370 4820
rect 9490 4768 9496 4820
rect 9548 4808 9554 4820
rect 10042 4808 10048 4820
rect 9548 4780 10048 4808
rect 9548 4768 9554 4780
rect 10042 4768 10048 4780
rect 10100 4768 10106 4820
rect 11330 4808 11336 4820
rect 10520 4780 11336 4808
rect 5626 4700 5632 4752
rect 5684 4740 5690 4752
rect 8956 4740 8984 4768
rect 5684 4712 8984 4740
rect 5684 4700 5690 4712
rect 6012 4623 6040 4712
rect 6270 4672 6276 4684
rect 6196 4644 6276 4672
rect 5997 4617 6055 4623
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4604 1823 4607
rect 3142 4604 3148 4616
rect 1811 4576 3148 4604
rect 1811 4573 1823 4576
rect 1765 4567 1823 4573
rect 3142 4564 3148 4576
rect 3200 4564 3206 4616
rect 5718 4564 5724 4616
rect 5776 4564 5782 4616
rect 5902 4564 5908 4616
rect 5960 4564 5966 4616
rect 5997 4583 6009 4617
rect 6043 4583 6055 4617
rect 6196 4613 6224 4644
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 8846 4632 8852 4684
rect 8904 4632 8910 4684
rect 9324 4681 9352 4768
rect 9309 4675 9367 4681
rect 9309 4641 9321 4675
rect 9355 4641 9367 4675
rect 9309 4635 9367 4641
rect 9766 4632 9772 4684
rect 9824 4632 9830 4684
rect 9953 4675 10011 4681
rect 9953 4641 9965 4675
rect 9999 4672 10011 4675
rect 10520 4672 10548 4780
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 11422 4768 11428 4820
rect 11480 4808 11486 4820
rect 11480 4780 12434 4808
rect 11480 4768 11486 4780
rect 12406 4740 12434 4780
rect 12894 4768 12900 4820
rect 12952 4808 12958 4820
rect 13538 4808 13544 4820
rect 12952 4780 13544 4808
rect 12952 4768 12958 4780
rect 13538 4768 13544 4780
rect 13596 4808 13602 4820
rect 13906 4808 13912 4820
rect 13596 4780 13912 4808
rect 13596 4768 13602 4780
rect 13906 4768 13912 4780
rect 13964 4768 13970 4820
rect 13998 4768 14004 4820
rect 14056 4808 14062 4820
rect 16577 4811 16635 4817
rect 16577 4808 16589 4811
rect 14056 4780 16589 4808
rect 14056 4768 14062 4780
rect 16577 4777 16589 4780
rect 16623 4777 16635 4811
rect 18782 4808 18788 4820
rect 16577 4771 16635 4777
rect 16868 4780 18788 4808
rect 16758 4740 16764 4752
rect 12406 4712 16764 4740
rect 16758 4700 16764 4712
rect 16816 4700 16822 4752
rect 9999 4644 10548 4672
rect 10597 4675 10655 4681
rect 9999 4641 10011 4644
rect 9953 4635 10011 4641
rect 10597 4641 10609 4675
rect 10643 4672 10655 4675
rect 10870 4672 10876 4684
rect 10643 4644 10876 4672
rect 10643 4641 10655 4644
rect 10597 4635 10655 4641
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 12897 4675 12955 4681
rect 12897 4641 12909 4675
rect 12943 4672 12955 4675
rect 12986 4672 12992 4684
rect 12943 4644 12992 4672
rect 12943 4641 12955 4644
rect 12897 4635 12955 4641
rect 12986 4632 12992 4644
rect 13044 4632 13050 4684
rect 13538 4632 13544 4684
rect 13596 4672 13602 4684
rect 13633 4675 13691 4681
rect 13633 4672 13645 4675
rect 13596 4644 13645 4672
rect 13596 4632 13602 4644
rect 13633 4641 13645 4644
rect 13679 4641 13691 4675
rect 16022 4672 16028 4684
rect 13633 4635 13691 4641
rect 15120 4644 16028 4672
rect 5997 4577 6055 4583
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4573 6975 4607
rect 6917 4567 6975 4573
rect 934 4496 940 4548
rect 992 4536 998 4548
rect 1397 4539 1455 4545
rect 1397 4536 1409 4539
rect 992 4508 1409 4536
rect 992 4496 998 4508
rect 1397 4505 1409 4508
rect 1443 4505 1455 4539
rect 6932 4536 6960 4567
rect 7098 4564 7104 4616
rect 7156 4564 7162 4616
rect 8864 4604 8892 4632
rect 9398 4604 9404 4616
rect 8864 4576 9404 4604
rect 9398 4564 9404 4576
rect 9456 4604 9462 4616
rect 9585 4607 9643 4613
rect 9585 4604 9597 4607
rect 9456 4576 9597 4604
rect 9456 4564 9462 4576
rect 9585 4573 9597 4576
rect 9631 4573 9643 4607
rect 9784 4604 9812 4632
rect 13360 4616 13412 4622
rect 12158 4604 12164 4616
rect 9784 4576 10180 4604
rect 12006 4576 12164 4604
rect 9585 4567 9643 4573
rect 10152 4536 10180 4576
rect 12158 4564 12164 4576
rect 12216 4564 12222 4616
rect 13360 4558 13412 4564
rect 10873 4539 10931 4545
rect 6932 4508 7696 4536
rect 10152 4508 10824 4536
rect 1397 4499 1455 4505
rect 7668 4480 7696 4508
rect 7650 4428 7656 4480
rect 7708 4428 7714 4480
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 10045 4471 10103 4477
rect 10045 4468 10057 4471
rect 9732 4440 10057 4468
rect 9732 4428 9738 4440
rect 10045 4437 10057 4440
rect 10091 4437 10103 4471
rect 10045 4431 10103 4437
rect 10410 4428 10416 4480
rect 10468 4428 10474 4480
rect 10796 4468 10824 4508
rect 10873 4505 10885 4539
rect 10919 4536 10931 4539
rect 11146 4536 11152 4548
rect 10919 4508 11152 4536
rect 10919 4505 10931 4508
rect 10873 4499 10931 4505
rect 11146 4496 11152 4508
rect 11204 4496 11210 4548
rect 12176 4508 13308 4536
rect 12176 4468 12204 4508
rect 10796 4440 12204 4468
rect 12342 4428 12348 4480
rect 12400 4428 12406 4480
rect 13280 4468 13308 4508
rect 15120 4468 15148 4644
rect 16022 4632 16028 4644
rect 16080 4672 16086 4684
rect 16117 4675 16175 4681
rect 16117 4672 16129 4675
rect 16080 4644 16129 4672
rect 16080 4632 16086 4644
rect 16117 4641 16129 4644
rect 16163 4672 16175 4675
rect 16868 4672 16896 4780
rect 18782 4768 18788 4780
rect 18840 4768 18846 4820
rect 18877 4811 18935 4817
rect 18877 4777 18889 4811
rect 18923 4808 18935 4811
rect 18966 4808 18972 4820
rect 18923 4780 18972 4808
rect 18923 4777 18935 4780
rect 18877 4771 18935 4777
rect 18966 4768 18972 4780
rect 19024 4768 19030 4820
rect 16163 4644 16896 4672
rect 16945 4675 17003 4681
rect 16163 4641 16175 4644
rect 16117 4635 16175 4641
rect 16945 4641 16957 4675
rect 16991 4672 17003 4675
rect 17034 4672 17040 4684
rect 16991 4644 17040 4672
rect 16991 4641 17003 4644
rect 16945 4635 17003 4641
rect 17034 4632 17040 4644
rect 17092 4632 17098 4684
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4604 16911 4607
rect 18046 4604 18052 4616
rect 16899 4576 18052 4604
rect 16899 4573 16911 4576
rect 16853 4567 16911 4573
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 19058 4564 19064 4616
rect 19116 4564 19122 4616
rect 16025 4539 16083 4545
rect 16025 4505 16037 4539
rect 16071 4536 16083 4539
rect 17770 4536 17776 4548
rect 16071 4508 17776 4536
rect 16071 4505 16083 4508
rect 16025 4499 16083 4505
rect 17770 4496 17776 4508
rect 17828 4496 17834 4548
rect 25593 4539 25651 4545
rect 25593 4536 25605 4539
rect 22066 4508 25605 4536
rect 13280 4440 15148 4468
rect 15194 4428 15200 4480
rect 15252 4468 15258 4480
rect 15565 4471 15623 4477
rect 15565 4468 15577 4471
rect 15252 4440 15577 4468
rect 15252 4428 15258 4440
rect 15565 4437 15577 4440
rect 15611 4437 15623 4471
rect 15565 4431 15623 4437
rect 15930 4428 15936 4480
rect 15988 4428 15994 4480
rect 16758 4428 16764 4480
rect 16816 4468 16822 4480
rect 22066 4468 22094 4508
rect 25593 4505 25605 4508
rect 25639 4505 25651 4539
rect 25593 4499 25651 4505
rect 16816 4440 22094 4468
rect 25869 4471 25927 4477
rect 16816 4428 16822 4440
rect 25869 4437 25881 4471
rect 25915 4468 25927 4471
rect 25958 4468 25964 4480
rect 25915 4440 25964 4468
rect 25915 4437 25927 4440
rect 25869 4431 25927 4437
rect 25958 4428 25964 4440
rect 26016 4428 26022 4480
rect 1104 4378 26472 4400
rect 1104 4326 7252 4378
rect 7304 4326 7316 4378
rect 7368 4326 7380 4378
rect 7432 4326 7444 4378
rect 7496 4326 7508 4378
rect 7560 4326 13554 4378
rect 13606 4326 13618 4378
rect 13670 4326 13682 4378
rect 13734 4326 13746 4378
rect 13798 4326 13810 4378
rect 13862 4326 19856 4378
rect 19908 4326 19920 4378
rect 19972 4326 19984 4378
rect 20036 4326 20048 4378
rect 20100 4326 20112 4378
rect 20164 4326 26158 4378
rect 26210 4326 26222 4378
rect 26274 4326 26286 4378
rect 26338 4326 26350 4378
rect 26402 4326 26414 4378
rect 26466 4326 26472 4378
rect 1104 4304 26472 4326
rect 6270 4224 6276 4276
rect 6328 4264 6334 4276
rect 6457 4267 6515 4273
rect 6457 4264 6469 4267
rect 6328 4236 6469 4264
rect 6328 4224 6334 4236
rect 6457 4233 6469 4236
rect 6503 4233 6515 4267
rect 6457 4227 6515 4233
rect 7650 4224 7656 4276
rect 7708 4264 7714 4276
rect 9493 4267 9551 4273
rect 9493 4264 9505 4267
rect 7708 4236 9505 4264
rect 7708 4224 7714 4236
rect 9493 4233 9505 4236
rect 9539 4233 9551 4267
rect 9493 4227 9551 4233
rect 9600 4236 10272 4264
rect 7098 4088 7104 4140
rect 7156 4088 7162 4140
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4128 7527 4131
rect 7668 4128 7696 4224
rect 9306 4196 9312 4208
rect 9154 4168 9312 4196
rect 9306 4156 9312 4168
rect 9364 4196 9370 4208
rect 9600 4196 9628 4236
rect 10244 4208 10272 4236
rect 10410 4224 10416 4276
rect 10468 4224 10474 4276
rect 10778 4224 10784 4276
rect 10836 4264 10842 4276
rect 10873 4267 10931 4273
rect 10873 4264 10885 4267
rect 10836 4236 10885 4264
rect 10836 4224 10842 4236
rect 10873 4233 10885 4236
rect 10919 4233 10931 4267
rect 10873 4227 10931 4233
rect 11146 4224 11152 4276
rect 11204 4264 11210 4276
rect 11517 4267 11575 4273
rect 11517 4264 11529 4267
rect 11204 4236 11529 4264
rect 11204 4224 11210 4236
rect 11517 4233 11529 4236
rect 11563 4233 11575 4267
rect 11517 4227 11575 4233
rect 13078 4224 13084 4276
rect 13136 4264 13142 4276
rect 13630 4264 13636 4276
rect 13136 4236 13636 4264
rect 13136 4224 13142 4236
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 9364 4168 9628 4196
rect 9364 4156 9370 4168
rect 9674 4156 9680 4208
rect 9732 4156 9738 4208
rect 10226 4156 10232 4208
rect 10284 4156 10290 4208
rect 7515 4100 7696 4128
rect 7515 4097 7527 4100
rect 7469 4091 7527 4097
rect 10042 4088 10048 4140
rect 10100 4088 10106 4140
rect 10321 4131 10379 4137
rect 10321 4097 10333 4131
rect 10367 4128 10379 4131
rect 10428 4128 10456 4224
rect 10965 4199 11023 4205
rect 10965 4165 10977 4199
rect 11011 4196 11023 4199
rect 11011 4168 11928 4196
rect 11011 4165 11023 4168
rect 10965 4159 11023 4165
rect 11701 4131 11759 4137
rect 11701 4128 11713 4131
rect 10367 4100 10456 4128
rect 11348 4100 11713 4128
rect 10367 4097 10379 4100
rect 10321 4091 10379 4097
rect 7653 4063 7711 4069
rect 7653 4029 7665 4063
rect 7699 4060 7711 4063
rect 7699 4032 7788 4060
rect 7699 4029 7711 4032
rect 7653 4023 7711 4029
rect 7760 3924 7788 4032
rect 7926 4020 7932 4072
rect 7984 4020 7990 4072
rect 10226 4060 10232 4072
rect 8956 4032 10232 4060
rect 8956 3924 8984 4032
rect 10226 4020 10232 4032
rect 10284 4020 10290 4072
rect 10689 4063 10747 4069
rect 10689 4029 10701 4063
rect 10735 4029 10747 4063
rect 10689 4023 10747 4029
rect 9398 3952 9404 4004
rect 9456 3992 9462 4004
rect 9456 3964 9720 3992
rect 9456 3952 9462 3964
rect 9692 3933 9720 3964
rect 7760 3896 8984 3924
rect 9677 3927 9735 3933
rect 9677 3893 9689 3927
rect 9723 3893 9735 3927
rect 9677 3887 9735 3893
rect 10134 3884 10140 3936
rect 10192 3884 10198 3936
rect 10704 3924 10732 4023
rect 11348 4001 11376 4100
rect 11701 4097 11713 4100
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 11900 4060 11928 4168
rect 13170 4156 13176 4208
rect 13228 4156 13234 4208
rect 15749 4199 15807 4205
rect 15749 4165 15761 4199
rect 15795 4196 15807 4199
rect 16114 4196 16120 4208
rect 15795 4168 16120 4196
rect 15795 4165 15807 4168
rect 15749 4159 15807 4165
rect 16114 4156 16120 4168
rect 16172 4156 16178 4208
rect 17037 4199 17095 4205
rect 17037 4165 17049 4199
rect 17083 4196 17095 4199
rect 17083 4168 18092 4196
rect 17083 4165 17095 4168
rect 17037 4159 17095 4165
rect 18064 4140 18092 4168
rect 21266 4156 21272 4208
rect 21324 4196 21330 4208
rect 21324 4168 22126 4196
rect 21324 4156 21330 4168
rect 11974 4088 11980 4140
rect 12032 4088 12038 4140
rect 12710 4088 12716 4140
rect 12768 4088 12774 4140
rect 13446 4088 13452 4140
rect 13504 4128 13510 4140
rect 13725 4131 13783 4137
rect 13725 4128 13737 4131
rect 13504 4100 13737 4128
rect 13504 4088 13510 4100
rect 13725 4097 13737 4100
rect 13771 4097 13783 4131
rect 13725 4091 13783 4097
rect 15197 4131 15255 4137
rect 15197 4097 15209 4131
rect 15243 4128 15255 4131
rect 15841 4131 15899 4137
rect 15243 4100 15424 4128
rect 15243 4097 15255 4100
rect 15197 4091 15255 4097
rect 12342 4060 12348 4072
rect 11900 4032 12348 4060
rect 12342 4020 12348 4032
rect 12400 4020 12406 4072
rect 13817 4063 13875 4069
rect 13817 4029 13829 4063
rect 13863 4029 13875 4063
rect 13817 4023 13875 4029
rect 11333 3995 11391 4001
rect 11333 3961 11345 3995
rect 11379 3961 11391 3995
rect 11882 3992 11888 4004
rect 11333 3955 11391 3961
rect 11440 3964 11888 3992
rect 11440 3924 11468 3964
rect 11882 3952 11888 3964
rect 11940 3992 11946 4004
rect 13832 3992 13860 4023
rect 15396 4001 15424 4100
rect 15841 4097 15853 4131
rect 15887 4128 15899 4131
rect 17126 4128 17132 4140
rect 15887 4100 17132 4128
rect 15887 4097 15899 4100
rect 15841 4091 15899 4097
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 17770 4088 17776 4140
rect 17828 4088 17834 4140
rect 17862 4088 17868 4140
rect 17920 4088 17926 4140
rect 18046 4088 18052 4140
rect 18104 4088 18110 4140
rect 23569 4131 23627 4137
rect 23569 4097 23581 4131
rect 23615 4128 23627 4131
rect 23658 4128 23664 4140
rect 23615 4100 23664 4128
rect 23615 4097 23627 4100
rect 23569 4091 23627 4097
rect 23658 4088 23664 4100
rect 23716 4088 23722 4140
rect 16022 4020 16028 4072
rect 16080 4020 16086 4072
rect 17221 4063 17279 4069
rect 17221 4060 17233 4063
rect 16316 4032 17233 4060
rect 15381 3995 15439 4001
rect 11940 3964 15332 3992
rect 11940 3952 11946 3964
rect 10704 3896 11468 3924
rect 11790 3884 11796 3936
rect 11848 3884 11854 3936
rect 13262 3884 13268 3936
rect 13320 3884 13326 3936
rect 15010 3884 15016 3936
rect 15068 3884 15074 3936
rect 15304 3924 15332 3964
rect 15381 3961 15393 3995
rect 15427 3961 15439 3995
rect 15381 3955 15439 3961
rect 16316 3924 16344 4032
rect 17221 4029 17233 4032
rect 17267 4060 17279 4063
rect 17589 4063 17647 4069
rect 17589 4060 17601 4063
rect 17267 4032 17601 4060
rect 17267 4029 17279 4032
rect 17221 4023 17279 4029
rect 17589 4029 17601 4032
rect 17635 4060 17647 4063
rect 18506 4060 18512 4072
rect 17635 4032 18512 4060
rect 17635 4029 17647 4032
rect 17589 4023 17647 4029
rect 18506 4020 18512 4032
rect 18564 4020 18570 4072
rect 21821 4063 21879 4069
rect 21821 4029 21833 4063
rect 21867 4060 21879 4063
rect 22554 4060 22560 4072
rect 21867 4032 22560 4060
rect 21867 4029 21879 4032
rect 21821 4023 21879 4029
rect 22554 4020 22560 4032
rect 22612 4020 22618 4072
rect 22830 4020 22836 4072
rect 22888 4060 22894 4072
rect 23293 4063 23351 4069
rect 23293 4060 23305 4063
rect 22888 4032 23305 4060
rect 22888 4020 22894 4032
rect 23293 4029 23305 4032
rect 23339 4029 23351 4063
rect 23293 4023 23351 4029
rect 15304 3896 16344 3924
rect 16390 3884 16396 3936
rect 16448 3924 16454 3936
rect 16669 3927 16727 3933
rect 16669 3924 16681 3927
rect 16448 3896 16681 3924
rect 16448 3884 16454 3896
rect 16669 3893 16681 3896
rect 16715 3893 16727 3927
rect 16669 3887 16727 3893
rect 18230 3884 18236 3936
rect 18288 3884 18294 3936
rect 1104 3834 26312 3856
rect 1104 3782 4101 3834
rect 4153 3782 4165 3834
rect 4217 3782 4229 3834
rect 4281 3782 4293 3834
rect 4345 3782 4357 3834
rect 4409 3782 10403 3834
rect 10455 3782 10467 3834
rect 10519 3782 10531 3834
rect 10583 3782 10595 3834
rect 10647 3782 10659 3834
rect 10711 3782 16705 3834
rect 16757 3782 16769 3834
rect 16821 3782 16833 3834
rect 16885 3782 16897 3834
rect 16949 3782 16961 3834
rect 17013 3782 23007 3834
rect 23059 3782 23071 3834
rect 23123 3782 23135 3834
rect 23187 3782 23199 3834
rect 23251 3782 23263 3834
rect 23315 3782 26312 3834
rect 1104 3760 26312 3782
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 7377 3723 7435 3729
rect 7377 3720 7389 3723
rect 7156 3692 7389 3720
rect 7156 3680 7162 3692
rect 7377 3689 7389 3692
rect 7423 3689 7435 3723
rect 7377 3683 7435 3689
rect 1394 3544 1400 3596
rect 1452 3584 1458 3596
rect 5629 3587 5687 3593
rect 5629 3584 5641 3587
rect 1452 3556 5641 3584
rect 1452 3544 1458 3556
rect 5629 3553 5641 3556
rect 5675 3553 5687 3587
rect 5629 3547 5687 3553
rect 7392 3516 7420 3683
rect 7926 3680 7932 3732
rect 7984 3720 7990 3732
rect 8297 3723 8355 3729
rect 8297 3720 8309 3723
rect 7984 3692 8309 3720
rect 7984 3680 7990 3692
rect 8297 3689 8309 3692
rect 8343 3689 8355 3723
rect 8297 3683 8355 3689
rect 10492 3723 10550 3729
rect 10492 3689 10504 3723
rect 10538 3720 10550 3723
rect 11790 3720 11796 3732
rect 10538 3692 11796 3720
rect 10538 3689 10550 3692
rect 10492 3683 10550 3689
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 11977 3723 12035 3729
rect 11977 3689 11989 3723
rect 12023 3720 12035 3723
rect 12434 3720 12440 3732
rect 12023 3692 12440 3720
rect 12023 3689 12035 3692
rect 11977 3683 12035 3689
rect 12434 3680 12440 3692
rect 12492 3720 12498 3732
rect 12986 3720 12992 3732
rect 12492 3692 12992 3720
rect 12492 3680 12498 3692
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 13446 3680 13452 3732
rect 13504 3680 13510 3732
rect 13630 3680 13636 3732
rect 13688 3720 13694 3732
rect 13817 3723 13875 3729
rect 13817 3720 13829 3723
rect 13688 3692 13829 3720
rect 13688 3680 13694 3692
rect 13817 3689 13829 3692
rect 13863 3689 13875 3723
rect 15194 3720 15200 3732
rect 13817 3683 13875 3689
rect 14200 3692 15200 3720
rect 11514 3612 11520 3664
rect 11572 3652 11578 3664
rect 11572 3624 12204 3652
rect 11572 3612 11578 3624
rect 7929 3587 7987 3593
rect 7929 3553 7941 3587
rect 7975 3584 7987 3587
rect 8018 3584 8024 3596
rect 7975 3556 8024 3584
rect 7975 3553 7987 3556
rect 7929 3547 7987 3553
rect 8018 3544 8024 3556
rect 8076 3544 8082 3596
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3584 8171 3587
rect 9493 3587 9551 3593
rect 9493 3584 9505 3587
rect 8159 3556 9505 3584
rect 8159 3553 8171 3556
rect 8113 3547 8171 3553
rect 9493 3553 9505 3556
rect 9539 3584 9551 3587
rect 9766 3584 9772 3596
rect 9539 3556 9772 3584
rect 9539 3553 9551 3556
rect 9493 3547 9551 3553
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 10226 3544 10232 3596
rect 10284 3584 10290 3596
rect 10870 3584 10876 3596
rect 10284 3556 10876 3584
rect 10284 3544 10290 3556
rect 10870 3544 10876 3556
rect 10928 3584 10934 3596
rect 12069 3587 12127 3593
rect 12069 3584 12081 3587
rect 10928 3556 12081 3584
rect 10928 3544 10934 3556
rect 12069 3553 12081 3556
rect 12115 3553 12127 3587
rect 12176 3584 12204 3624
rect 13464 3584 13492 3680
rect 12176 3556 13492 3584
rect 12069 3547 12127 3553
rect 7837 3519 7895 3525
rect 7837 3516 7849 3519
rect 7392 3488 7849 3516
rect 7837 3485 7849 3488
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3516 8539 3519
rect 9309 3519 9367 3525
rect 8527 3488 8984 3516
rect 8527 3485 8539 3488
rect 8481 3479 8539 3485
rect 5902 3408 5908 3460
rect 5960 3408 5966 3460
rect 6012 3420 6394 3448
rect 3418 3340 3424 3392
rect 3476 3380 3482 3392
rect 6012 3380 6040 3420
rect 3476 3352 6040 3380
rect 7469 3383 7527 3389
rect 3476 3340 3482 3352
rect 7469 3349 7481 3383
rect 7515 3380 7527 3383
rect 7650 3380 7656 3392
rect 7515 3352 7656 3380
rect 7515 3349 7527 3352
rect 7469 3343 7527 3349
rect 7650 3340 7656 3352
rect 7708 3340 7714 3392
rect 8956 3389 8984 3488
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9398 3516 9404 3528
rect 9355 3488 9404 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 14200 3525 14228 3692
rect 15194 3680 15200 3692
rect 15252 3680 15258 3732
rect 15930 3680 15936 3732
rect 15988 3720 15994 3732
rect 16209 3723 16267 3729
rect 16209 3720 16221 3723
rect 15988 3692 16221 3720
rect 15988 3680 15994 3692
rect 16209 3689 16221 3692
rect 16255 3689 16267 3723
rect 16209 3683 16267 3689
rect 18046 3680 18052 3732
rect 18104 3680 18110 3732
rect 22465 3723 22523 3729
rect 22465 3689 22477 3723
rect 22511 3720 22523 3723
rect 22830 3720 22836 3732
rect 22511 3692 22836 3720
rect 22511 3689 22523 3692
rect 22465 3683 22523 3689
rect 22830 3680 22836 3692
rect 22888 3680 22894 3732
rect 16301 3587 16359 3593
rect 16301 3584 16313 3587
rect 14476 3556 16313 3584
rect 14185 3519 14243 3525
rect 14185 3485 14197 3519
rect 14231 3485 14243 3519
rect 14185 3479 14243 3485
rect 14366 3476 14372 3528
rect 14424 3516 14430 3528
rect 14476 3525 14504 3556
rect 16301 3553 16313 3556
rect 16347 3584 16359 3587
rect 18874 3584 18880 3596
rect 16347 3556 18880 3584
rect 16347 3553 16359 3556
rect 16301 3547 16359 3553
rect 18874 3544 18880 3556
rect 18932 3584 18938 3596
rect 19705 3587 19763 3593
rect 19705 3584 19717 3587
rect 18932 3556 19717 3584
rect 18932 3544 18938 3556
rect 19705 3553 19717 3556
rect 19751 3553 19763 3587
rect 19705 3547 19763 3553
rect 21453 3587 21511 3593
rect 21453 3553 21465 3587
rect 21499 3584 21511 3587
rect 21821 3587 21879 3593
rect 21821 3584 21833 3587
rect 21499 3556 21833 3584
rect 21499 3553 21511 3556
rect 21453 3547 21511 3553
rect 21821 3553 21833 3556
rect 21867 3553 21879 3587
rect 21821 3547 21879 3553
rect 14461 3519 14519 3525
rect 14461 3516 14473 3519
rect 14424 3488 14473 3516
rect 14424 3476 14430 3488
rect 14461 3485 14473 3488
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 18141 3519 18199 3525
rect 18141 3485 18153 3519
rect 18187 3516 18199 3519
rect 18230 3516 18236 3528
rect 18187 3488 18236 3516
rect 18187 3485 18199 3488
rect 18141 3479 18199 3485
rect 18230 3476 18236 3488
rect 18288 3476 18294 3528
rect 11730 3420 11836 3448
rect 8941 3383 8999 3389
rect 8941 3349 8953 3383
rect 8987 3349 8999 3383
rect 8941 3343 8999 3349
rect 9401 3383 9459 3389
rect 9401 3349 9413 3383
rect 9447 3380 9459 3383
rect 11514 3380 11520 3392
rect 9447 3352 11520 3380
rect 9447 3349 9459 3352
rect 9401 3343 9459 3349
rect 11514 3340 11520 3352
rect 11572 3340 11578 3392
rect 11808 3380 11836 3420
rect 12342 3408 12348 3460
rect 12400 3408 12406 3460
rect 14737 3451 14795 3457
rect 12544 3420 12834 3448
rect 12158 3380 12164 3392
rect 11808 3352 12164 3380
rect 12158 3340 12164 3352
rect 12216 3380 12222 3392
rect 12544 3380 12572 3420
rect 14737 3417 14749 3451
rect 14783 3417 14795 3451
rect 15194 3448 15200 3460
rect 14737 3411 14795 3417
rect 15120 3420 15200 3448
rect 12216 3352 12572 3380
rect 14369 3383 14427 3389
rect 12216 3340 12222 3352
rect 14369 3349 14381 3383
rect 14415 3380 14427 3383
rect 14752 3380 14780 3411
rect 14415 3352 14780 3380
rect 15120 3380 15148 3420
rect 15194 3408 15200 3420
rect 15252 3408 15258 3460
rect 16574 3408 16580 3460
rect 16632 3408 16638 3460
rect 17034 3448 17040 3460
rect 16960 3420 17040 3448
rect 16960 3380 16988 3420
rect 17034 3408 17040 3420
rect 17092 3408 17098 3460
rect 19981 3451 20039 3457
rect 19981 3417 19993 3451
rect 20027 3448 20039 3451
rect 20254 3448 20260 3460
rect 20027 3420 20260 3448
rect 20027 3417 20039 3420
rect 19981 3411 20039 3417
rect 20254 3408 20260 3420
rect 20312 3408 20318 3460
rect 21266 3448 21272 3460
rect 21206 3420 21272 3448
rect 21266 3408 21272 3420
rect 21324 3408 21330 3460
rect 15120 3352 16988 3380
rect 14415 3349 14427 3352
rect 14369 3343 14427 3349
rect 18322 3340 18328 3392
rect 18380 3340 18386 3392
rect 1104 3290 26472 3312
rect 1104 3238 7252 3290
rect 7304 3238 7316 3290
rect 7368 3238 7380 3290
rect 7432 3238 7444 3290
rect 7496 3238 7508 3290
rect 7560 3238 13554 3290
rect 13606 3238 13618 3290
rect 13670 3238 13682 3290
rect 13734 3238 13746 3290
rect 13798 3238 13810 3290
rect 13862 3238 19856 3290
rect 19908 3238 19920 3290
rect 19972 3238 19984 3290
rect 20036 3238 20048 3290
rect 20100 3238 20112 3290
rect 20164 3238 26158 3290
rect 26210 3238 26222 3290
rect 26274 3238 26286 3290
rect 26338 3238 26350 3290
rect 26402 3238 26414 3290
rect 26466 3238 26472 3290
rect 1104 3216 26472 3238
rect 5902 3136 5908 3188
rect 5960 3176 5966 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 5960 3148 6561 3176
rect 5960 3136 5966 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 7650 3136 7656 3188
rect 7708 3136 7714 3188
rect 8389 3179 8447 3185
rect 8389 3145 8401 3179
rect 8435 3176 8447 3179
rect 9674 3176 9680 3188
rect 8435 3148 9680 3176
rect 8435 3145 8447 3148
rect 8389 3139 8447 3145
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 10134 3176 10140 3188
rect 9876 3148 10140 3176
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3040 6791 3043
rect 7668 3040 7696 3136
rect 9306 3068 9312 3120
rect 9364 3068 9370 3120
rect 9876 3117 9904 3148
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 11974 3136 11980 3188
rect 12032 3176 12038 3188
rect 12253 3179 12311 3185
rect 12253 3176 12265 3179
rect 12032 3148 12265 3176
rect 12032 3136 12038 3148
rect 12253 3145 12265 3148
rect 12299 3145 12311 3179
rect 12253 3139 12311 3145
rect 12342 3136 12348 3188
rect 12400 3176 12406 3188
rect 12529 3179 12587 3185
rect 12529 3176 12541 3179
rect 12400 3148 12541 3176
rect 12400 3136 12406 3148
rect 12529 3145 12541 3148
rect 12575 3145 12587 3179
rect 12529 3139 12587 3145
rect 13262 3136 13268 3188
rect 13320 3136 13326 3188
rect 15010 3136 15016 3188
rect 15068 3136 15074 3188
rect 16114 3136 16120 3188
rect 16172 3136 16178 3188
rect 16390 3136 16396 3188
rect 16448 3136 16454 3188
rect 16485 3179 16543 3185
rect 16485 3145 16497 3179
rect 16531 3176 16543 3179
rect 16574 3176 16580 3188
rect 16531 3148 16580 3176
rect 16531 3145 16543 3148
rect 16485 3139 16543 3145
rect 16574 3136 16580 3148
rect 16632 3136 16638 3188
rect 17129 3179 17187 3185
rect 17129 3145 17141 3179
rect 17175 3176 17187 3179
rect 17862 3176 17868 3188
rect 17175 3148 17868 3176
rect 17175 3145 17187 3148
rect 17129 3139 17187 3145
rect 17862 3136 17868 3148
rect 17920 3136 17926 3188
rect 18322 3136 18328 3188
rect 18380 3136 18386 3188
rect 9861 3111 9919 3117
rect 9861 3077 9873 3111
rect 9907 3077 9919 3111
rect 11793 3111 11851 3117
rect 11793 3108 11805 3111
rect 9861 3071 9919 3077
rect 10336 3080 11805 3108
rect 6779 3012 7696 3040
rect 10137 3043 10195 3049
rect 6779 3009 6791 3012
rect 6733 3003 6791 3009
rect 10137 3009 10149 3043
rect 10183 3040 10195 3043
rect 10226 3040 10232 3052
rect 10183 3012 10232 3040
rect 10183 3009 10195 3012
rect 10137 3003 10195 3009
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 8018 2932 8024 2984
rect 8076 2972 8082 2984
rect 10336 2972 10364 3080
rect 11793 3077 11805 3080
rect 11839 3077 11851 3111
rect 11793 3071 11851 3077
rect 11885 3111 11943 3117
rect 11885 3077 11897 3111
rect 11931 3108 11943 3111
rect 12434 3108 12440 3120
rect 11931 3080 12440 3108
rect 11931 3077 11943 3080
rect 11885 3071 11943 3077
rect 12434 3068 12440 3080
rect 12492 3068 12498 3120
rect 12713 3043 12771 3049
rect 11716 3012 11928 3040
rect 11716 2981 11744 3012
rect 11900 2984 11928 3012
rect 12713 3009 12725 3043
rect 12759 3040 12771 3043
rect 13280 3040 13308 3136
rect 14645 3111 14703 3117
rect 14645 3077 14657 3111
rect 14691 3108 14703 3111
rect 15028 3108 15056 3136
rect 14691 3080 15056 3108
rect 14691 3077 14703 3080
rect 14645 3071 14703 3077
rect 15286 3068 15292 3120
rect 15344 3068 15350 3120
rect 12759 3012 13308 3040
rect 12759 3009 12771 3012
rect 12713 3003 12771 3009
rect 14366 3000 14372 3052
rect 14424 3000 14430 3052
rect 16301 3043 16359 3049
rect 16301 3009 16313 3043
rect 16347 3040 16359 3043
rect 16408 3040 16436 3136
rect 17034 3068 17040 3120
rect 17092 3108 17098 3120
rect 18340 3108 18368 3136
rect 18601 3111 18659 3117
rect 18601 3108 18613 3111
rect 17092 3080 17434 3108
rect 18340 3080 18613 3108
rect 17092 3068 17098 3080
rect 18601 3077 18613 3080
rect 18647 3077 18659 3111
rect 18601 3071 18659 3077
rect 16347 3012 16436 3040
rect 16347 3009 16359 3012
rect 16301 3003 16359 3009
rect 8076 2944 10364 2972
rect 11701 2975 11759 2981
rect 8076 2932 8082 2944
rect 11701 2941 11713 2975
rect 11747 2941 11759 2975
rect 11701 2935 11759 2941
rect 11882 2932 11888 2984
rect 11940 2932 11946 2984
rect 18874 2932 18880 2984
rect 18932 2932 18938 2984
rect 1104 2746 26312 2768
rect 1104 2694 4101 2746
rect 4153 2694 4165 2746
rect 4217 2694 4229 2746
rect 4281 2694 4293 2746
rect 4345 2694 4357 2746
rect 4409 2694 10403 2746
rect 10455 2694 10467 2746
rect 10519 2694 10531 2746
rect 10583 2694 10595 2746
rect 10647 2694 10659 2746
rect 10711 2694 16705 2746
rect 16757 2694 16769 2746
rect 16821 2694 16833 2746
rect 16885 2694 16897 2746
rect 16949 2694 16961 2746
rect 17013 2694 23007 2746
rect 23059 2694 23071 2746
rect 23123 2694 23135 2746
rect 23187 2694 23199 2746
rect 23251 2694 23263 2746
rect 23315 2694 26312 2746
rect 1104 2672 26312 2694
rect 20073 2635 20131 2641
rect 20073 2601 20085 2635
rect 20119 2632 20131 2635
rect 20254 2632 20260 2644
rect 20119 2604 20260 2632
rect 20119 2601 20131 2604
rect 20073 2595 20131 2601
rect 20254 2592 20260 2604
rect 20312 2592 20318 2644
rect 25130 2592 25136 2644
rect 25188 2632 25194 2644
rect 25777 2635 25835 2641
rect 25777 2632 25789 2635
rect 25188 2604 25789 2632
rect 25188 2592 25194 2604
rect 25777 2601 25789 2604
rect 25823 2601 25835 2635
rect 25777 2595 25835 2601
rect 3510 2456 3516 2508
rect 3568 2496 3574 2508
rect 3568 2468 6914 2496
rect 3568 2456 3574 2468
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2428 1823 2431
rect 2222 2428 2228 2440
rect 1811 2400 2228 2428
rect 1811 2397 1823 2400
rect 1765 2391 1823 2397
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 4890 2428 4896 2440
rect 4387 2400 4896 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 6886 2428 6914 2468
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 6886 2400 7941 2428
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 14182 2428 14188 2440
rect 12115 2400 14188 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 15930 2388 15936 2440
rect 15988 2388 15994 2440
rect 20254 2388 20260 2440
rect 20312 2388 20318 2440
rect 25961 2431 26019 2437
rect 25961 2428 25973 2431
rect 24780 2400 25973 2428
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 72 2332 1409 2360
rect 72 2320 78 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 3970 2320 3976 2372
rect 4028 2320 4034 2372
rect 11698 2320 11704 2372
rect 11756 2320 11762 2372
rect 15562 2320 15568 2372
rect 15620 2320 15626 2372
rect 16390 2320 16396 2372
rect 16448 2360 16454 2372
rect 24489 2363 24547 2369
rect 24489 2360 24501 2363
rect 16448 2332 24501 2360
rect 16448 2320 16454 2332
rect 24489 2329 24501 2332
rect 24535 2329 24547 2363
rect 24489 2323 24547 2329
rect 24780 2304 24808 2400
rect 25961 2397 25973 2400
rect 26007 2397 26019 2431
rect 25961 2391 26019 2397
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7800 2264 8033 2292
rect 7800 2252 7806 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 23842 2252 23848 2304
rect 23900 2292 23906 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 23900 2264 24593 2292
rect 23900 2252 23906 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 24762 2252 24768 2304
rect 24820 2252 24826 2304
rect 1104 2202 26472 2224
rect 1104 2150 7252 2202
rect 7304 2150 7316 2202
rect 7368 2150 7380 2202
rect 7432 2150 7444 2202
rect 7496 2150 7508 2202
rect 7560 2150 13554 2202
rect 13606 2150 13618 2202
rect 13670 2150 13682 2202
rect 13734 2150 13746 2202
rect 13798 2150 13810 2202
rect 13862 2150 19856 2202
rect 19908 2150 19920 2202
rect 19972 2150 19984 2202
rect 20036 2150 20048 2202
rect 20100 2150 20112 2202
rect 20164 2150 26158 2202
rect 26210 2150 26222 2202
rect 26274 2150 26286 2202
rect 26338 2150 26350 2202
rect 26402 2150 26414 2202
rect 26466 2150 26472 2202
rect 1104 2128 26472 2150
<< via1 >>
rect 7252 27174 7304 27226
rect 7316 27174 7368 27226
rect 7380 27174 7432 27226
rect 7444 27174 7496 27226
rect 7508 27174 7560 27226
rect 13554 27174 13606 27226
rect 13618 27174 13670 27226
rect 13682 27174 13734 27226
rect 13746 27174 13798 27226
rect 13810 27174 13862 27226
rect 19856 27174 19908 27226
rect 19920 27174 19972 27226
rect 19984 27174 20036 27226
rect 20048 27174 20100 27226
rect 20112 27174 20164 27226
rect 26158 27174 26210 27226
rect 26222 27174 26274 27226
rect 26286 27174 26338 27226
rect 26350 27174 26402 27226
rect 26414 27174 26466 27226
rect 2780 27072 2832 27124
rect 3240 27072 3292 27124
rect 7104 27072 7156 27124
rect 11612 27072 11664 27124
rect 1768 26979 1820 26988
rect 1768 26945 1777 26979
rect 1777 26945 1811 26979
rect 1811 26945 1820 26979
rect 1768 26936 1820 26945
rect 5080 26936 5132 26988
rect 10968 26979 11020 26988
rect 10968 26945 10977 26979
rect 10977 26945 11011 26979
rect 11011 26945 11020 26979
rect 10968 26936 11020 26945
rect 11336 26936 11388 26988
rect 15200 27072 15252 27124
rect 15752 27115 15804 27124
rect 15752 27081 15761 27115
rect 15761 27081 15795 27115
rect 15795 27081 15804 27115
rect 15752 27072 15804 27081
rect 19340 27072 19392 27124
rect 23480 27072 23532 27124
rect 13452 27004 13504 27056
rect 14004 26936 14056 26988
rect 15660 26979 15712 26988
rect 15660 26945 15669 26979
rect 15669 26945 15703 26979
rect 15703 26945 15712 26979
rect 15660 26936 15712 26945
rect 17132 26936 17184 26988
rect 20996 26979 21048 26988
rect 14924 26868 14976 26920
rect 15384 26868 15436 26920
rect 20996 26945 21005 26979
rect 21005 26945 21039 26979
rect 21039 26945 21048 26979
rect 20996 26936 21048 26945
rect 20720 26911 20772 26920
rect 20720 26877 20729 26911
rect 20729 26877 20763 26911
rect 20763 26877 20772 26911
rect 20720 26868 20772 26877
rect 7196 26775 7248 26784
rect 7196 26741 7205 26775
rect 7205 26741 7239 26775
rect 7239 26741 7248 26775
rect 7196 26732 7248 26741
rect 9772 26732 9824 26784
rect 10784 26732 10836 26784
rect 11428 26732 11480 26784
rect 12256 26732 12308 26784
rect 12440 26732 12492 26784
rect 17040 26732 17092 26784
rect 19616 26775 19668 26784
rect 19616 26741 19625 26775
rect 19625 26741 19659 26775
rect 19659 26741 19668 26775
rect 19616 26732 19668 26741
rect 22468 26732 22520 26784
rect 4101 26630 4153 26682
rect 4165 26630 4217 26682
rect 4229 26630 4281 26682
rect 4293 26630 4345 26682
rect 4357 26630 4409 26682
rect 10403 26630 10455 26682
rect 10467 26630 10519 26682
rect 10531 26630 10583 26682
rect 10595 26630 10647 26682
rect 10659 26630 10711 26682
rect 16705 26630 16757 26682
rect 16769 26630 16821 26682
rect 16833 26630 16885 26682
rect 16897 26630 16949 26682
rect 16961 26630 17013 26682
rect 23007 26630 23059 26682
rect 23071 26630 23123 26682
rect 23135 26630 23187 26682
rect 23199 26630 23251 26682
rect 23263 26630 23315 26682
rect 7196 26528 7248 26580
rect 10784 26528 10836 26580
rect 14924 26528 14976 26580
rect 8484 26324 8536 26376
rect 11336 26367 11388 26376
rect 11336 26333 11345 26367
rect 11345 26333 11379 26367
rect 11379 26333 11388 26367
rect 11336 26324 11388 26333
rect 11796 26324 11848 26376
rect 15292 26460 15344 26512
rect 15476 26460 15528 26512
rect 14556 26392 14608 26444
rect 4988 26188 5040 26240
rect 7656 26256 7708 26308
rect 8852 26256 8904 26308
rect 13912 26324 13964 26376
rect 8024 26188 8076 26240
rect 8208 26188 8260 26240
rect 15200 26367 15252 26376
rect 15200 26333 15209 26367
rect 15209 26333 15243 26367
rect 15243 26333 15252 26367
rect 15200 26324 15252 26333
rect 20904 26392 20956 26444
rect 17316 26324 17368 26376
rect 17500 26367 17552 26376
rect 17500 26333 17509 26367
rect 17509 26333 17543 26367
rect 17543 26333 17552 26367
rect 17500 26324 17552 26333
rect 17684 26324 17736 26376
rect 18420 26324 18472 26376
rect 22836 26392 22888 26444
rect 9956 26188 10008 26240
rect 11888 26231 11940 26240
rect 11888 26197 11897 26231
rect 11897 26197 11931 26231
rect 11931 26197 11940 26231
rect 11888 26188 11940 26197
rect 12532 26188 12584 26240
rect 13452 26188 13504 26240
rect 14556 26188 14608 26240
rect 14832 26188 14884 26240
rect 18512 26256 18564 26308
rect 15568 26231 15620 26240
rect 15568 26197 15577 26231
rect 15577 26197 15611 26231
rect 15611 26197 15620 26231
rect 15568 26188 15620 26197
rect 17408 26188 17460 26240
rect 22100 26256 22152 26308
rect 22744 26188 22796 26240
rect 7252 26086 7304 26138
rect 7316 26086 7368 26138
rect 7380 26086 7432 26138
rect 7444 26086 7496 26138
rect 7508 26086 7560 26138
rect 13554 26086 13606 26138
rect 13618 26086 13670 26138
rect 13682 26086 13734 26138
rect 13746 26086 13798 26138
rect 13810 26086 13862 26138
rect 19856 26086 19908 26138
rect 19920 26086 19972 26138
rect 19984 26086 20036 26138
rect 20048 26086 20100 26138
rect 20112 26086 20164 26138
rect 26158 26086 26210 26138
rect 26222 26086 26274 26138
rect 26286 26086 26338 26138
rect 26350 26086 26402 26138
rect 26414 26086 26466 26138
rect 11336 25984 11388 26036
rect 7472 25916 7524 25968
rect 8024 25916 8076 25968
rect 5908 25780 5960 25832
rect 6920 25780 6972 25832
rect 8484 25823 8536 25832
rect 8484 25789 8493 25823
rect 8493 25789 8527 25823
rect 8527 25789 8536 25823
rect 8484 25780 8536 25789
rect 8760 25823 8812 25832
rect 8760 25789 8769 25823
rect 8769 25789 8803 25823
rect 8803 25789 8812 25823
rect 8760 25780 8812 25789
rect 11336 25891 11388 25900
rect 11336 25857 11345 25891
rect 11345 25857 11379 25891
rect 11379 25857 11388 25891
rect 11336 25848 11388 25857
rect 12348 25916 12400 25968
rect 12532 25916 12584 25968
rect 13912 26027 13964 26036
rect 13912 25993 13921 26027
rect 13921 25993 13955 26027
rect 13955 25993 13964 26027
rect 13912 25984 13964 25993
rect 14004 26027 14056 26036
rect 14004 25993 14013 26027
rect 14013 25993 14047 26027
rect 14047 25993 14056 26027
rect 14004 25984 14056 25993
rect 15384 25984 15436 26036
rect 14648 25916 14700 25968
rect 17040 25916 17092 25968
rect 18236 25916 18288 25968
rect 18512 25916 18564 25968
rect 22468 25916 22520 25968
rect 22744 25916 22796 25968
rect 14464 25848 14516 25900
rect 20812 25848 20864 25900
rect 10876 25823 10928 25832
rect 10876 25789 10885 25823
rect 10885 25789 10919 25823
rect 10919 25789 10928 25823
rect 10876 25780 10928 25789
rect 11980 25780 12032 25832
rect 14556 25823 14608 25832
rect 14556 25789 14565 25823
rect 14565 25789 14599 25823
rect 14599 25789 14608 25823
rect 14556 25780 14608 25789
rect 15568 25780 15620 25832
rect 16580 25780 16632 25832
rect 18420 25823 18472 25832
rect 18420 25789 18429 25823
rect 18429 25789 18463 25823
rect 18463 25789 18472 25823
rect 18420 25780 18472 25789
rect 5356 25644 5408 25696
rect 7472 25644 7524 25696
rect 10784 25644 10836 25696
rect 12164 25644 12216 25696
rect 12624 25644 12676 25696
rect 17684 25644 17736 25696
rect 20628 25823 20680 25832
rect 20628 25789 20637 25823
rect 20637 25789 20671 25823
rect 20671 25789 20680 25823
rect 20628 25780 20680 25789
rect 20904 25780 20956 25832
rect 19248 25644 19300 25696
rect 20260 25687 20312 25696
rect 20260 25653 20269 25687
rect 20269 25653 20303 25687
rect 20303 25653 20312 25687
rect 20260 25644 20312 25653
rect 21180 25687 21232 25696
rect 21180 25653 21189 25687
rect 21189 25653 21223 25687
rect 21223 25653 21232 25687
rect 21180 25644 21232 25653
rect 21456 25687 21508 25696
rect 21456 25653 21465 25687
rect 21465 25653 21499 25687
rect 21499 25653 21508 25687
rect 21456 25644 21508 25653
rect 23664 25687 23716 25696
rect 23664 25653 23673 25687
rect 23673 25653 23707 25687
rect 23707 25653 23716 25687
rect 23664 25644 23716 25653
rect 4101 25542 4153 25594
rect 4165 25542 4217 25594
rect 4229 25542 4281 25594
rect 4293 25542 4345 25594
rect 4357 25542 4409 25594
rect 10403 25542 10455 25594
rect 10467 25542 10519 25594
rect 10531 25542 10583 25594
rect 10595 25542 10647 25594
rect 10659 25542 10711 25594
rect 16705 25542 16757 25594
rect 16769 25542 16821 25594
rect 16833 25542 16885 25594
rect 16897 25542 16949 25594
rect 16961 25542 17013 25594
rect 23007 25542 23059 25594
rect 23071 25542 23123 25594
rect 23135 25542 23187 25594
rect 23199 25542 23251 25594
rect 23263 25542 23315 25594
rect 8760 25440 8812 25492
rect 10784 25440 10836 25492
rect 11796 25483 11848 25492
rect 11796 25449 11805 25483
rect 11805 25449 11839 25483
rect 11839 25449 11848 25483
rect 11796 25440 11848 25449
rect 11980 25440 12032 25492
rect 12164 25483 12216 25492
rect 12164 25449 12194 25483
rect 12194 25449 12216 25483
rect 12164 25440 12216 25449
rect 12256 25440 12308 25492
rect 5356 25304 5408 25356
rect 940 25236 992 25288
rect 4436 25236 4488 25288
rect 4988 25279 5040 25288
rect 4988 25245 4997 25279
rect 4997 25245 5031 25279
rect 5031 25245 5040 25279
rect 4988 25236 5040 25245
rect 6276 25168 6328 25220
rect 8208 25304 8260 25356
rect 8576 25279 8628 25288
rect 8576 25245 8585 25279
rect 8585 25245 8619 25279
rect 8619 25245 8628 25279
rect 8576 25236 8628 25245
rect 8852 25236 8904 25288
rect 9588 25304 9640 25356
rect 9956 25304 10008 25356
rect 14556 25440 14608 25492
rect 15292 25440 15344 25492
rect 14464 25347 14516 25356
rect 14464 25313 14473 25347
rect 14473 25313 14507 25347
rect 14507 25313 14516 25347
rect 14464 25304 14516 25313
rect 15200 25304 15252 25356
rect 17132 25440 17184 25492
rect 17500 25440 17552 25492
rect 22100 25440 22152 25492
rect 23664 25440 23716 25492
rect 16304 25304 16356 25356
rect 6920 25168 6972 25220
rect 7104 25100 7156 25152
rect 10876 25168 10928 25220
rect 12624 25168 12676 25220
rect 17316 25279 17368 25288
rect 17316 25245 17325 25279
rect 17325 25245 17359 25279
rect 17359 25245 17368 25279
rect 17316 25236 17368 25245
rect 17408 25279 17460 25288
rect 17408 25245 17417 25279
rect 17417 25245 17451 25279
rect 17451 25245 17460 25279
rect 17408 25236 17460 25245
rect 17776 25347 17828 25356
rect 17776 25313 17785 25347
rect 17785 25313 17819 25347
rect 17819 25313 17828 25347
rect 17776 25304 17828 25313
rect 18328 25279 18380 25288
rect 18328 25245 18337 25279
rect 18337 25245 18371 25279
rect 18371 25245 18380 25279
rect 18328 25236 18380 25245
rect 18420 25236 18472 25288
rect 19616 25304 19668 25356
rect 20720 25304 20772 25356
rect 20904 25304 20956 25356
rect 21456 25304 21508 25356
rect 22560 25304 22612 25356
rect 26332 25372 26384 25424
rect 9496 25100 9548 25152
rect 15108 25100 15160 25152
rect 17684 25168 17736 25220
rect 19248 25279 19300 25288
rect 19248 25245 19257 25279
rect 19257 25245 19291 25279
rect 19291 25245 19300 25279
rect 19248 25236 19300 25245
rect 25688 25279 25740 25288
rect 25688 25245 25697 25279
rect 25697 25245 25731 25279
rect 25731 25245 25740 25279
rect 25688 25236 25740 25245
rect 18052 25100 18104 25152
rect 18144 25100 18196 25152
rect 22652 25168 22704 25220
rect 18972 25100 19024 25152
rect 21364 25100 21416 25152
rect 24400 25143 24452 25152
rect 24400 25109 24409 25143
rect 24409 25109 24443 25143
rect 24443 25109 24452 25143
rect 24400 25100 24452 25109
rect 7252 24998 7304 25050
rect 7316 24998 7368 25050
rect 7380 24998 7432 25050
rect 7444 24998 7496 25050
rect 7508 24998 7560 25050
rect 13554 24998 13606 25050
rect 13618 24998 13670 25050
rect 13682 24998 13734 25050
rect 13746 24998 13798 25050
rect 13810 24998 13862 25050
rect 19856 24998 19908 25050
rect 19920 24998 19972 25050
rect 19984 24998 20036 25050
rect 20048 24998 20100 25050
rect 20112 24998 20164 25050
rect 26158 24998 26210 25050
rect 26222 24998 26274 25050
rect 26286 24998 26338 25050
rect 26350 24998 26402 25050
rect 26414 24998 26466 25050
rect 8576 24896 8628 24948
rect 9772 24896 9824 24948
rect 11336 24896 11388 24948
rect 11888 24939 11940 24948
rect 11888 24905 11897 24939
rect 11897 24905 11931 24939
rect 11931 24905 11940 24939
rect 11888 24896 11940 24905
rect 6000 24828 6052 24880
rect 6276 24828 6328 24880
rect 7656 24828 7708 24880
rect 6460 24803 6512 24812
rect 6460 24769 6469 24803
rect 6469 24769 6503 24803
rect 6503 24769 6512 24803
rect 6460 24760 6512 24769
rect 6920 24760 6972 24812
rect 7104 24760 7156 24812
rect 7196 24803 7248 24812
rect 7196 24769 7205 24803
rect 7205 24769 7239 24803
rect 7239 24769 7248 24803
rect 7196 24760 7248 24769
rect 8484 24760 8536 24812
rect 4436 24735 4488 24744
rect 4436 24701 4445 24735
rect 4445 24701 4479 24735
rect 4479 24701 4488 24735
rect 4436 24692 4488 24701
rect 4712 24735 4764 24744
rect 4712 24701 4721 24735
rect 4721 24701 4755 24735
rect 4755 24701 4764 24735
rect 4712 24692 4764 24701
rect 10876 24760 10928 24812
rect 13176 24896 13228 24948
rect 14280 24896 14332 24948
rect 14556 24760 14608 24812
rect 9404 24735 9456 24744
rect 9404 24701 9413 24735
rect 9413 24701 9447 24735
rect 9447 24701 9456 24735
rect 9404 24692 9456 24701
rect 9496 24692 9548 24744
rect 9864 24735 9916 24744
rect 9864 24701 9873 24735
rect 9873 24701 9907 24735
rect 9907 24701 9916 24735
rect 9864 24692 9916 24701
rect 11060 24692 11112 24744
rect 12348 24692 12400 24744
rect 13268 24735 13320 24744
rect 13268 24701 13277 24735
rect 13277 24701 13311 24735
rect 13311 24701 13320 24735
rect 13268 24692 13320 24701
rect 13820 24692 13872 24744
rect 14924 24692 14976 24744
rect 15476 24760 15528 24812
rect 16028 24760 16080 24812
rect 17500 24828 17552 24880
rect 18236 24828 18288 24880
rect 20904 24896 20956 24948
rect 20720 24828 20772 24880
rect 18880 24760 18932 24812
rect 24400 24828 24452 24880
rect 7564 24667 7616 24676
rect 7564 24633 7573 24667
rect 7573 24633 7607 24667
rect 7607 24633 7616 24667
rect 7564 24624 7616 24633
rect 15200 24624 15252 24676
rect 11520 24556 11572 24608
rect 13084 24556 13136 24608
rect 15752 24556 15804 24608
rect 16488 24556 16540 24608
rect 17868 24692 17920 24744
rect 17960 24556 18012 24608
rect 19248 24692 19300 24744
rect 19708 24735 19760 24744
rect 19708 24701 19717 24735
rect 19717 24701 19751 24735
rect 19751 24701 19760 24735
rect 19708 24692 19760 24701
rect 21272 24735 21324 24744
rect 21272 24701 21281 24735
rect 21281 24701 21315 24735
rect 21315 24701 21324 24735
rect 21272 24692 21324 24701
rect 18420 24624 18472 24676
rect 21916 24803 21968 24812
rect 21916 24769 21925 24803
rect 21925 24769 21959 24803
rect 21959 24769 21968 24803
rect 21916 24760 21968 24769
rect 22744 24760 22796 24812
rect 18788 24556 18840 24608
rect 19156 24556 19208 24608
rect 20628 24556 20680 24608
rect 22100 24556 22152 24608
rect 22376 24599 22428 24608
rect 22376 24565 22385 24599
rect 22385 24565 22419 24599
rect 22419 24565 22428 24599
rect 22376 24556 22428 24565
rect 23388 24556 23440 24608
rect 4101 24454 4153 24506
rect 4165 24454 4217 24506
rect 4229 24454 4281 24506
rect 4293 24454 4345 24506
rect 4357 24454 4409 24506
rect 10403 24454 10455 24506
rect 10467 24454 10519 24506
rect 10531 24454 10583 24506
rect 10595 24454 10647 24506
rect 10659 24454 10711 24506
rect 16705 24454 16757 24506
rect 16769 24454 16821 24506
rect 16833 24454 16885 24506
rect 16897 24454 16949 24506
rect 16961 24454 17013 24506
rect 23007 24454 23059 24506
rect 23071 24454 23123 24506
rect 23135 24454 23187 24506
rect 23199 24454 23251 24506
rect 23263 24454 23315 24506
rect 7196 24352 7248 24404
rect 9864 24352 9916 24404
rect 11060 24352 11112 24404
rect 11704 24352 11756 24404
rect 13268 24352 13320 24404
rect 16488 24352 16540 24404
rect 17500 24352 17552 24404
rect 20812 24395 20864 24404
rect 20812 24361 20821 24395
rect 20821 24361 20855 24395
rect 20855 24361 20864 24395
rect 20812 24352 20864 24361
rect 21272 24352 21324 24404
rect 9496 24284 9548 24336
rect 8300 24216 8352 24268
rect 11520 24284 11572 24336
rect 11244 24259 11296 24268
rect 11244 24225 11253 24259
rect 11253 24225 11287 24259
rect 11287 24225 11296 24259
rect 11244 24216 11296 24225
rect 5448 24148 5500 24200
rect 5816 24191 5868 24200
rect 5816 24157 5825 24191
rect 5825 24157 5859 24191
rect 5859 24157 5868 24191
rect 5816 24148 5868 24157
rect 4436 24012 4488 24064
rect 6460 24012 6512 24064
rect 6828 24012 6880 24064
rect 7104 24012 7156 24064
rect 11428 24191 11480 24200
rect 11428 24157 11437 24191
rect 11437 24157 11471 24191
rect 11471 24157 11480 24191
rect 11428 24148 11480 24157
rect 11520 24191 11572 24200
rect 11520 24157 11530 24191
rect 11530 24157 11564 24191
rect 11564 24157 11572 24191
rect 11520 24148 11572 24157
rect 11796 24191 11848 24200
rect 11796 24157 11805 24191
rect 11805 24157 11839 24191
rect 11839 24157 11848 24191
rect 11796 24148 11848 24157
rect 12072 24148 12124 24200
rect 12348 24148 12400 24200
rect 17868 24284 17920 24336
rect 15108 24216 15160 24268
rect 15292 24216 15344 24268
rect 15844 24259 15896 24268
rect 15844 24225 15853 24259
rect 15853 24225 15887 24259
rect 15887 24225 15896 24259
rect 15844 24216 15896 24225
rect 13820 24148 13872 24200
rect 13912 24148 13964 24200
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 12992 24080 13044 24132
rect 17868 24148 17920 24200
rect 17960 24148 18012 24200
rect 18604 24259 18656 24268
rect 18604 24225 18613 24259
rect 18613 24225 18647 24259
rect 18647 24225 18656 24259
rect 18604 24216 18656 24225
rect 18696 24148 18748 24200
rect 21180 24259 21232 24268
rect 21180 24225 21189 24259
rect 21189 24225 21223 24259
rect 21223 24225 21232 24259
rect 21180 24216 21232 24225
rect 22008 24216 22060 24268
rect 12532 24012 12584 24064
rect 13452 24055 13504 24064
rect 13452 24021 13461 24055
rect 13461 24021 13495 24055
rect 13495 24021 13504 24055
rect 13452 24012 13504 24021
rect 13912 24055 13964 24064
rect 13912 24021 13921 24055
rect 13921 24021 13955 24055
rect 13955 24021 13964 24055
rect 13912 24012 13964 24021
rect 14096 24055 14148 24064
rect 14096 24021 14105 24055
rect 14105 24021 14139 24055
rect 14139 24021 14148 24055
rect 14096 24012 14148 24021
rect 15568 24055 15620 24064
rect 15568 24021 15577 24055
rect 15577 24021 15611 24055
rect 15611 24021 15620 24055
rect 15568 24012 15620 24021
rect 17316 24012 17368 24064
rect 19340 24012 19392 24064
rect 22192 24148 22244 24200
rect 22928 24148 22980 24200
rect 22100 24080 22152 24132
rect 20352 24055 20404 24064
rect 20352 24021 20361 24055
rect 20361 24021 20395 24055
rect 20395 24021 20404 24055
rect 20352 24012 20404 24021
rect 20628 24012 20680 24064
rect 21732 24055 21784 24064
rect 21732 24021 21741 24055
rect 21741 24021 21775 24055
rect 21775 24021 21784 24055
rect 21732 24012 21784 24021
rect 23664 24012 23716 24064
rect 7252 23910 7304 23962
rect 7316 23910 7368 23962
rect 7380 23910 7432 23962
rect 7444 23910 7496 23962
rect 7508 23910 7560 23962
rect 13554 23910 13606 23962
rect 13618 23910 13670 23962
rect 13682 23910 13734 23962
rect 13746 23910 13798 23962
rect 13810 23910 13862 23962
rect 19856 23910 19908 23962
rect 19920 23910 19972 23962
rect 19984 23910 20036 23962
rect 20048 23910 20100 23962
rect 20112 23910 20164 23962
rect 26158 23910 26210 23962
rect 26222 23910 26274 23962
rect 26286 23910 26338 23962
rect 26350 23910 26402 23962
rect 26414 23910 26466 23962
rect 4712 23808 4764 23860
rect 7656 23808 7708 23860
rect 4712 23647 4764 23656
rect 4712 23613 4721 23647
rect 4721 23613 4755 23647
rect 4755 23613 4764 23647
rect 4712 23604 4764 23613
rect 4988 23604 5040 23656
rect 5356 23672 5408 23724
rect 6460 23672 6512 23724
rect 8300 23851 8352 23860
rect 8300 23817 8309 23851
rect 8309 23817 8343 23851
rect 8343 23817 8352 23851
rect 8300 23808 8352 23817
rect 14096 23808 14148 23860
rect 14924 23851 14976 23860
rect 14924 23817 14933 23851
rect 14933 23817 14967 23851
rect 14967 23817 14976 23851
rect 14924 23808 14976 23817
rect 15200 23808 15252 23860
rect 15568 23808 15620 23860
rect 15108 23740 15160 23792
rect 9036 23715 9088 23724
rect 9036 23681 9045 23715
rect 9045 23681 9079 23715
rect 9079 23681 9088 23715
rect 9036 23672 9088 23681
rect 4528 23511 4580 23520
rect 4528 23477 4537 23511
rect 4537 23477 4571 23511
rect 4571 23477 4580 23511
rect 4528 23468 4580 23477
rect 5448 23604 5500 23656
rect 6920 23604 6972 23656
rect 9312 23715 9364 23724
rect 9312 23681 9321 23715
rect 9321 23681 9355 23715
rect 9355 23681 9364 23715
rect 9312 23672 9364 23681
rect 11520 23672 11572 23724
rect 13084 23672 13136 23724
rect 13176 23715 13228 23724
rect 13176 23681 13185 23715
rect 13185 23681 13219 23715
rect 13219 23681 13228 23715
rect 13176 23672 13228 23681
rect 14924 23672 14976 23724
rect 17960 23808 18012 23860
rect 17960 23672 18012 23724
rect 19708 23808 19760 23860
rect 21732 23808 21784 23860
rect 22652 23808 22704 23860
rect 23664 23808 23716 23860
rect 18236 23740 18288 23792
rect 19156 23740 19208 23792
rect 12532 23604 12584 23656
rect 12624 23647 12676 23656
rect 12624 23613 12633 23647
rect 12633 23613 12667 23647
rect 12667 23613 12676 23647
rect 12624 23604 12676 23613
rect 17040 23604 17092 23656
rect 17316 23604 17368 23656
rect 18972 23604 19024 23656
rect 19340 23715 19392 23724
rect 19340 23681 19350 23715
rect 19350 23681 19384 23715
rect 19384 23681 19392 23715
rect 19340 23672 19392 23681
rect 6276 23468 6328 23520
rect 8484 23468 8536 23520
rect 9128 23511 9180 23520
rect 9128 23477 9137 23511
rect 9137 23477 9171 23511
rect 9171 23477 9180 23511
rect 9128 23468 9180 23477
rect 10324 23468 10376 23520
rect 11980 23511 12032 23520
rect 11980 23477 11989 23511
rect 11989 23477 12023 23511
rect 12023 23477 12032 23511
rect 11980 23468 12032 23477
rect 12992 23511 13044 23520
rect 12992 23477 13001 23511
rect 13001 23477 13035 23511
rect 13035 23477 13044 23511
rect 12992 23468 13044 23477
rect 13452 23468 13504 23520
rect 15936 23468 15988 23520
rect 18144 23468 18196 23520
rect 18512 23511 18564 23520
rect 18512 23477 18521 23511
rect 18521 23477 18555 23511
rect 18555 23477 18564 23511
rect 18512 23468 18564 23477
rect 18880 23468 18932 23520
rect 19064 23468 19116 23520
rect 20352 23672 20404 23724
rect 20812 23672 20864 23724
rect 22100 23715 22152 23724
rect 22100 23681 22109 23715
rect 22109 23681 22143 23715
rect 22143 23681 22152 23715
rect 22100 23672 22152 23681
rect 22008 23604 22060 23656
rect 22376 23715 22428 23724
rect 22376 23681 22385 23715
rect 22385 23681 22419 23715
rect 22419 23681 22428 23715
rect 22376 23672 22428 23681
rect 22652 23672 22704 23724
rect 22744 23604 22796 23656
rect 19892 23511 19944 23520
rect 19892 23477 19901 23511
rect 19901 23477 19935 23511
rect 19935 23477 19944 23511
rect 19892 23468 19944 23477
rect 20076 23468 20128 23520
rect 21916 23511 21968 23520
rect 21916 23477 21925 23511
rect 21925 23477 21959 23511
rect 21959 23477 21968 23511
rect 21916 23468 21968 23477
rect 22652 23536 22704 23588
rect 22560 23468 22612 23520
rect 23388 23468 23440 23520
rect 4101 23366 4153 23418
rect 4165 23366 4217 23418
rect 4229 23366 4281 23418
rect 4293 23366 4345 23418
rect 4357 23366 4409 23418
rect 10403 23366 10455 23418
rect 10467 23366 10519 23418
rect 10531 23366 10583 23418
rect 10595 23366 10647 23418
rect 10659 23366 10711 23418
rect 16705 23366 16757 23418
rect 16769 23366 16821 23418
rect 16833 23366 16885 23418
rect 16897 23366 16949 23418
rect 16961 23366 17013 23418
rect 23007 23366 23059 23418
rect 23071 23366 23123 23418
rect 23135 23366 23187 23418
rect 23199 23366 23251 23418
rect 23263 23366 23315 23418
rect 6460 23264 6512 23316
rect 6920 23239 6972 23248
rect 6920 23205 6929 23239
rect 6929 23205 6963 23239
rect 6963 23205 6972 23239
rect 6920 23196 6972 23205
rect 4436 23128 4488 23180
rect 9036 23264 9088 23316
rect 10324 23264 10376 23316
rect 12072 23264 12124 23316
rect 12808 23264 12860 23316
rect 16028 23264 16080 23316
rect 17040 23264 17092 23316
rect 18696 23264 18748 23316
rect 8300 23128 8352 23180
rect 12624 23128 12676 23180
rect 13360 23128 13412 23180
rect 16212 23128 16264 23180
rect 17316 23128 17368 23180
rect 17408 23171 17460 23180
rect 17408 23137 17417 23171
rect 17417 23137 17451 23171
rect 17451 23137 17460 23171
rect 17408 23128 17460 23137
rect 5448 23060 5500 23112
rect 6000 23060 6052 23112
rect 6276 22992 6328 23044
rect 4528 22924 4580 22976
rect 6920 23060 6972 23112
rect 10232 23103 10284 23112
rect 10232 23069 10241 23103
rect 10241 23069 10275 23103
rect 10275 23069 10284 23103
rect 10232 23060 10284 23069
rect 6552 23035 6604 23044
rect 6552 23001 6561 23035
rect 6561 23001 6595 23035
rect 6595 23001 6604 23035
rect 6552 22992 6604 23001
rect 7196 22992 7248 23044
rect 6828 22924 6880 22976
rect 7104 22924 7156 22976
rect 10140 22992 10192 23044
rect 7656 22924 7708 22976
rect 10876 22924 10928 22976
rect 11428 22924 11480 22976
rect 12808 23103 12860 23112
rect 12808 23069 12817 23103
rect 12817 23069 12851 23103
rect 12851 23069 12860 23103
rect 12808 23060 12860 23069
rect 12900 23103 12952 23112
rect 12900 23069 12909 23103
rect 12909 23069 12943 23103
rect 12943 23069 12952 23103
rect 12900 23060 12952 23069
rect 13084 23103 13136 23112
rect 13084 23069 13093 23103
rect 13093 23069 13127 23103
rect 13127 23069 13136 23103
rect 13084 23060 13136 23069
rect 16396 23103 16448 23112
rect 16396 23069 16405 23103
rect 16405 23069 16439 23103
rect 16439 23069 16448 23103
rect 16396 23060 16448 23069
rect 17776 23060 17828 23112
rect 18512 23060 18564 23112
rect 18788 23060 18840 23112
rect 20076 23264 20128 23316
rect 22008 23264 22060 23316
rect 20628 23196 20680 23248
rect 20260 23128 20312 23180
rect 19248 23103 19300 23112
rect 19248 23069 19257 23103
rect 19257 23069 19291 23103
rect 19291 23069 19300 23103
rect 19248 23060 19300 23069
rect 22376 23264 22428 23316
rect 22928 23264 22980 23316
rect 22560 23196 22612 23248
rect 22192 23060 22244 23112
rect 15936 22992 15988 23044
rect 15476 22924 15528 22976
rect 15844 22924 15896 22976
rect 16304 23035 16356 23044
rect 16304 23001 16313 23035
rect 16313 23001 16347 23035
rect 16347 23001 16356 23035
rect 16304 22992 16356 23001
rect 18788 22967 18840 22976
rect 18788 22933 18797 22967
rect 18797 22933 18831 22967
rect 18831 22933 18840 22967
rect 18788 22924 18840 22933
rect 20996 22992 21048 23044
rect 21088 22967 21140 22976
rect 21088 22933 21097 22967
rect 21097 22933 21131 22967
rect 21131 22933 21140 22967
rect 21088 22924 21140 22933
rect 21456 22992 21508 23044
rect 22468 22924 22520 22976
rect 22744 23128 22796 23180
rect 22744 22924 22796 22976
rect 7252 22822 7304 22874
rect 7316 22822 7368 22874
rect 7380 22822 7432 22874
rect 7444 22822 7496 22874
rect 7508 22822 7560 22874
rect 13554 22822 13606 22874
rect 13618 22822 13670 22874
rect 13682 22822 13734 22874
rect 13746 22822 13798 22874
rect 13810 22822 13862 22874
rect 19856 22822 19908 22874
rect 19920 22822 19972 22874
rect 19984 22822 20036 22874
rect 20048 22822 20100 22874
rect 20112 22822 20164 22874
rect 26158 22822 26210 22874
rect 26222 22822 26274 22874
rect 26286 22822 26338 22874
rect 26350 22822 26402 22874
rect 26414 22822 26466 22874
rect 3148 22720 3200 22772
rect 5356 22720 5408 22772
rect 7104 22720 7156 22772
rect 8300 22720 8352 22772
rect 5448 22652 5500 22704
rect 6184 22652 6236 22704
rect 9128 22720 9180 22772
rect 11520 22763 11572 22772
rect 11520 22729 11529 22763
rect 11529 22729 11563 22763
rect 11563 22729 11572 22763
rect 11520 22720 11572 22729
rect 11980 22720 12032 22772
rect 14832 22720 14884 22772
rect 16304 22720 16356 22772
rect 16396 22720 16448 22772
rect 18788 22720 18840 22772
rect 4988 22627 5040 22636
rect 4988 22593 4997 22627
rect 4997 22593 5031 22627
rect 5031 22593 5040 22627
rect 4988 22584 5040 22593
rect 2688 22559 2740 22568
rect 2688 22525 2697 22559
rect 2697 22525 2731 22559
rect 2731 22525 2740 22559
rect 2688 22516 2740 22525
rect 3516 22516 3568 22568
rect 4712 22516 4764 22568
rect 5816 22627 5868 22636
rect 5816 22593 5825 22627
rect 5825 22593 5859 22627
rect 5859 22593 5868 22627
rect 5816 22584 5868 22593
rect 6828 22584 6880 22636
rect 7104 22627 7156 22636
rect 7104 22593 7113 22627
rect 7113 22593 7147 22627
rect 7147 22593 7156 22627
rect 7104 22584 7156 22593
rect 9864 22652 9916 22704
rect 11244 22652 11296 22704
rect 11152 22627 11204 22636
rect 11152 22593 11161 22627
rect 11161 22593 11195 22627
rect 11195 22593 11204 22627
rect 11152 22584 11204 22593
rect 8484 22516 8536 22568
rect 9772 22516 9824 22568
rect 10324 22516 10376 22568
rect 11980 22559 12032 22568
rect 11980 22525 11989 22559
rect 11989 22525 12023 22559
rect 12023 22525 12032 22559
rect 11980 22516 12032 22525
rect 15292 22652 15344 22704
rect 15568 22584 15620 22636
rect 12440 22516 12492 22568
rect 14740 22559 14792 22568
rect 14740 22525 14749 22559
rect 14749 22525 14783 22559
rect 14783 22525 14792 22559
rect 14740 22516 14792 22525
rect 15016 22516 15068 22568
rect 16028 22559 16080 22568
rect 16028 22525 16037 22559
rect 16037 22525 16071 22559
rect 16071 22525 16080 22559
rect 16028 22516 16080 22525
rect 19248 22652 19300 22704
rect 20812 22763 20864 22772
rect 20812 22729 20821 22763
rect 20821 22729 20855 22763
rect 20855 22729 20864 22763
rect 20812 22720 20864 22729
rect 21456 22720 21508 22772
rect 21272 22584 21324 22636
rect 22192 22652 22244 22704
rect 22100 22584 22152 22636
rect 23388 22720 23440 22772
rect 22468 22652 22520 22704
rect 5908 22380 5960 22432
rect 6276 22380 6328 22432
rect 9956 22423 10008 22432
rect 9956 22389 9965 22423
rect 9965 22389 9999 22423
rect 9999 22389 10008 22423
rect 9956 22380 10008 22389
rect 10968 22423 11020 22432
rect 10968 22389 10977 22423
rect 10977 22389 11011 22423
rect 11011 22389 11020 22423
rect 10968 22380 11020 22389
rect 12348 22423 12400 22432
rect 12348 22389 12357 22423
rect 12357 22389 12391 22423
rect 12391 22389 12400 22423
rect 12348 22380 12400 22389
rect 14004 22380 14056 22432
rect 15476 22423 15528 22432
rect 15476 22389 15485 22423
rect 15485 22389 15519 22423
rect 15519 22389 15528 22423
rect 15476 22380 15528 22389
rect 15844 22380 15896 22432
rect 16304 22380 16356 22432
rect 20904 22423 20956 22432
rect 20904 22389 20913 22423
rect 20913 22389 20947 22423
rect 20947 22389 20956 22423
rect 20904 22380 20956 22389
rect 22560 22380 22612 22432
rect 4101 22278 4153 22330
rect 4165 22278 4217 22330
rect 4229 22278 4281 22330
rect 4293 22278 4345 22330
rect 4357 22278 4409 22330
rect 10403 22278 10455 22330
rect 10467 22278 10519 22330
rect 10531 22278 10583 22330
rect 10595 22278 10647 22330
rect 10659 22278 10711 22330
rect 16705 22278 16757 22330
rect 16769 22278 16821 22330
rect 16833 22278 16885 22330
rect 16897 22278 16949 22330
rect 16961 22278 17013 22330
rect 23007 22278 23059 22330
rect 23071 22278 23123 22330
rect 23135 22278 23187 22330
rect 23199 22278 23251 22330
rect 23263 22278 23315 22330
rect 6920 22176 6972 22228
rect 7656 22176 7708 22228
rect 9588 22176 9640 22228
rect 6828 22040 6880 22092
rect 5540 22015 5592 22024
rect 5540 21981 5549 22015
rect 5549 21981 5583 22015
rect 5583 21981 5592 22015
rect 5540 21972 5592 21981
rect 6920 21972 6972 22024
rect 12992 22176 13044 22228
rect 14832 22176 14884 22228
rect 10232 22040 10284 22092
rect 13176 22040 13228 22092
rect 5816 21947 5868 21956
rect 5816 21913 5825 21947
rect 5825 21913 5859 21947
rect 5859 21913 5868 21947
rect 5816 21904 5868 21913
rect 8024 21836 8076 21888
rect 8576 21836 8628 21888
rect 10048 22015 10100 22024
rect 10048 21981 10057 22015
rect 10057 21981 10091 22015
rect 10091 21981 10100 22015
rect 10048 21972 10100 21981
rect 10600 21972 10652 22024
rect 12072 21972 12124 22024
rect 15476 22176 15528 22228
rect 16120 22176 16172 22228
rect 17868 22176 17920 22228
rect 22192 22176 22244 22228
rect 22376 22151 22428 22160
rect 22376 22117 22385 22151
rect 22385 22117 22419 22151
rect 22419 22117 22428 22151
rect 22376 22108 22428 22117
rect 15568 22083 15620 22092
rect 15568 22049 15577 22083
rect 15577 22049 15611 22083
rect 15611 22049 15620 22083
rect 15568 22040 15620 22049
rect 18512 22040 18564 22092
rect 19248 22040 19300 22092
rect 9772 21904 9824 21956
rect 10232 21947 10284 21956
rect 10232 21913 10241 21947
rect 10241 21913 10275 21947
rect 10275 21913 10284 21947
rect 10232 21904 10284 21913
rect 10324 21947 10376 21956
rect 10324 21913 10333 21947
rect 10333 21913 10367 21947
rect 10367 21913 10376 21947
rect 10324 21904 10376 21913
rect 9588 21879 9640 21888
rect 9588 21845 9597 21879
rect 9597 21845 9631 21879
rect 9631 21845 9640 21879
rect 9588 21836 9640 21845
rect 9956 21836 10008 21888
rect 10968 21947 11020 21956
rect 10968 21913 10977 21947
rect 10977 21913 11011 21947
rect 11011 21913 11020 21947
rect 10968 21904 11020 21913
rect 12532 21947 12584 21956
rect 10600 21879 10652 21888
rect 10600 21845 10609 21879
rect 10609 21845 10643 21879
rect 10643 21845 10652 21879
rect 10600 21836 10652 21845
rect 10784 21836 10836 21888
rect 11060 21836 11112 21888
rect 12532 21913 12541 21947
rect 12541 21913 12575 21947
rect 12575 21913 12584 21947
rect 12532 21904 12584 21913
rect 14372 21947 14424 21956
rect 14372 21913 14381 21947
rect 14381 21913 14415 21947
rect 14415 21913 14424 21947
rect 14372 21904 14424 21913
rect 14464 21947 14516 21956
rect 14464 21913 14473 21947
rect 14473 21913 14507 21947
rect 14507 21913 14516 21947
rect 14464 21904 14516 21913
rect 14740 21972 14792 22024
rect 16120 22015 16172 22024
rect 16120 21981 16129 22015
rect 16129 21981 16163 22015
rect 16163 21981 16172 22015
rect 16120 21972 16172 21981
rect 16212 21972 16264 22024
rect 15200 21904 15252 21956
rect 17500 21972 17552 22024
rect 18696 21972 18748 22024
rect 20720 22015 20772 22024
rect 20720 21981 20729 22015
rect 20729 21981 20763 22015
rect 20763 21981 20772 22015
rect 20720 21972 20772 21981
rect 22560 22040 22612 22092
rect 12440 21879 12492 21888
rect 12440 21845 12449 21879
rect 12449 21845 12483 21879
rect 12483 21845 12492 21879
rect 12440 21836 12492 21845
rect 13912 21879 13964 21888
rect 13912 21845 13921 21879
rect 13921 21845 13955 21879
rect 13955 21845 13964 21879
rect 13912 21836 13964 21845
rect 14096 21879 14148 21888
rect 14096 21845 14105 21879
rect 14105 21845 14139 21879
rect 14139 21845 14148 21879
rect 14096 21836 14148 21845
rect 16488 21879 16540 21888
rect 16488 21845 16497 21879
rect 16497 21845 16531 21879
rect 16531 21845 16540 21879
rect 16488 21836 16540 21845
rect 19340 21904 19392 21956
rect 21548 21947 21600 21956
rect 21548 21913 21557 21947
rect 21557 21913 21591 21947
rect 21591 21913 21600 21947
rect 21548 21904 21600 21913
rect 21916 22015 21968 22024
rect 21916 21981 21925 22015
rect 21925 21981 21959 22015
rect 21959 21981 21968 22015
rect 21916 21972 21968 21981
rect 22560 21904 22612 21956
rect 22744 21904 22796 21956
rect 17040 21879 17092 21888
rect 17040 21845 17049 21879
rect 17049 21845 17083 21879
rect 17083 21845 17092 21879
rect 17040 21836 17092 21845
rect 17408 21879 17460 21888
rect 17408 21845 17417 21879
rect 17417 21845 17451 21879
rect 17451 21845 17460 21879
rect 17408 21836 17460 21845
rect 20352 21879 20404 21888
rect 20352 21845 20361 21879
rect 20361 21845 20395 21879
rect 20395 21845 20404 21879
rect 20352 21836 20404 21845
rect 22836 21879 22888 21888
rect 22836 21845 22845 21879
rect 22845 21845 22879 21879
rect 22879 21845 22888 21879
rect 22836 21836 22888 21845
rect 7252 21734 7304 21786
rect 7316 21734 7368 21786
rect 7380 21734 7432 21786
rect 7444 21734 7496 21786
rect 7508 21734 7560 21786
rect 13554 21734 13606 21786
rect 13618 21734 13670 21786
rect 13682 21734 13734 21786
rect 13746 21734 13798 21786
rect 13810 21734 13862 21786
rect 19856 21734 19908 21786
rect 19920 21734 19972 21786
rect 19984 21734 20036 21786
rect 20048 21734 20100 21786
rect 20112 21734 20164 21786
rect 26158 21734 26210 21786
rect 26222 21734 26274 21786
rect 26286 21734 26338 21786
rect 26350 21734 26402 21786
rect 26414 21734 26466 21786
rect 2688 21564 2740 21616
rect 5540 21632 5592 21684
rect 1952 21496 2004 21548
rect 3148 21564 3200 21616
rect 10140 21632 10192 21684
rect 11060 21632 11112 21684
rect 11152 21632 11204 21684
rect 12348 21632 12400 21684
rect 12440 21632 12492 21684
rect 8576 21607 8628 21616
rect 8576 21573 8585 21607
rect 8585 21573 8619 21607
rect 8619 21573 8628 21607
rect 8576 21564 8628 21573
rect 10048 21564 10100 21616
rect 10600 21564 10652 21616
rect 6276 21496 6328 21548
rect 8300 21539 8352 21548
rect 8300 21505 8309 21539
rect 8309 21505 8343 21539
rect 8343 21505 8352 21539
rect 8300 21496 8352 21505
rect 9588 21496 9640 21548
rect 9864 21496 9916 21548
rect 10784 21496 10836 21548
rect 11980 21539 12032 21548
rect 11980 21505 11989 21539
rect 11989 21505 12023 21539
rect 12023 21505 12032 21539
rect 11980 21496 12032 21505
rect 12808 21564 12860 21616
rect 13360 21539 13412 21548
rect 13360 21505 13370 21539
rect 13370 21505 13404 21539
rect 13404 21505 13412 21539
rect 13360 21496 13412 21505
rect 13544 21607 13596 21616
rect 13544 21573 13553 21607
rect 13553 21573 13587 21607
rect 13587 21573 13596 21607
rect 13544 21564 13596 21573
rect 14372 21632 14424 21684
rect 16212 21632 16264 21684
rect 13912 21564 13964 21616
rect 14924 21564 14976 21616
rect 16488 21564 16540 21616
rect 17960 21564 18012 21616
rect 3056 21471 3108 21480
rect 3056 21437 3065 21471
rect 3065 21437 3099 21471
rect 3099 21437 3108 21471
rect 3056 21428 3108 21437
rect 4804 21471 4856 21480
rect 4804 21437 4813 21471
rect 4813 21437 4847 21471
rect 4847 21437 4856 21471
rect 4804 21428 4856 21437
rect 6368 21428 6420 21480
rect 7472 21428 7524 21480
rect 8024 21471 8076 21480
rect 8024 21437 8033 21471
rect 8033 21437 8067 21471
rect 8067 21437 8076 21471
rect 8024 21428 8076 21437
rect 10324 21428 10376 21480
rect 11428 21428 11480 21480
rect 12072 21428 12124 21480
rect 12256 21428 12308 21480
rect 12808 21428 12860 21480
rect 13176 21428 13228 21480
rect 14740 21428 14792 21480
rect 16028 21428 16080 21480
rect 16580 21496 16632 21548
rect 17040 21428 17092 21480
rect 20352 21632 20404 21684
rect 22836 21632 22888 21684
rect 20996 21564 21048 21616
rect 19248 21496 19300 21548
rect 21272 21496 21324 21548
rect 20904 21428 20956 21480
rect 22652 21496 22704 21548
rect 23388 21496 23440 21548
rect 25688 21539 25740 21548
rect 25688 21505 25697 21539
rect 25697 21505 25731 21539
rect 25731 21505 25740 21539
rect 25688 21496 25740 21505
rect 940 21292 992 21344
rect 6000 21292 6052 21344
rect 7288 21292 7340 21344
rect 7380 21335 7432 21344
rect 7380 21301 7389 21335
rect 7389 21301 7423 21335
rect 7423 21301 7432 21335
rect 7380 21292 7432 21301
rect 10140 21335 10192 21344
rect 10140 21301 10149 21335
rect 10149 21301 10183 21335
rect 10183 21301 10192 21335
rect 10140 21292 10192 21301
rect 12440 21292 12492 21344
rect 13912 21335 13964 21344
rect 13912 21301 13921 21335
rect 13921 21301 13955 21335
rect 13955 21301 13964 21335
rect 13912 21292 13964 21301
rect 18696 21292 18748 21344
rect 25872 21335 25924 21344
rect 25872 21301 25881 21335
rect 25881 21301 25915 21335
rect 25915 21301 25924 21335
rect 25872 21292 25924 21301
rect 4101 21190 4153 21242
rect 4165 21190 4217 21242
rect 4229 21190 4281 21242
rect 4293 21190 4345 21242
rect 4357 21190 4409 21242
rect 10403 21190 10455 21242
rect 10467 21190 10519 21242
rect 10531 21190 10583 21242
rect 10595 21190 10647 21242
rect 10659 21190 10711 21242
rect 16705 21190 16757 21242
rect 16769 21190 16821 21242
rect 16833 21190 16885 21242
rect 16897 21190 16949 21242
rect 16961 21190 17013 21242
rect 23007 21190 23059 21242
rect 23071 21190 23123 21242
rect 23135 21190 23187 21242
rect 23199 21190 23251 21242
rect 23263 21190 23315 21242
rect 3056 21088 3108 21140
rect 5816 21088 5868 21140
rect 6552 21088 6604 21140
rect 6736 21088 6788 21140
rect 4160 20952 4212 21004
rect 5264 20952 5316 21004
rect 4804 20884 4856 20936
rect 4804 20748 4856 20800
rect 5264 20816 5316 20868
rect 6184 20884 6236 20936
rect 9312 21088 9364 21140
rect 10140 21088 10192 21140
rect 6644 20952 6696 21004
rect 7380 20952 7432 21004
rect 7104 20884 7156 20936
rect 6184 20748 6236 20800
rect 6552 20748 6604 20800
rect 7196 20816 7248 20868
rect 7288 20859 7340 20868
rect 7288 20825 7297 20859
rect 7297 20825 7331 20859
rect 7331 20825 7340 20859
rect 7288 20816 7340 20825
rect 7472 20859 7524 20868
rect 7472 20825 7481 20859
rect 7481 20825 7515 20859
rect 7515 20825 7524 20859
rect 9404 20952 9456 21004
rect 7472 20816 7524 20825
rect 8116 20816 8168 20868
rect 15108 21088 15160 21140
rect 16120 21088 16172 21140
rect 16396 21088 16448 21140
rect 20996 21088 21048 21140
rect 23388 21088 23440 21140
rect 17960 21020 18012 21072
rect 16396 20952 16448 21004
rect 16488 20995 16540 21004
rect 16488 20961 16497 20995
rect 16497 20961 16531 20995
rect 16531 20961 16540 20995
rect 16488 20952 16540 20961
rect 17408 20952 17460 21004
rect 12532 20927 12584 20936
rect 12532 20893 12541 20927
rect 12541 20893 12575 20927
rect 12575 20893 12584 20927
rect 12532 20884 12584 20893
rect 14004 20884 14056 20936
rect 13084 20816 13136 20868
rect 17776 20884 17828 20936
rect 18972 20952 19024 21004
rect 21088 20952 21140 21004
rect 22100 20952 22152 21004
rect 18420 20884 18472 20936
rect 21456 20927 21508 20936
rect 21456 20893 21465 20927
rect 21465 20893 21499 20927
rect 21499 20893 21508 20927
rect 21456 20884 21508 20893
rect 9956 20748 10008 20800
rect 14556 20748 14608 20800
rect 15844 20816 15896 20868
rect 18052 20816 18104 20868
rect 21272 20816 21324 20868
rect 20996 20791 21048 20800
rect 20996 20757 21005 20791
rect 21005 20757 21039 20791
rect 21039 20757 21048 20791
rect 20996 20748 21048 20757
rect 7252 20646 7304 20698
rect 7316 20646 7368 20698
rect 7380 20646 7432 20698
rect 7444 20646 7496 20698
rect 7508 20646 7560 20698
rect 13554 20646 13606 20698
rect 13618 20646 13670 20698
rect 13682 20646 13734 20698
rect 13746 20646 13798 20698
rect 13810 20646 13862 20698
rect 19856 20646 19908 20698
rect 19920 20646 19972 20698
rect 19984 20646 20036 20698
rect 20048 20646 20100 20698
rect 20112 20646 20164 20698
rect 26158 20646 26210 20698
rect 26222 20646 26274 20698
rect 26286 20646 26338 20698
rect 26350 20646 26402 20698
rect 26414 20646 26466 20698
rect 5356 20544 5408 20596
rect 6644 20544 6696 20596
rect 6736 20587 6788 20596
rect 6736 20553 6745 20587
rect 6745 20553 6779 20587
rect 6779 20553 6788 20587
rect 6736 20544 6788 20553
rect 4896 20476 4948 20528
rect 7104 20544 7156 20596
rect 2780 20340 2832 20392
rect 4804 20408 4856 20460
rect 5448 20408 5500 20460
rect 6000 20408 6052 20460
rect 6184 20451 6236 20460
rect 6184 20417 6193 20451
rect 6193 20417 6227 20451
rect 6227 20417 6236 20451
rect 6184 20408 6236 20417
rect 3332 20383 3384 20392
rect 3332 20349 3341 20383
rect 3341 20349 3375 20383
rect 3375 20349 3384 20383
rect 3332 20340 3384 20349
rect 3976 20340 4028 20392
rect 4160 20340 4212 20392
rect 4436 20340 4488 20392
rect 6644 20408 6696 20460
rect 12440 20544 12492 20596
rect 14740 20544 14792 20596
rect 9956 20476 10008 20528
rect 14924 20476 14976 20528
rect 15476 20476 15528 20528
rect 5632 20272 5684 20324
rect 5724 20315 5776 20324
rect 5724 20281 5733 20315
rect 5733 20281 5767 20315
rect 5767 20281 5776 20315
rect 5724 20272 5776 20281
rect 5816 20272 5868 20324
rect 12900 20408 12952 20460
rect 16120 20544 16172 20596
rect 17040 20587 17092 20596
rect 17040 20553 17049 20587
rect 17049 20553 17083 20587
rect 17083 20553 17092 20587
rect 17040 20544 17092 20553
rect 17500 20587 17552 20596
rect 17500 20553 17509 20587
rect 17509 20553 17543 20587
rect 17543 20553 17552 20587
rect 17500 20544 17552 20553
rect 15936 20476 15988 20528
rect 16396 20476 16448 20528
rect 19340 20544 19392 20596
rect 16120 20451 16172 20460
rect 16120 20417 16129 20451
rect 16129 20417 16163 20451
rect 16163 20417 16172 20451
rect 16120 20408 16172 20417
rect 16212 20451 16264 20460
rect 16212 20417 16221 20451
rect 16221 20417 16255 20451
rect 16255 20417 16264 20451
rect 16212 20408 16264 20417
rect 18420 20476 18472 20528
rect 22100 20476 22152 20528
rect 23296 20587 23348 20596
rect 23296 20553 23305 20587
rect 23305 20553 23339 20587
rect 23339 20553 23348 20587
rect 23296 20544 23348 20553
rect 25688 20544 25740 20596
rect 23388 20476 23440 20528
rect 17592 20451 17644 20460
rect 9680 20340 9732 20392
rect 10784 20340 10836 20392
rect 12256 20383 12308 20392
rect 12256 20349 12265 20383
rect 12265 20349 12299 20383
rect 12299 20349 12308 20383
rect 12256 20340 12308 20349
rect 12440 20340 12492 20392
rect 13084 20383 13136 20392
rect 13084 20349 13093 20383
rect 13093 20349 13127 20383
rect 13127 20349 13136 20383
rect 13084 20340 13136 20349
rect 14096 20340 14148 20392
rect 17040 20340 17092 20392
rect 17592 20417 17601 20451
rect 17601 20417 17635 20451
rect 17635 20417 17644 20451
rect 17592 20408 17644 20417
rect 17684 20408 17736 20460
rect 18052 20408 18104 20460
rect 9864 20272 9916 20324
rect 10968 20272 11020 20324
rect 12072 20272 12124 20324
rect 12532 20272 12584 20324
rect 18696 20451 18748 20460
rect 18696 20417 18706 20451
rect 18706 20417 18740 20451
rect 18740 20417 18748 20451
rect 18696 20408 18748 20417
rect 18880 20451 18932 20460
rect 18880 20417 18889 20451
rect 18889 20417 18923 20451
rect 18923 20417 18932 20451
rect 18880 20408 18932 20417
rect 18972 20451 19024 20460
rect 18972 20417 18981 20451
rect 18981 20417 19015 20451
rect 19015 20417 19024 20451
rect 18972 20408 19024 20417
rect 19064 20451 19116 20460
rect 19064 20417 19097 20451
rect 19097 20417 19116 20451
rect 19064 20408 19116 20417
rect 20260 20408 20312 20460
rect 22836 20408 22888 20460
rect 23848 20451 23900 20460
rect 23848 20417 23857 20451
rect 23857 20417 23891 20451
rect 23891 20417 23900 20451
rect 23848 20408 23900 20417
rect 23940 20451 23992 20460
rect 23940 20417 23949 20451
rect 23949 20417 23983 20451
rect 23983 20417 23992 20451
rect 23940 20408 23992 20417
rect 24032 20451 24084 20460
rect 24032 20417 24041 20451
rect 24041 20417 24075 20451
rect 24075 20417 24084 20451
rect 24032 20408 24084 20417
rect 18328 20340 18380 20392
rect 22652 20340 22704 20392
rect 25136 20408 25188 20460
rect 2136 20247 2188 20256
rect 2136 20213 2145 20247
rect 2145 20213 2179 20247
rect 2179 20213 2188 20247
rect 2136 20204 2188 20213
rect 2412 20247 2464 20256
rect 2412 20213 2421 20247
rect 2421 20213 2455 20247
rect 2455 20213 2464 20247
rect 2412 20204 2464 20213
rect 9220 20204 9272 20256
rect 11612 20247 11664 20256
rect 11612 20213 11621 20247
rect 11621 20213 11655 20247
rect 11655 20213 11664 20247
rect 11612 20204 11664 20213
rect 16580 20204 16632 20256
rect 17684 20204 17736 20256
rect 18972 20204 19024 20256
rect 20996 20204 21048 20256
rect 21364 20204 21416 20256
rect 21456 20204 21508 20256
rect 23664 20247 23716 20256
rect 23664 20213 23673 20247
rect 23673 20213 23707 20247
rect 23707 20213 23716 20247
rect 23664 20204 23716 20213
rect 4101 20102 4153 20154
rect 4165 20102 4217 20154
rect 4229 20102 4281 20154
rect 4293 20102 4345 20154
rect 4357 20102 4409 20154
rect 10403 20102 10455 20154
rect 10467 20102 10519 20154
rect 10531 20102 10583 20154
rect 10595 20102 10647 20154
rect 10659 20102 10711 20154
rect 16705 20102 16757 20154
rect 16769 20102 16821 20154
rect 16833 20102 16885 20154
rect 16897 20102 16949 20154
rect 16961 20102 17013 20154
rect 23007 20102 23059 20154
rect 23071 20102 23123 20154
rect 23135 20102 23187 20154
rect 23199 20102 23251 20154
rect 23263 20102 23315 20154
rect 4436 20043 4488 20052
rect 4436 20009 4445 20043
rect 4445 20009 4479 20043
rect 4479 20009 4488 20043
rect 4436 20000 4488 20009
rect 4896 20043 4948 20052
rect 4896 20009 4905 20043
rect 4905 20009 4939 20043
rect 4939 20009 4948 20043
rect 4896 20000 4948 20009
rect 5448 20000 5500 20052
rect 2412 19864 2464 19916
rect 1584 19839 1636 19848
rect 1584 19805 1593 19839
rect 1593 19805 1627 19839
rect 1627 19805 1636 19839
rect 1584 19796 1636 19805
rect 4620 19864 4672 19916
rect 6000 20000 6052 20052
rect 6184 20000 6236 20052
rect 6920 20000 6972 20052
rect 3148 19728 3200 19780
rect 5264 19796 5316 19848
rect 5356 19839 5408 19848
rect 5356 19805 5365 19839
rect 5365 19805 5399 19839
rect 5399 19805 5408 19839
rect 5356 19796 5408 19805
rect 5632 19796 5684 19848
rect 5724 19839 5776 19848
rect 5724 19805 5733 19839
rect 5733 19805 5767 19839
rect 5767 19805 5776 19839
rect 5724 19796 5776 19805
rect 6184 19907 6236 19916
rect 6184 19873 6193 19907
rect 6193 19873 6227 19907
rect 6227 19873 6236 19907
rect 6184 19864 6236 19873
rect 6276 19907 6328 19916
rect 6276 19873 6285 19907
rect 6285 19873 6319 19907
rect 6319 19873 6328 19907
rect 6276 19864 6328 19873
rect 6552 19864 6604 19916
rect 8024 20043 8076 20052
rect 8024 20009 8033 20043
rect 8033 20009 8067 20043
rect 8067 20009 8076 20043
rect 8024 20000 8076 20009
rect 9956 20000 10008 20052
rect 10784 20000 10836 20052
rect 8300 19864 8352 19916
rect 9220 19907 9272 19916
rect 9220 19873 9229 19907
rect 9229 19873 9263 19907
rect 9263 19873 9272 19907
rect 9220 19864 9272 19873
rect 8116 19796 8168 19848
rect 8760 19839 8812 19848
rect 8760 19805 8769 19839
rect 8769 19805 8803 19839
rect 8803 19805 8812 19839
rect 8760 19796 8812 19805
rect 11612 20000 11664 20052
rect 12900 20000 12952 20052
rect 15844 20000 15896 20052
rect 18604 20000 18656 20052
rect 23388 20000 23440 20052
rect 24492 20000 24544 20052
rect 12440 19864 12492 19916
rect 13360 19932 13412 19984
rect 17868 19907 17920 19916
rect 17868 19873 17877 19907
rect 17877 19873 17911 19907
rect 17911 19873 17920 19907
rect 17868 19864 17920 19873
rect 10968 19796 11020 19848
rect 12532 19796 12584 19848
rect 12900 19796 12952 19848
rect 13268 19796 13320 19848
rect 16488 19796 16540 19848
rect 18788 19796 18840 19848
rect 22652 19864 22704 19916
rect 22100 19796 22152 19848
rect 23020 19796 23072 19848
rect 23480 19796 23532 19848
rect 23848 19796 23900 19848
rect 24492 19796 24544 19848
rect 24768 19796 24820 19848
rect 25228 19839 25280 19848
rect 25228 19805 25237 19839
rect 25237 19805 25271 19839
rect 25271 19805 25280 19839
rect 25228 19796 25280 19805
rect 5816 19771 5868 19780
rect 5816 19737 5825 19771
rect 5825 19737 5859 19771
rect 5859 19737 5868 19771
rect 5816 19728 5868 19737
rect 6460 19728 6512 19780
rect 4804 19660 4856 19712
rect 5172 19660 5224 19712
rect 7012 19728 7064 19780
rect 8576 19703 8628 19712
rect 8576 19669 8585 19703
rect 8585 19669 8619 19703
rect 8619 19669 8628 19703
rect 8576 19660 8628 19669
rect 11152 19660 11204 19712
rect 12808 19660 12860 19712
rect 16304 19703 16356 19712
rect 16304 19669 16313 19703
rect 16313 19669 16347 19703
rect 16347 19669 16356 19703
rect 16304 19660 16356 19669
rect 17316 19703 17368 19712
rect 17316 19669 17325 19703
rect 17325 19669 17359 19703
rect 17359 19669 17368 19703
rect 17316 19660 17368 19669
rect 17684 19703 17736 19712
rect 17684 19669 17693 19703
rect 17693 19669 17727 19703
rect 17727 19669 17736 19703
rect 17684 19660 17736 19669
rect 20720 19703 20772 19712
rect 20720 19669 20729 19703
rect 20729 19669 20763 19703
rect 20763 19669 20772 19703
rect 20720 19660 20772 19669
rect 23848 19660 23900 19712
rect 24124 19660 24176 19712
rect 25412 19703 25464 19712
rect 25412 19669 25421 19703
rect 25421 19669 25455 19703
rect 25455 19669 25464 19703
rect 25412 19660 25464 19669
rect 7252 19558 7304 19610
rect 7316 19558 7368 19610
rect 7380 19558 7432 19610
rect 7444 19558 7496 19610
rect 7508 19558 7560 19610
rect 13554 19558 13606 19610
rect 13618 19558 13670 19610
rect 13682 19558 13734 19610
rect 13746 19558 13798 19610
rect 13810 19558 13862 19610
rect 19856 19558 19908 19610
rect 19920 19558 19972 19610
rect 19984 19558 20036 19610
rect 20048 19558 20100 19610
rect 20112 19558 20164 19610
rect 26158 19558 26210 19610
rect 26222 19558 26274 19610
rect 26286 19558 26338 19610
rect 26350 19558 26402 19610
rect 26414 19558 26466 19610
rect 2688 19456 2740 19508
rect 2780 19456 2832 19508
rect 2136 19388 2188 19440
rect 3332 19388 3384 19440
rect 4620 19456 4672 19508
rect 5356 19456 5408 19508
rect 5816 19456 5868 19508
rect 3976 19388 4028 19440
rect 1584 19363 1636 19372
rect 1584 19329 1593 19363
rect 1593 19329 1627 19363
rect 1627 19329 1636 19363
rect 1584 19320 1636 19329
rect 3148 19320 3200 19372
rect 5172 19320 5224 19372
rect 5632 19363 5684 19372
rect 5632 19329 5641 19363
rect 5641 19329 5675 19363
rect 5675 19329 5684 19363
rect 5632 19320 5684 19329
rect 6092 19456 6144 19508
rect 6460 19456 6512 19508
rect 6184 19363 6236 19372
rect 6184 19329 6193 19363
rect 6193 19329 6227 19363
rect 6227 19329 6236 19363
rect 6184 19320 6236 19329
rect 6368 19363 6420 19372
rect 6368 19329 6377 19363
rect 6377 19329 6411 19363
rect 6411 19329 6420 19363
rect 6368 19320 6420 19329
rect 8576 19388 8628 19440
rect 9680 19388 9732 19440
rect 8024 19320 8076 19372
rect 8300 19320 8352 19372
rect 11152 19363 11204 19372
rect 11152 19329 11161 19363
rect 11161 19329 11195 19363
rect 11195 19329 11204 19363
rect 11152 19320 11204 19329
rect 12440 19456 12492 19508
rect 16488 19499 16540 19508
rect 16488 19465 16497 19499
rect 16497 19465 16531 19499
rect 16531 19465 16540 19499
rect 16488 19456 16540 19465
rect 16580 19456 16632 19508
rect 17316 19456 17368 19508
rect 17776 19456 17828 19508
rect 18420 19456 18472 19508
rect 22100 19456 22152 19508
rect 24032 19456 24084 19508
rect 15476 19388 15528 19440
rect 12900 19320 12952 19372
rect 14740 19363 14792 19372
rect 14740 19329 14749 19363
rect 14749 19329 14783 19363
rect 14783 19329 14792 19363
rect 14740 19320 14792 19329
rect 9404 19252 9456 19304
rect 10324 19252 10376 19304
rect 12164 19252 12216 19304
rect 14648 19252 14700 19304
rect 15108 19252 15160 19304
rect 22836 19431 22888 19440
rect 22836 19397 22845 19431
rect 22845 19397 22879 19431
rect 22879 19397 22888 19431
rect 22836 19388 22888 19397
rect 21272 19320 21324 19372
rect 21916 19320 21968 19372
rect 22744 19320 22796 19372
rect 23020 19320 23072 19372
rect 23664 19320 23716 19372
rect 25228 19320 25280 19372
rect 17132 19295 17184 19304
rect 17132 19261 17141 19295
rect 17141 19261 17175 19295
rect 17175 19261 17184 19295
rect 17132 19252 17184 19261
rect 6000 19116 6052 19168
rect 10232 19159 10284 19168
rect 10232 19125 10241 19159
rect 10241 19125 10275 19159
rect 10275 19125 10284 19159
rect 10232 19116 10284 19125
rect 13268 19227 13320 19236
rect 13268 19193 13277 19227
rect 13277 19193 13311 19227
rect 13311 19193 13320 19227
rect 13268 19184 13320 19193
rect 18880 19252 18932 19304
rect 12164 19116 12216 19168
rect 12256 19116 12308 19168
rect 16948 19116 17000 19168
rect 18144 19116 18196 19168
rect 18788 19116 18840 19168
rect 19616 19116 19668 19168
rect 20720 19252 20772 19304
rect 22008 19252 22060 19304
rect 23480 19295 23532 19304
rect 23480 19261 23489 19295
rect 23489 19261 23523 19295
rect 23523 19261 23532 19295
rect 23480 19252 23532 19261
rect 24492 19252 24544 19304
rect 20720 19116 20772 19168
rect 22100 19116 22152 19168
rect 23664 19159 23716 19168
rect 23664 19125 23673 19159
rect 23673 19125 23707 19159
rect 23707 19125 23716 19159
rect 23664 19116 23716 19125
rect 4101 19014 4153 19066
rect 4165 19014 4217 19066
rect 4229 19014 4281 19066
rect 4293 19014 4345 19066
rect 4357 19014 4409 19066
rect 10403 19014 10455 19066
rect 10467 19014 10519 19066
rect 10531 19014 10583 19066
rect 10595 19014 10647 19066
rect 10659 19014 10711 19066
rect 16705 19014 16757 19066
rect 16769 19014 16821 19066
rect 16833 19014 16885 19066
rect 16897 19014 16949 19066
rect 16961 19014 17013 19066
rect 23007 19014 23059 19066
rect 23071 19014 23123 19066
rect 23135 19014 23187 19066
rect 23199 19014 23251 19066
rect 23263 19014 23315 19066
rect 5172 18955 5224 18964
rect 5172 18921 5181 18955
rect 5181 18921 5215 18955
rect 5215 18921 5224 18955
rect 5172 18912 5224 18921
rect 5632 18912 5684 18964
rect 8760 18912 8812 18964
rect 10784 18912 10836 18964
rect 10876 18912 10928 18964
rect 1584 18819 1636 18828
rect 1584 18785 1593 18819
rect 1593 18785 1627 18819
rect 1627 18785 1636 18819
rect 1584 18776 1636 18785
rect 6000 18819 6052 18828
rect 4160 18708 4212 18760
rect 4988 18708 5040 18760
rect 6000 18785 6009 18819
rect 6009 18785 6043 18819
rect 6043 18785 6052 18819
rect 6000 18776 6052 18785
rect 9404 18776 9456 18828
rect 1860 18683 1912 18692
rect 1860 18649 1869 18683
rect 1869 18649 1903 18683
rect 1903 18649 1912 18683
rect 1860 18640 1912 18649
rect 3240 18640 3292 18692
rect 5632 18751 5684 18760
rect 5632 18717 5641 18751
rect 5641 18717 5675 18751
rect 5675 18717 5684 18751
rect 5632 18708 5684 18717
rect 5816 18751 5868 18760
rect 5816 18717 5825 18751
rect 5825 18717 5859 18751
rect 5859 18717 5868 18751
rect 5816 18708 5868 18717
rect 10232 18708 10284 18760
rect 10324 18708 10376 18760
rect 9956 18640 10008 18692
rect 6184 18572 6236 18624
rect 10232 18572 10284 18624
rect 10784 18751 10836 18760
rect 10784 18717 10793 18751
rect 10793 18717 10827 18751
rect 10827 18717 10836 18751
rect 12532 18887 12584 18896
rect 12532 18853 12541 18887
rect 12541 18853 12575 18887
rect 12575 18853 12584 18887
rect 12532 18844 12584 18853
rect 15108 18912 15160 18964
rect 15384 18844 15436 18896
rect 15568 18887 15620 18896
rect 15568 18853 15577 18887
rect 15577 18853 15611 18887
rect 15611 18853 15620 18887
rect 15568 18844 15620 18853
rect 10784 18708 10836 18717
rect 13268 18776 13320 18828
rect 16212 18912 16264 18964
rect 12716 18708 12768 18760
rect 15016 18751 15068 18760
rect 15016 18717 15025 18751
rect 15025 18717 15059 18751
rect 15059 18717 15068 18751
rect 15016 18708 15068 18717
rect 15384 18751 15436 18760
rect 15384 18717 15393 18751
rect 15393 18717 15427 18751
rect 15427 18717 15436 18751
rect 16212 18819 16264 18828
rect 16212 18785 16221 18819
rect 16221 18785 16255 18819
rect 16255 18785 16264 18819
rect 16212 18776 16264 18785
rect 15384 18708 15436 18717
rect 16304 18708 16356 18760
rect 16488 18751 16540 18760
rect 16488 18717 16497 18751
rect 16497 18717 16531 18751
rect 16531 18717 16540 18751
rect 16488 18708 16540 18717
rect 19340 18912 19392 18964
rect 23480 18912 23532 18964
rect 18512 18844 18564 18896
rect 17132 18819 17184 18828
rect 17132 18785 17141 18819
rect 17141 18785 17175 18819
rect 17175 18785 17184 18819
rect 17132 18776 17184 18785
rect 17776 18776 17828 18828
rect 20720 18776 20772 18828
rect 22008 18776 22060 18828
rect 23664 18776 23716 18828
rect 19616 18751 19668 18760
rect 19616 18717 19625 18751
rect 19625 18717 19659 18751
rect 19659 18717 19668 18751
rect 19616 18708 19668 18717
rect 25228 18708 25280 18760
rect 12164 18683 12216 18692
rect 12164 18649 12173 18683
rect 12173 18649 12207 18683
rect 12207 18649 12216 18683
rect 12164 18640 12216 18649
rect 12808 18640 12860 18692
rect 10600 18572 10652 18624
rect 15292 18683 15344 18692
rect 15292 18649 15301 18683
rect 15301 18649 15335 18683
rect 15335 18649 15344 18683
rect 15292 18640 15344 18649
rect 15568 18640 15620 18692
rect 16580 18640 16632 18692
rect 16672 18683 16724 18692
rect 16672 18649 16681 18683
rect 16681 18649 16715 18683
rect 16715 18649 16724 18683
rect 16672 18640 16724 18649
rect 15936 18572 15988 18624
rect 16120 18615 16172 18624
rect 16120 18581 16129 18615
rect 16129 18581 16163 18615
rect 16163 18581 16172 18615
rect 16120 18572 16172 18581
rect 17040 18615 17092 18624
rect 17040 18581 17049 18615
rect 17049 18581 17083 18615
rect 17083 18581 17092 18615
rect 17040 18572 17092 18581
rect 17408 18683 17460 18692
rect 17408 18649 17417 18683
rect 17417 18649 17451 18683
rect 17451 18649 17460 18683
rect 17408 18640 17460 18649
rect 18420 18640 18472 18692
rect 20996 18640 21048 18692
rect 18144 18572 18196 18624
rect 18880 18615 18932 18624
rect 18880 18581 18889 18615
rect 18889 18581 18923 18615
rect 18923 18581 18932 18615
rect 18880 18572 18932 18581
rect 19248 18615 19300 18624
rect 19248 18581 19257 18615
rect 19257 18581 19291 18615
rect 19291 18581 19300 18615
rect 19248 18572 19300 18581
rect 22008 18572 22060 18624
rect 24492 18615 24544 18624
rect 24492 18581 24501 18615
rect 24501 18581 24535 18615
rect 24535 18581 24544 18615
rect 24492 18572 24544 18581
rect 7252 18470 7304 18522
rect 7316 18470 7368 18522
rect 7380 18470 7432 18522
rect 7444 18470 7496 18522
rect 7508 18470 7560 18522
rect 13554 18470 13606 18522
rect 13618 18470 13670 18522
rect 13682 18470 13734 18522
rect 13746 18470 13798 18522
rect 13810 18470 13862 18522
rect 19856 18470 19908 18522
rect 19920 18470 19972 18522
rect 19984 18470 20036 18522
rect 20048 18470 20100 18522
rect 20112 18470 20164 18522
rect 26158 18470 26210 18522
rect 26222 18470 26274 18522
rect 26286 18470 26338 18522
rect 26350 18470 26402 18522
rect 26414 18470 26466 18522
rect 1860 18368 1912 18420
rect 3516 18411 3568 18420
rect 3516 18377 3525 18411
rect 3525 18377 3559 18411
rect 3559 18377 3568 18411
rect 3516 18368 3568 18377
rect 4160 18368 4212 18420
rect 6920 18411 6972 18420
rect 6920 18377 6929 18411
rect 6929 18377 6963 18411
rect 6963 18377 6972 18411
rect 6920 18368 6972 18377
rect 8208 18368 8260 18420
rect 3516 18232 3568 18284
rect 4620 18232 4672 18284
rect 5908 18232 5960 18284
rect 6368 18232 6420 18284
rect 6828 18232 6880 18284
rect 9680 18300 9732 18352
rect 9496 18232 9548 18284
rect 16120 18368 16172 18420
rect 17408 18411 17460 18420
rect 17408 18377 17417 18411
rect 17417 18377 17451 18411
rect 17451 18377 17460 18411
rect 17408 18368 17460 18377
rect 10600 18343 10652 18352
rect 10600 18309 10609 18343
rect 10609 18309 10643 18343
rect 10643 18309 10652 18343
rect 10600 18300 10652 18309
rect 12164 18300 12216 18352
rect 3332 18207 3384 18216
rect 3332 18173 3341 18207
rect 3341 18173 3375 18207
rect 3375 18173 3384 18207
rect 3332 18164 3384 18173
rect 3976 18164 4028 18216
rect 4436 18164 4488 18216
rect 6184 18164 6236 18216
rect 6460 18207 6512 18216
rect 6460 18173 6469 18207
rect 6469 18173 6503 18207
rect 6503 18173 6512 18207
rect 6460 18164 6512 18173
rect 1952 18096 2004 18148
rect 8024 18207 8076 18216
rect 8024 18173 8033 18207
rect 8033 18173 8067 18207
rect 8067 18173 8076 18207
rect 8024 18164 8076 18173
rect 10140 18164 10192 18216
rect 10784 18275 10836 18284
rect 10784 18241 10793 18275
rect 10793 18241 10827 18275
rect 10827 18241 10836 18275
rect 10784 18232 10836 18241
rect 10876 18232 10928 18284
rect 15476 18300 15528 18352
rect 15936 18300 15988 18352
rect 16672 18300 16724 18352
rect 17776 18300 17828 18352
rect 5540 18071 5592 18080
rect 5540 18037 5549 18071
rect 5549 18037 5583 18071
rect 5583 18037 5592 18071
rect 5540 18028 5592 18037
rect 12624 18275 12676 18284
rect 12624 18241 12633 18275
rect 12633 18241 12667 18275
rect 12667 18241 12676 18275
rect 12624 18232 12676 18241
rect 12716 18275 12768 18284
rect 12716 18241 12730 18275
rect 12730 18241 12764 18275
rect 12764 18241 12768 18275
rect 12716 18232 12768 18241
rect 15292 18232 15344 18284
rect 15844 18275 15896 18284
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 15844 18232 15896 18241
rect 19248 18368 19300 18420
rect 20996 18411 21048 18420
rect 20996 18377 21005 18411
rect 21005 18377 21039 18411
rect 21039 18377 21048 18411
rect 20996 18368 21048 18377
rect 18420 18232 18472 18284
rect 24492 18368 24544 18420
rect 22100 18300 22152 18352
rect 23756 18300 23808 18352
rect 8484 18028 8536 18080
rect 9680 18071 9732 18080
rect 9680 18037 9689 18071
rect 9689 18037 9723 18071
rect 9723 18037 9732 18071
rect 9680 18028 9732 18037
rect 12440 18028 12492 18080
rect 12808 18028 12860 18080
rect 13360 18207 13412 18216
rect 13360 18173 13369 18207
rect 13369 18173 13403 18207
rect 13403 18173 13412 18207
rect 13360 18164 13412 18173
rect 13636 18207 13688 18216
rect 13636 18173 13645 18207
rect 13645 18173 13679 18207
rect 13679 18173 13688 18207
rect 13636 18164 13688 18173
rect 15016 18164 15068 18216
rect 17684 18164 17736 18216
rect 18144 18164 18196 18216
rect 21364 18232 21416 18284
rect 21916 18232 21968 18284
rect 14832 18096 14884 18148
rect 15476 18096 15528 18148
rect 19524 18207 19576 18216
rect 19524 18173 19533 18207
rect 19533 18173 19567 18207
rect 19567 18173 19576 18207
rect 19524 18164 19576 18173
rect 20720 18164 20772 18216
rect 22652 18164 22704 18216
rect 22836 18164 22888 18216
rect 24860 18164 24912 18216
rect 13452 18028 13504 18080
rect 15292 18071 15344 18080
rect 15292 18037 15301 18071
rect 15301 18037 15335 18071
rect 15335 18037 15344 18071
rect 15292 18028 15344 18037
rect 16580 18028 16632 18080
rect 18052 18071 18104 18080
rect 18052 18037 18061 18071
rect 18061 18037 18095 18071
rect 18095 18037 18104 18071
rect 18052 18028 18104 18037
rect 19892 18071 19944 18080
rect 19892 18037 19901 18071
rect 19901 18037 19935 18071
rect 19935 18037 19944 18071
rect 19892 18028 19944 18037
rect 22100 18028 22152 18080
rect 4101 17926 4153 17978
rect 4165 17926 4217 17978
rect 4229 17926 4281 17978
rect 4293 17926 4345 17978
rect 4357 17926 4409 17978
rect 10403 17926 10455 17978
rect 10467 17926 10519 17978
rect 10531 17926 10583 17978
rect 10595 17926 10647 17978
rect 10659 17926 10711 17978
rect 16705 17926 16757 17978
rect 16769 17926 16821 17978
rect 16833 17926 16885 17978
rect 16897 17926 16949 17978
rect 16961 17926 17013 17978
rect 23007 17926 23059 17978
rect 23071 17926 23123 17978
rect 23135 17926 23187 17978
rect 23199 17926 23251 17978
rect 23263 17926 23315 17978
rect 6092 17824 6144 17876
rect 6460 17824 6512 17876
rect 8024 17824 8076 17876
rect 9772 17824 9824 17876
rect 6368 17756 6420 17808
rect 6552 17756 6604 17808
rect 6736 17756 6788 17808
rect 5632 17688 5684 17740
rect 3516 17620 3568 17672
rect 4528 17620 4580 17672
rect 4988 17663 5040 17672
rect 4988 17629 4997 17663
rect 4997 17629 5031 17663
rect 5031 17629 5040 17663
rect 4988 17620 5040 17629
rect 5264 17663 5316 17672
rect 5264 17629 5273 17663
rect 5273 17629 5307 17663
rect 5307 17629 5316 17663
rect 5264 17620 5316 17629
rect 5356 17663 5408 17672
rect 5356 17629 5365 17663
rect 5365 17629 5399 17663
rect 5399 17629 5408 17663
rect 5356 17620 5408 17629
rect 5724 17620 5776 17672
rect 6000 17663 6052 17672
rect 6000 17629 6009 17663
rect 6009 17629 6043 17663
rect 6043 17629 6052 17663
rect 6000 17620 6052 17629
rect 6276 17620 6328 17672
rect 6368 17663 6420 17672
rect 6368 17629 6377 17663
rect 6377 17629 6411 17663
rect 6411 17629 6420 17663
rect 6368 17620 6420 17629
rect 6552 17663 6604 17672
rect 6552 17629 6561 17663
rect 6561 17629 6595 17663
rect 6595 17629 6604 17663
rect 6552 17620 6604 17629
rect 7104 17620 7156 17672
rect 11796 17756 11848 17808
rect 8116 17688 8168 17740
rect 12256 17688 12308 17740
rect 9680 17620 9732 17672
rect 10876 17663 10928 17672
rect 10876 17629 10885 17663
rect 10885 17629 10919 17663
rect 10919 17629 10928 17663
rect 10876 17620 10928 17629
rect 13636 17867 13688 17876
rect 13636 17833 13645 17867
rect 13645 17833 13679 17867
rect 13679 17833 13688 17867
rect 13636 17824 13688 17833
rect 15844 17867 15896 17876
rect 15844 17833 15853 17867
rect 15853 17833 15887 17867
rect 15887 17833 15896 17867
rect 15844 17824 15896 17833
rect 12624 17688 12676 17740
rect 13176 17731 13228 17740
rect 13176 17697 13185 17731
rect 13185 17697 13219 17731
rect 13219 17697 13228 17731
rect 13176 17688 13228 17697
rect 13360 17688 13412 17740
rect 14740 17688 14792 17740
rect 15016 17688 15068 17740
rect 16212 17688 16264 17740
rect 5172 17484 5224 17536
rect 6644 17484 6696 17536
rect 7932 17484 7984 17536
rect 10232 17527 10284 17536
rect 10232 17493 10241 17527
rect 10241 17493 10275 17527
rect 10275 17493 10284 17527
rect 10232 17484 10284 17493
rect 11520 17484 11572 17536
rect 14004 17620 14056 17672
rect 15476 17620 15528 17672
rect 16580 17620 16632 17672
rect 13452 17484 13504 17536
rect 18328 17824 18380 17876
rect 19524 17824 19576 17876
rect 17040 17663 17092 17672
rect 17040 17629 17049 17663
rect 17049 17629 17083 17663
rect 17083 17629 17092 17663
rect 17040 17620 17092 17629
rect 18880 17756 18932 17808
rect 22192 17824 22244 17876
rect 22376 17824 22428 17876
rect 22652 17824 22704 17876
rect 17408 17688 17460 17740
rect 17500 17663 17552 17672
rect 17500 17629 17514 17663
rect 17514 17629 17548 17663
rect 17548 17629 17552 17663
rect 17500 17620 17552 17629
rect 18052 17620 18104 17672
rect 20812 17688 20864 17740
rect 23756 17867 23808 17876
rect 23756 17833 23765 17867
rect 23765 17833 23799 17867
rect 23799 17833 23808 17867
rect 23756 17824 23808 17833
rect 24124 17824 24176 17876
rect 16396 17527 16448 17536
rect 16396 17493 16405 17527
rect 16405 17493 16439 17527
rect 16439 17493 16448 17527
rect 16396 17484 16448 17493
rect 17960 17484 18012 17536
rect 18144 17484 18196 17536
rect 19892 17620 19944 17672
rect 21732 17620 21784 17672
rect 22100 17620 22152 17672
rect 20904 17552 20956 17604
rect 22468 17663 22520 17672
rect 22468 17629 22477 17663
rect 22477 17629 22511 17663
rect 22511 17629 22520 17663
rect 22468 17620 22520 17629
rect 22652 17663 22704 17672
rect 22652 17629 22661 17663
rect 22661 17629 22695 17663
rect 22695 17629 22704 17663
rect 22652 17620 22704 17629
rect 22836 17663 22888 17672
rect 22836 17629 22845 17663
rect 22845 17629 22879 17663
rect 22879 17629 22888 17663
rect 22836 17620 22888 17629
rect 25412 17688 25464 17740
rect 23388 17620 23440 17672
rect 23940 17620 23992 17672
rect 22192 17484 22244 17536
rect 23664 17484 23716 17536
rect 7252 17382 7304 17434
rect 7316 17382 7368 17434
rect 7380 17382 7432 17434
rect 7444 17382 7496 17434
rect 7508 17382 7560 17434
rect 13554 17382 13606 17434
rect 13618 17382 13670 17434
rect 13682 17382 13734 17434
rect 13746 17382 13798 17434
rect 13810 17382 13862 17434
rect 19856 17382 19908 17434
rect 19920 17382 19972 17434
rect 19984 17382 20036 17434
rect 20048 17382 20100 17434
rect 20112 17382 20164 17434
rect 26158 17382 26210 17434
rect 26222 17382 26274 17434
rect 26286 17382 26338 17434
rect 26350 17382 26402 17434
rect 26414 17382 26466 17434
rect 5356 17280 5408 17332
rect 6368 17280 6420 17332
rect 10232 17280 10284 17332
rect 3240 17144 3292 17196
rect 1584 17119 1636 17128
rect 1584 17085 1593 17119
rect 1593 17085 1627 17119
rect 1627 17085 1636 17119
rect 1584 17076 1636 17085
rect 1860 17119 1912 17128
rect 1860 17085 1869 17119
rect 1869 17085 1903 17119
rect 1903 17085 1912 17119
rect 1860 17076 1912 17085
rect 6552 17255 6604 17264
rect 6552 17221 6561 17255
rect 6561 17221 6595 17255
rect 6595 17221 6604 17255
rect 6552 17212 6604 17221
rect 9588 17212 9640 17264
rect 11520 17280 11572 17332
rect 12716 17280 12768 17332
rect 4988 17187 5040 17196
rect 4988 17153 4997 17187
rect 4997 17153 5031 17187
rect 5031 17153 5040 17187
rect 4988 17144 5040 17153
rect 5172 17144 5224 17196
rect 5356 17187 5408 17196
rect 5356 17153 5365 17187
rect 5365 17153 5399 17187
rect 5399 17153 5408 17187
rect 5356 17144 5408 17153
rect 5448 17144 5500 17196
rect 5540 17187 5592 17196
rect 5540 17153 5549 17187
rect 5549 17153 5583 17187
rect 5583 17153 5592 17187
rect 5540 17144 5592 17153
rect 6276 17144 6328 17196
rect 6368 17187 6420 17196
rect 6368 17153 6377 17187
rect 6377 17153 6411 17187
rect 6411 17153 6420 17187
rect 6368 17144 6420 17153
rect 4712 17076 4764 17128
rect 5816 17076 5868 17128
rect 4804 17008 4856 17060
rect 6644 17076 6696 17128
rect 7012 17144 7064 17196
rect 9036 17187 9088 17196
rect 9036 17153 9045 17187
rect 9045 17153 9079 17187
rect 9079 17153 9088 17187
rect 9036 17144 9088 17153
rect 7104 17111 7156 17128
rect 7104 17077 7113 17111
rect 7113 17077 7147 17111
rect 7147 17077 7156 17111
rect 7104 17076 7156 17077
rect 9772 17076 9824 17128
rect 6276 17008 6328 17060
rect 6828 17008 6880 17060
rect 8760 17008 8812 17060
rect 11152 17144 11204 17196
rect 11888 17212 11940 17264
rect 13176 17280 13228 17332
rect 14004 17280 14056 17332
rect 15292 17280 15344 17332
rect 16396 17212 16448 17264
rect 12900 17144 12952 17196
rect 14004 17144 14056 17196
rect 18512 17280 18564 17332
rect 18788 17212 18840 17264
rect 22468 17280 22520 17332
rect 11796 17119 11848 17128
rect 11796 17085 11805 17119
rect 11805 17085 11839 17119
rect 11839 17085 11848 17119
rect 11796 17076 11848 17085
rect 11888 17076 11940 17128
rect 4988 16940 5040 16992
rect 6092 16940 6144 16992
rect 6184 16983 6236 16992
rect 6184 16949 6193 16983
rect 6193 16949 6227 16983
rect 6227 16949 6236 16983
rect 6184 16940 6236 16949
rect 6460 16940 6512 16992
rect 8852 16983 8904 16992
rect 8852 16949 8861 16983
rect 8861 16949 8895 16983
rect 8895 16949 8904 16983
rect 8852 16940 8904 16949
rect 10324 16940 10376 16992
rect 10784 16940 10836 16992
rect 12900 17008 12952 17060
rect 13360 17076 13412 17128
rect 13452 17076 13504 17128
rect 15108 17008 15160 17060
rect 15292 17076 15344 17128
rect 18512 17187 18564 17196
rect 18512 17153 18521 17187
rect 18521 17153 18555 17187
rect 18555 17153 18564 17187
rect 18512 17144 18564 17153
rect 19064 17187 19116 17196
rect 19064 17153 19073 17187
rect 19073 17153 19107 17187
rect 19107 17153 19116 17187
rect 19064 17144 19116 17153
rect 19432 17144 19484 17196
rect 21364 17187 21416 17196
rect 21364 17153 21373 17187
rect 21373 17153 21407 17187
rect 21407 17153 21416 17187
rect 21364 17144 21416 17153
rect 21548 17187 21600 17196
rect 21548 17153 21557 17187
rect 21557 17153 21591 17187
rect 21591 17153 21600 17187
rect 21548 17144 21600 17153
rect 23940 17187 23992 17196
rect 23940 17153 23949 17187
rect 23949 17153 23983 17187
rect 23983 17153 23992 17187
rect 23940 17144 23992 17153
rect 24768 17144 24820 17196
rect 17040 17076 17092 17128
rect 17868 17076 17920 17128
rect 26332 17076 26384 17128
rect 17408 17008 17460 17060
rect 13268 16940 13320 16992
rect 15200 16983 15252 16992
rect 15200 16949 15209 16983
rect 15209 16949 15243 16983
rect 15243 16949 15252 16983
rect 15200 16940 15252 16949
rect 19708 16940 19760 16992
rect 19984 16983 20036 16992
rect 19984 16949 19993 16983
rect 19993 16949 20027 16983
rect 20027 16949 20036 16983
rect 19984 16940 20036 16949
rect 22100 16940 22152 16992
rect 25596 16940 25648 16992
rect 4101 16838 4153 16890
rect 4165 16838 4217 16890
rect 4229 16838 4281 16890
rect 4293 16838 4345 16890
rect 4357 16838 4409 16890
rect 10403 16838 10455 16890
rect 10467 16838 10519 16890
rect 10531 16838 10583 16890
rect 10595 16838 10647 16890
rect 10659 16838 10711 16890
rect 16705 16838 16757 16890
rect 16769 16838 16821 16890
rect 16833 16838 16885 16890
rect 16897 16838 16949 16890
rect 16961 16838 17013 16890
rect 23007 16838 23059 16890
rect 23071 16838 23123 16890
rect 23135 16838 23187 16890
rect 23199 16838 23251 16890
rect 23263 16838 23315 16890
rect 1860 16736 1912 16788
rect 5264 16736 5316 16788
rect 6092 16779 6144 16788
rect 6092 16745 6101 16779
rect 6101 16745 6135 16779
rect 6135 16745 6144 16779
rect 6092 16736 6144 16745
rect 10324 16736 10376 16788
rect 10876 16736 10928 16788
rect 11152 16736 11204 16788
rect 4712 16668 4764 16720
rect 5908 16668 5960 16720
rect 1492 16643 1544 16652
rect 1492 16609 1501 16643
rect 1501 16609 1535 16643
rect 1535 16609 1544 16643
rect 1492 16600 1544 16609
rect 3332 16643 3384 16652
rect 3332 16609 3341 16643
rect 3341 16609 3375 16643
rect 3375 16609 3384 16643
rect 3332 16600 3384 16609
rect 5356 16600 5408 16652
rect 6460 16600 6512 16652
rect 7656 16600 7708 16652
rect 8116 16600 8168 16652
rect 10784 16643 10836 16652
rect 10784 16609 10793 16643
rect 10793 16609 10827 16643
rect 10827 16609 10836 16643
rect 10784 16600 10836 16609
rect 2228 16464 2280 16516
rect 5172 16575 5224 16584
rect 5172 16541 5181 16575
rect 5181 16541 5215 16575
rect 5215 16541 5224 16575
rect 5172 16532 5224 16541
rect 5540 16532 5592 16584
rect 6368 16532 6420 16584
rect 6552 16575 6604 16584
rect 6552 16541 6561 16575
rect 6561 16541 6595 16575
rect 6595 16541 6604 16575
rect 6552 16532 6604 16541
rect 6736 16575 6788 16584
rect 6736 16541 6745 16575
rect 6745 16541 6779 16575
rect 6779 16541 6788 16575
rect 6736 16532 6788 16541
rect 8760 16532 8812 16584
rect 8944 16575 8996 16584
rect 8944 16541 8953 16575
rect 8953 16541 8987 16575
rect 8987 16541 8996 16575
rect 8944 16532 8996 16541
rect 12440 16736 12492 16788
rect 12900 16736 12952 16788
rect 13268 16736 13320 16788
rect 16396 16736 16448 16788
rect 15016 16643 15068 16652
rect 15016 16609 15025 16643
rect 15025 16609 15059 16643
rect 15059 16609 15068 16643
rect 15016 16600 15068 16609
rect 18512 16736 18564 16788
rect 19340 16779 19392 16788
rect 19340 16745 19349 16779
rect 19349 16745 19383 16779
rect 19383 16745 19392 16779
rect 19340 16736 19392 16745
rect 23940 16736 23992 16788
rect 3056 16439 3108 16448
rect 3056 16405 3065 16439
rect 3065 16405 3099 16439
rect 3099 16405 3108 16439
rect 3056 16396 3108 16405
rect 3608 16396 3660 16448
rect 4620 16507 4672 16516
rect 4620 16473 4629 16507
rect 4629 16473 4663 16507
rect 4663 16473 4672 16507
rect 4620 16464 4672 16473
rect 4712 16464 4764 16516
rect 6920 16464 6972 16516
rect 5632 16396 5684 16448
rect 6276 16396 6328 16448
rect 6368 16439 6420 16448
rect 6368 16405 6377 16439
rect 6377 16405 6411 16439
rect 6411 16405 6420 16439
rect 6368 16396 6420 16405
rect 9496 16464 9548 16516
rect 12072 16396 12124 16448
rect 12716 16464 12768 16516
rect 14740 16439 14792 16448
rect 14740 16405 14749 16439
rect 14749 16405 14783 16439
rect 14783 16405 14792 16439
rect 14740 16396 14792 16405
rect 14924 16575 14976 16584
rect 14924 16541 14933 16575
rect 14933 16541 14967 16575
rect 14967 16541 14976 16575
rect 14924 16532 14976 16541
rect 17408 16643 17460 16652
rect 17408 16609 17417 16643
rect 17417 16609 17451 16643
rect 17451 16609 17460 16643
rect 17408 16600 17460 16609
rect 17776 16600 17828 16652
rect 17040 16532 17092 16584
rect 18420 16600 18472 16652
rect 18512 16600 18564 16652
rect 20904 16600 20956 16652
rect 23480 16600 23532 16652
rect 18788 16532 18840 16584
rect 19340 16532 19392 16584
rect 15568 16464 15620 16516
rect 19708 16464 19760 16516
rect 19984 16464 20036 16516
rect 20812 16532 20864 16584
rect 20996 16464 21048 16516
rect 18880 16396 18932 16448
rect 21824 16575 21876 16584
rect 21824 16541 21833 16575
rect 21833 16541 21867 16575
rect 21867 16541 21876 16575
rect 21824 16532 21876 16541
rect 23572 16464 23624 16516
rect 23388 16396 23440 16448
rect 7252 16294 7304 16346
rect 7316 16294 7368 16346
rect 7380 16294 7432 16346
rect 7444 16294 7496 16346
rect 7508 16294 7560 16346
rect 13554 16294 13606 16346
rect 13618 16294 13670 16346
rect 13682 16294 13734 16346
rect 13746 16294 13798 16346
rect 13810 16294 13862 16346
rect 19856 16294 19908 16346
rect 19920 16294 19972 16346
rect 19984 16294 20036 16346
rect 20048 16294 20100 16346
rect 20112 16294 20164 16346
rect 26158 16294 26210 16346
rect 26222 16294 26274 16346
rect 26286 16294 26338 16346
rect 26350 16294 26402 16346
rect 26414 16294 26466 16346
rect 5632 16235 5684 16244
rect 5632 16201 5641 16235
rect 5641 16201 5675 16235
rect 5675 16201 5684 16235
rect 5632 16192 5684 16201
rect 6552 16192 6604 16244
rect 6920 16235 6972 16244
rect 6920 16201 6929 16235
rect 6929 16201 6963 16235
rect 6963 16201 6972 16235
rect 6920 16192 6972 16201
rect 3516 16124 3568 16176
rect 4988 16124 5040 16176
rect 9496 16192 9548 16244
rect 2504 16099 2556 16108
rect 2504 16065 2513 16099
rect 2513 16065 2547 16099
rect 2547 16065 2556 16099
rect 2504 16056 2556 16065
rect 3056 16099 3108 16108
rect 3056 16065 3065 16099
rect 3065 16065 3099 16099
rect 3099 16065 3108 16099
rect 3056 16056 3108 16065
rect 3332 15988 3384 16040
rect 5172 16056 5224 16108
rect 5264 16056 5316 16108
rect 5724 16056 5776 16108
rect 6276 16056 6328 16108
rect 6736 16056 6788 16108
rect 6920 16056 6972 16108
rect 8944 16124 8996 16176
rect 2044 15895 2096 15904
rect 2044 15861 2053 15895
rect 2053 15861 2087 15895
rect 2087 15861 2096 15895
rect 2044 15852 2096 15861
rect 2320 15895 2372 15904
rect 2320 15861 2329 15895
rect 2329 15861 2363 15895
rect 2363 15861 2372 15895
rect 2320 15852 2372 15861
rect 7012 15988 7064 16040
rect 7104 15988 7156 16040
rect 5356 15920 5408 15972
rect 6828 15920 6880 15972
rect 7840 15852 7892 15904
rect 8024 16031 8076 16040
rect 8024 15997 8033 16031
rect 8033 15997 8067 16031
rect 8067 15997 8076 16031
rect 8024 15988 8076 15997
rect 10140 16235 10192 16244
rect 10140 16201 10149 16235
rect 10149 16201 10183 16235
rect 10183 16201 10192 16235
rect 10140 16192 10192 16201
rect 14740 16192 14792 16244
rect 16948 16192 17000 16244
rect 17040 16192 17092 16244
rect 17224 16192 17276 16244
rect 15476 16124 15528 16176
rect 16580 16056 16632 16108
rect 21364 16192 21416 16244
rect 21824 16192 21876 16244
rect 24860 16192 24912 16244
rect 17868 16167 17920 16176
rect 17868 16133 17877 16167
rect 17877 16133 17911 16167
rect 17911 16133 17920 16167
rect 17868 16124 17920 16133
rect 19432 16124 19484 16176
rect 20720 16124 20772 16176
rect 14004 15988 14056 16040
rect 14096 15988 14148 16040
rect 14832 15988 14884 16040
rect 17500 16056 17552 16108
rect 18420 16099 18472 16108
rect 18420 16065 18429 16099
rect 18429 16065 18463 16099
rect 18463 16065 18472 16099
rect 18420 16056 18472 16065
rect 18880 16099 18932 16108
rect 18880 16065 18889 16099
rect 18889 16065 18923 16099
rect 18923 16065 18932 16099
rect 18880 16056 18932 16065
rect 19156 16097 19165 16108
rect 19165 16097 19199 16108
rect 19199 16097 19208 16108
rect 19156 16056 19208 16097
rect 18788 15988 18840 16040
rect 20628 16056 20680 16108
rect 19984 15920 20036 15972
rect 8024 15852 8076 15904
rect 8852 15852 8904 15904
rect 10232 15895 10284 15904
rect 10232 15861 10241 15895
rect 10241 15861 10275 15895
rect 10275 15861 10284 15895
rect 10232 15852 10284 15861
rect 17316 15895 17368 15904
rect 17316 15861 17325 15895
rect 17325 15861 17359 15895
rect 17359 15861 17368 15895
rect 17316 15852 17368 15861
rect 18328 15852 18380 15904
rect 18696 15852 18748 15904
rect 20444 15988 20496 16040
rect 22100 16167 22152 16176
rect 22100 16133 22109 16167
rect 22109 16133 22143 16167
rect 22143 16133 22152 16167
rect 22100 16124 22152 16133
rect 23388 16124 23440 16176
rect 25504 16167 25556 16176
rect 25504 16133 25513 16167
rect 25513 16133 25547 16167
rect 25547 16133 25556 16167
rect 25504 16124 25556 16133
rect 21732 15988 21784 16040
rect 23572 16056 23624 16108
rect 24492 16056 24544 16108
rect 25780 16031 25832 16040
rect 25780 15997 25789 16031
rect 25789 15997 25823 16031
rect 25823 15997 25832 16031
rect 25780 15988 25832 15997
rect 21824 15920 21876 15972
rect 21364 15852 21416 15904
rect 24032 15895 24084 15904
rect 24032 15861 24041 15895
rect 24041 15861 24075 15895
rect 24075 15861 24084 15895
rect 24032 15852 24084 15861
rect 4101 15750 4153 15802
rect 4165 15750 4217 15802
rect 4229 15750 4281 15802
rect 4293 15750 4345 15802
rect 4357 15750 4409 15802
rect 10403 15750 10455 15802
rect 10467 15750 10519 15802
rect 10531 15750 10583 15802
rect 10595 15750 10647 15802
rect 10659 15750 10711 15802
rect 16705 15750 16757 15802
rect 16769 15750 16821 15802
rect 16833 15750 16885 15802
rect 16897 15750 16949 15802
rect 16961 15750 17013 15802
rect 23007 15750 23059 15802
rect 23071 15750 23123 15802
rect 23135 15750 23187 15802
rect 23199 15750 23251 15802
rect 23263 15750 23315 15802
rect 2320 15648 2372 15700
rect 2504 15648 2556 15700
rect 4160 15648 4212 15700
rect 4712 15648 4764 15700
rect 6920 15691 6972 15700
rect 6920 15657 6929 15691
rect 6929 15657 6963 15691
rect 6963 15657 6972 15691
rect 6920 15648 6972 15657
rect 7012 15648 7064 15700
rect 8024 15648 8076 15700
rect 9036 15648 9088 15700
rect 10232 15648 10284 15700
rect 10324 15648 10376 15700
rect 11704 15648 11756 15700
rect 18144 15648 18196 15700
rect 19064 15648 19116 15700
rect 19340 15648 19392 15700
rect 21732 15648 21784 15700
rect 1584 15555 1636 15564
rect 1584 15521 1593 15555
rect 1593 15521 1627 15555
rect 1627 15521 1636 15555
rect 1584 15512 1636 15521
rect 2596 15512 2648 15564
rect 3240 15444 3292 15496
rect 3332 15444 3384 15496
rect 4068 15444 4120 15496
rect 4712 15512 4764 15564
rect 4988 15444 5040 15496
rect 7840 15512 7892 15564
rect 9404 15512 9456 15564
rect 3608 15419 3660 15428
rect 3608 15385 3617 15419
rect 3617 15385 3651 15419
rect 3651 15385 3660 15419
rect 3608 15376 3660 15385
rect 4344 15308 4396 15360
rect 4620 15308 4672 15360
rect 5908 15376 5960 15428
rect 6368 15308 6420 15360
rect 9496 15444 9548 15496
rect 19984 15623 20036 15632
rect 19984 15589 19993 15623
rect 19993 15589 20027 15623
rect 20027 15589 20036 15623
rect 19984 15580 20036 15589
rect 12348 15512 12400 15564
rect 17776 15512 17828 15564
rect 18420 15512 18472 15564
rect 11428 15444 11480 15496
rect 7196 15376 7248 15428
rect 8024 15308 8076 15360
rect 8852 15308 8904 15360
rect 9588 15308 9640 15360
rect 11336 15351 11388 15360
rect 11336 15317 11345 15351
rect 11345 15317 11379 15351
rect 11379 15317 11388 15351
rect 11336 15308 11388 15317
rect 11704 15351 11756 15360
rect 11704 15317 11713 15351
rect 11713 15317 11747 15351
rect 11747 15317 11756 15351
rect 11704 15308 11756 15317
rect 14188 15444 14240 15496
rect 16212 15444 16264 15496
rect 18512 15487 18564 15496
rect 18512 15453 18521 15487
rect 18521 15453 18555 15487
rect 18555 15453 18564 15487
rect 18512 15444 18564 15453
rect 18696 15444 18748 15496
rect 18880 15487 18932 15496
rect 18880 15453 18890 15487
rect 18890 15453 18924 15487
rect 18924 15453 18932 15487
rect 18880 15444 18932 15453
rect 19340 15444 19392 15496
rect 19432 15444 19484 15496
rect 20352 15487 20404 15496
rect 20352 15453 20361 15487
rect 20361 15453 20395 15487
rect 20395 15453 20404 15487
rect 20352 15444 20404 15453
rect 20444 15487 20496 15496
rect 20444 15453 20453 15487
rect 20453 15453 20487 15487
rect 20487 15453 20496 15487
rect 20444 15444 20496 15453
rect 21824 15444 21876 15496
rect 12532 15376 12584 15428
rect 13452 15308 13504 15360
rect 14372 15308 14424 15360
rect 17224 15308 17276 15360
rect 17684 15419 17736 15428
rect 17684 15385 17693 15419
rect 17693 15385 17727 15419
rect 17727 15385 17736 15419
rect 17684 15376 17736 15385
rect 17868 15419 17920 15428
rect 17868 15385 17877 15419
rect 17877 15385 17911 15419
rect 17911 15385 17920 15419
rect 17868 15376 17920 15385
rect 19156 15376 19208 15428
rect 20720 15419 20772 15428
rect 20720 15385 20729 15419
rect 20729 15385 20763 15419
rect 20763 15385 20772 15419
rect 20720 15376 20772 15385
rect 22560 15648 22612 15700
rect 23480 15691 23532 15700
rect 23480 15657 23489 15691
rect 23489 15657 23523 15691
rect 23523 15657 23532 15691
rect 23480 15648 23532 15657
rect 24032 15648 24084 15700
rect 22284 15555 22336 15564
rect 22284 15521 22293 15555
rect 22293 15521 22327 15555
rect 22327 15521 22336 15555
rect 22284 15512 22336 15521
rect 18236 15308 18288 15360
rect 18328 15308 18380 15360
rect 19432 15351 19484 15360
rect 19432 15317 19441 15351
rect 19441 15317 19475 15351
rect 19475 15317 19484 15351
rect 19432 15308 19484 15317
rect 19616 15308 19668 15360
rect 22928 15351 22980 15360
rect 22928 15317 22937 15351
rect 22937 15317 22971 15351
rect 22971 15317 22980 15351
rect 22928 15308 22980 15317
rect 23112 15308 23164 15360
rect 25228 15308 25280 15360
rect 7252 15206 7304 15258
rect 7316 15206 7368 15258
rect 7380 15206 7432 15258
rect 7444 15206 7496 15258
rect 7508 15206 7560 15258
rect 13554 15206 13606 15258
rect 13618 15206 13670 15258
rect 13682 15206 13734 15258
rect 13746 15206 13798 15258
rect 13810 15206 13862 15258
rect 19856 15206 19908 15258
rect 19920 15206 19972 15258
rect 19984 15206 20036 15258
rect 20048 15206 20100 15258
rect 20112 15206 20164 15258
rect 26158 15206 26210 15258
rect 26222 15206 26274 15258
rect 26286 15206 26338 15258
rect 26350 15206 26402 15258
rect 26414 15206 26466 15258
rect 2044 15104 2096 15156
rect 4068 15104 4120 15156
rect 4160 15147 4212 15156
rect 4160 15113 4169 15147
rect 4169 15113 4203 15147
rect 4203 15113 4212 15147
rect 4160 15104 4212 15113
rect 5724 15104 5776 15156
rect 6460 15147 6512 15156
rect 6460 15113 6469 15147
rect 6469 15113 6503 15147
rect 6503 15113 6512 15147
rect 6460 15104 6512 15113
rect 7104 15104 7156 15156
rect 3240 15036 3292 15088
rect 1584 15011 1636 15020
rect 1584 14977 1593 15011
rect 1593 14977 1627 15011
rect 1627 14977 1636 15011
rect 1584 14968 1636 14977
rect 3516 14968 3568 15020
rect 3976 14968 4028 15020
rect 7380 15036 7432 15088
rect 7656 15036 7708 15088
rect 6184 14968 6236 15020
rect 6552 14968 6604 15020
rect 7196 15011 7248 15020
rect 7196 14977 7205 15011
rect 7205 14977 7239 15011
rect 7239 14977 7248 15011
rect 7196 14968 7248 14977
rect 8852 15011 8904 15020
rect 8852 14977 8861 15011
rect 8861 14977 8895 15011
rect 8895 14977 8904 15011
rect 8852 14968 8904 14977
rect 11428 15104 11480 15156
rect 6736 14900 6788 14952
rect 11428 14968 11480 15020
rect 11704 15036 11756 15088
rect 12072 15036 12124 15088
rect 12256 15036 12308 15088
rect 14096 15036 14148 15088
rect 27068 15104 27120 15156
rect 16764 15036 16816 15088
rect 17776 15036 17828 15088
rect 18236 15036 18288 15088
rect 19156 15036 19208 15088
rect 4344 14832 4396 14884
rect 4804 14832 4856 14884
rect 11060 14900 11112 14952
rect 11244 14900 11296 14952
rect 12808 14900 12860 14952
rect 18144 14900 18196 14952
rect 20444 14968 20496 15020
rect 20996 14968 21048 15020
rect 24492 15036 24544 15088
rect 25228 15036 25280 15088
rect 21364 15011 21416 15020
rect 21364 14977 21373 15011
rect 21373 14977 21407 15011
rect 21407 14977 21416 15011
rect 21364 14968 21416 14977
rect 21548 14968 21600 15020
rect 23112 14968 23164 15020
rect 25780 15011 25832 15020
rect 25780 14977 25789 15011
rect 25789 14977 25823 15011
rect 25823 14977 25832 15011
rect 25780 14968 25832 14977
rect 19708 14943 19760 14952
rect 19708 14909 19717 14943
rect 19717 14909 19751 14943
rect 19751 14909 19760 14943
rect 19708 14900 19760 14909
rect 17684 14832 17736 14884
rect 3700 14807 3752 14816
rect 3700 14773 3709 14807
rect 3709 14773 3743 14807
rect 3743 14773 3752 14807
rect 3700 14764 3752 14773
rect 4896 14764 4948 14816
rect 9588 14764 9640 14816
rect 10140 14764 10192 14816
rect 13452 14764 13504 14816
rect 14004 14807 14056 14816
rect 14004 14773 14013 14807
rect 14013 14773 14047 14807
rect 14047 14773 14056 14807
rect 14004 14764 14056 14773
rect 17592 14764 17644 14816
rect 20720 14832 20772 14884
rect 21272 14943 21324 14952
rect 21272 14909 21281 14943
rect 21281 14909 21315 14943
rect 21315 14909 21324 14943
rect 21272 14900 21324 14909
rect 23388 14764 23440 14816
rect 25044 14764 25096 14816
rect 4101 14662 4153 14714
rect 4165 14662 4217 14714
rect 4229 14662 4281 14714
rect 4293 14662 4345 14714
rect 4357 14662 4409 14714
rect 10403 14662 10455 14714
rect 10467 14662 10519 14714
rect 10531 14662 10583 14714
rect 10595 14662 10647 14714
rect 10659 14662 10711 14714
rect 16705 14662 16757 14714
rect 16769 14662 16821 14714
rect 16833 14662 16885 14714
rect 16897 14662 16949 14714
rect 16961 14662 17013 14714
rect 23007 14662 23059 14714
rect 23071 14662 23123 14714
rect 23135 14662 23187 14714
rect 23199 14662 23251 14714
rect 23263 14662 23315 14714
rect 3700 14560 3752 14612
rect 6460 14560 6512 14612
rect 7196 14560 7248 14612
rect 3148 14399 3200 14408
rect 3148 14365 3157 14399
rect 3157 14365 3191 14399
rect 3191 14365 3200 14399
rect 3148 14356 3200 14365
rect 3976 14424 4028 14476
rect 6552 14467 6604 14476
rect 6552 14433 6561 14467
rect 6561 14433 6595 14467
rect 6595 14433 6604 14467
rect 6552 14424 6604 14433
rect 7748 14492 7800 14544
rect 8116 14492 8168 14544
rect 10692 14492 10744 14544
rect 6736 14467 6788 14476
rect 6736 14433 6745 14467
rect 6745 14433 6779 14467
rect 6779 14433 6788 14467
rect 6736 14424 6788 14433
rect 5908 14356 5960 14408
rect 6920 14356 6972 14408
rect 10600 14424 10652 14476
rect 11060 14560 11112 14612
rect 18144 14560 18196 14612
rect 12348 14492 12400 14544
rect 11336 14424 11388 14476
rect 11612 14424 11664 14476
rect 11980 14424 12032 14476
rect 14372 14467 14424 14476
rect 14372 14433 14381 14467
rect 14381 14433 14415 14467
rect 14415 14433 14424 14467
rect 14372 14424 14424 14433
rect 18236 14424 18288 14476
rect 18880 14492 18932 14544
rect 19616 14560 19668 14612
rect 19432 14492 19484 14544
rect 23296 14560 23348 14612
rect 23388 14603 23440 14612
rect 23388 14569 23397 14603
rect 23397 14569 23431 14603
rect 23431 14569 23440 14603
rect 23388 14560 23440 14569
rect 24584 14603 24636 14612
rect 24584 14569 24593 14603
rect 24593 14569 24627 14603
rect 24627 14569 24636 14603
rect 24584 14560 24636 14569
rect 20352 14467 20404 14476
rect 9956 14288 10008 14340
rect 3148 14220 3200 14272
rect 3332 14263 3384 14272
rect 3332 14229 3341 14263
rect 3341 14229 3375 14263
rect 3375 14229 3384 14263
rect 3332 14220 3384 14229
rect 8208 14220 8260 14272
rect 8300 14263 8352 14272
rect 8300 14229 8309 14263
rect 8309 14229 8343 14263
rect 8343 14229 8352 14263
rect 8300 14220 8352 14229
rect 9312 14220 9364 14272
rect 9864 14263 9916 14272
rect 9864 14229 9873 14263
rect 9873 14229 9907 14263
rect 9907 14229 9916 14263
rect 9864 14220 9916 14229
rect 10232 14356 10284 14408
rect 10416 14288 10468 14340
rect 10324 14220 10376 14272
rect 12256 14356 12308 14408
rect 14096 14399 14148 14408
rect 14096 14365 14105 14399
rect 14105 14365 14139 14399
rect 14139 14365 14148 14399
rect 14096 14356 14148 14365
rect 15476 14356 15528 14408
rect 20352 14433 20361 14467
rect 20361 14433 20395 14467
rect 20395 14433 20404 14467
rect 20352 14424 20404 14433
rect 21456 14424 21508 14476
rect 23480 14424 23532 14476
rect 11244 14288 11296 14340
rect 19156 14288 19208 14340
rect 21824 14331 21876 14340
rect 21824 14297 21833 14331
rect 21833 14297 21867 14331
rect 21867 14297 21876 14331
rect 21824 14288 21876 14297
rect 14464 14220 14516 14272
rect 19248 14263 19300 14272
rect 19248 14229 19257 14263
rect 19257 14229 19291 14263
rect 19291 14229 19300 14263
rect 19248 14220 19300 14229
rect 20260 14220 20312 14272
rect 21640 14220 21692 14272
rect 22468 14399 22520 14408
rect 22468 14365 22477 14399
rect 22477 14365 22511 14399
rect 22511 14365 22520 14399
rect 22468 14356 22520 14365
rect 22744 14356 22796 14408
rect 23204 14399 23256 14408
rect 23204 14365 23213 14399
rect 23213 14365 23247 14399
rect 23247 14365 23256 14399
rect 23204 14356 23256 14365
rect 24216 14356 24268 14408
rect 24676 14399 24728 14408
rect 24676 14365 24685 14399
rect 24685 14365 24719 14399
rect 24719 14365 24728 14399
rect 24676 14356 24728 14365
rect 25044 14399 25096 14408
rect 25044 14365 25053 14399
rect 25053 14365 25087 14399
rect 25087 14365 25096 14399
rect 25044 14356 25096 14365
rect 23296 14288 23348 14340
rect 23388 14220 23440 14272
rect 24952 14263 25004 14272
rect 24952 14229 24961 14263
rect 24961 14229 24995 14263
rect 24995 14229 25004 14263
rect 24952 14220 25004 14229
rect 25688 14263 25740 14272
rect 25688 14229 25697 14263
rect 25697 14229 25731 14263
rect 25731 14229 25740 14263
rect 25688 14220 25740 14229
rect 7252 14118 7304 14170
rect 7316 14118 7368 14170
rect 7380 14118 7432 14170
rect 7444 14118 7496 14170
rect 7508 14118 7560 14170
rect 13554 14118 13606 14170
rect 13618 14118 13670 14170
rect 13682 14118 13734 14170
rect 13746 14118 13798 14170
rect 13810 14118 13862 14170
rect 19856 14118 19908 14170
rect 19920 14118 19972 14170
rect 19984 14118 20036 14170
rect 20048 14118 20100 14170
rect 20112 14118 20164 14170
rect 26158 14118 26210 14170
rect 26222 14118 26274 14170
rect 26286 14118 26338 14170
rect 26350 14118 26402 14170
rect 26414 14118 26466 14170
rect 3332 13948 3384 14000
rect 2596 13880 2648 13932
rect 3148 13812 3200 13864
rect 4896 13880 4948 13932
rect 5080 13880 5132 13932
rect 4804 13855 4856 13864
rect 4804 13821 4813 13855
rect 4813 13821 4847 13855
rect 4847 13821 4856 13855
rect 4804 13812 4856 13821
rect 5632 13719 5684 13728
rect 5632 13685 5641 13719
rect 5641 13685 5675 13719
rect 5675 13685 5684 13719
rect 5632 13676 5684 13685
rect 6184 13923 6236 13932
rect 6184 13889 6193 13923
rect 6193 13889 6227 13923
rect 6227 13889 6236 13923
rect 6184 13880 6236 13889
rect 8300 14016 8352 14068
rect 8944 14016 8996 14068
rect 7748 13948 7800 14000
rect 9128 13948 9180 14000
rect 9312 13948 9364 14000
rect 6000 13744 6052 13796
rect 6920 13855 6972 13864
rect 6920 13821 6929 13855
rect 6929 13821 6963 13855
rect 6963 13821 6972 13855
rect 6920 13812 6972 13821
rect 7012 13855 7064 13864
rect 7012 13821 7021 13855
rect 7021 13821 7055 13855
rect 7055 13821 7064 13855
rect 7012 13812 7064 13821
rect 8208 13812 8260 13864
rect 10600 14016 10652 14068
rect 14188 14016 14240 14068
rect 14464 14059 14516 14068
rect 14464 14025 14473 14059
rect 14473 14025 14507 14059
rect 14507 14025 14516 14059
rect 14464 14016 14516 14025
rect 15844 14016 15896 14068
rect 9864 13991 9916 14000
rect 9864 13957 9873 13991
rect 9873 13957 9907 13991
rect 9907 13957 9916 13991
rect 9864 13948 9916 13957
rect 10140 13948 10192 14000
rect 11152 13948 11204 14000
rect 13912 13948 13964 14000
rect 7380 13676 7432 13728
rect 7932 13676 7984 13728
rect 9128 13676 9180 13728
rect 10232 13812 10284 13864
rect 10324 13812 10376 13864
rect 14280 13880 14332 13932
rect 17316 14016 17368 14068
rect 18328 13948 18380 14000
rect 17040 13923 17092 13932
rect 17040 13889 17049 13923
rect 17049 13889 17083 13923
rect 17083 13889 17092 13923
rect 17040 13880 17092 13889
rect 19156 13948 19208 14000
rect 19708 14016 19760 14068
rect 21824 14016 21876 14068
rect 20812 13948 20864 14000
rect 21456 13948 21508 14000
rect 21732 13948 21784 14000
rect 12348 13744 12400 13796
rect 17868 13744 17920 13796
rect 20444 13812 20496 13864
rect 21640 13923 21692 13932
rect 21640 13889 21649 13923
rect 21649 13889 21683 13923
rect 21683 13889 21692 13923
rect 21640 13880 21692 13889
rect 24584 14016 24636 14068
rect 21548 13812 21600 13864
rect 24032 13948 24084 14000
rect 25688 13948 25740 14000
rect 22192 13744 22244 13796
rect 22744 13880 22796 13932
rect 22836 13923 22888 13932
rect 22836 13889 22845 13923
rect 22845 13889 22879 13923
rect 22879 13889 22888 13923
rect 22836 13880 22888 13889
rect 23388 13880 23440 13932
rect 22468 13855 22520 13864
rect 22468 13821 22477 13855
rect 22477 13821 22511 13855
rect 22511 13821 22520 13855
rect 22468 13812 22520 13821
rect 23204 13812 23256 13864
rect 24400 13812 24452 13864
rect 25688 13855 25740 13864
rect 25688 13821 25697 13855
rect 25697 13821 25731 13855
rect 25731 13821 25740 13855
rect 25688 13812 25740 13821
rect 15016 13719 15068 13728
rect 15016 13685 15025 13719
rect 15025 13685 15059 13719
rect 15059 13685 15068 13719
rect 15016 13676 15068 13685
rect 16304 13676 16356 13728
rect 22468 13676 22520 13728
rect 22652 13676 22704 13728
rect 23388 13676 23440 13728
rect 25320 13676 25372 13728
rect 4101 13574 4153 13626
rect 4165 13574 4217 13626
rect 4229 13574 4281 13626
rect 4293 13574 4345 13626
rect 4357 13574 4409 13626
rect 10403 13574 10455 13626
rect 10467 13574 10519 13626
rect 10531 13574 10583 13626
rect 10595 13574 10647 13626
rect 10659 13574 10711 13626
rect 16705 13574 16757 13626
rect 16769 13574 16821 13626
rect 16833 13574 16885 13626
rect 16897 13574 16949 13626
rect 16961 13574 17013 13626
rect 23007 13574 23059 13626
rect 23071 13574 23123 13626
rect 23135 13574 23187 13626
rect 23199 13574 23251 13626
rect 23263 13574 23315 13626
rect 4988 13472 5040 13524
rect 5632 13472 5684 13524
rect 5724 13472 5776 13524
rect 6092 13472 6144 13524
rect 6368 13472 6420 13524
rect 6828 13515 6880 13524
rect 6828 13481 6837 13515
rect 6837 13481 6871 13515
rect 6871 13481 6880 13515
rect 6828 13472 6880 13481
rect 4344 13404 4396 13456
rect 6184 13404 6236 13456
rect 6460 13404 6512 13456
rect 11060 13472 11112 13524
rect 13912 13515 13964 13524
rect 13912 13481 13921 13515
rect 13921 13481 13955 13515
rect 13955 13481 13964 13515
rect 13912 13472 13964 13481
rect 7380 13447 7432 13456
rect 7380 13413 7389 13447
rect 7389 13413 7423 13447
rect 7423 13413 7432 13447
rect 7380 13404 7432 13413
rect 8484 13404 8536 13456
rect 14740 13404 14792 13456
rect 3148 13268 3200 13320
rect 1584 13200 1636 13252
rect 1676 13243 1728 13252
rect 1676 13209 1685 13243
rect 1685 13209 1719 13243
rect 1719 13209 1728 13243
rect 1676 13200 1728 13209
rect 4896 13200 4948 13252
rect 5724 13268 5776 13320
rect 6920 13336 6972 13388
rect 6000 13268 6052 13320
rect 6276 13268 6328 13320
rect 6828 13268 6880 13320
rect 7656 13336 7708 13388
rect 7748 13268 7800 13320
rect 8208 13311 8260 13320
rect 8208 13277 8217 13311
rect 8217 13277 8251 13311
rect 8251 13277 8260 13311
rect 8208 13268 8260 13277
rect 8760 13311 8812 13320
rect 8760 13277 8769 13311
rect 8769 13277 8803 13311
rect 8803 13277 8812 13311
rect 8760 13268 8812 13277
rect 12532 13268 12584 13320
rect 13176 13311 13228 13320
rect 13176 13277 13185 13311
rect 13185 13277 13219 13311
rect 13219 13277 13228 13311
rect 13176 13268 13228 13277
rect 14464 13336 14516 13388
rect 17040 13472 17092 13524
rect 17776 13515 17828 13524
rect 17776 13481 17785 13515
rect 17785 13481 17819 13515
rect 17819 13481 17828 13515
rect 17776 13472 17828 13481
rect 21732 13515 21784 13524
rect 21732 13481 21741 13515
rect 21741 13481 21775 13515
rect 21775 13481 21784 13515
rect 21732 13472 21784 13481
rect 16304 13379 16356 13388
rect 16304 13345 16313 13379
rect 16313 13345 16347 13379
rect 16347 13345 16356 13379
rect 16304 13336 16356 13345
rect 18512 13379 18564 13388
rect 9036 13243 9088 13252
rect 9036 13209 9045 13243
rect 9045 13209 9079 13243
rect 9079 13209 9088 13243
rect 9036 13200 9088 13209
rect 9404 13243 9456 13252
rect 9404 13209 9413 13243
rect 9413 13209 9447 13243
rect 9447 13209 9456 13243
rect 9404 13200 9456 13209
rect 14280 13268 14332 13320
rect 14096 13200 14148 13252
rect 5448 13132 5500 13184
rect 6276 13175 6328 13184
rect 6276 13141 6285 13175
rect 6285 13141 6319 13175
rect 6319 13141 6328 13175
rect 6276 13132 6328 13141
rect 8392 13132 8444 13184
rect 14924 13200 14976 13252
rect 15384 13311 15436 13320
rect 15384 13277 15393 13311
rect 15393 13277 15427 13311
rect 15427 13277 15436 13311
rect 15384 13268 15436 13277
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 18512 13345 18521 13379
rect 18521 13345 18555 13379
rect 18555 13345 18564 13379
rect 18512 13336 18564 13345
rect 19156 13336 19208 13388
rect 22192 13472 22244 13524
rect 22836 13472 22888 13524
rect 24216 13515 24268 13524
rect 24216 13481 24225 13515
rect 24225 13481 24259 13515
rect 24259 13481 24268 13515
rect 24216 13472 24268 13481
rect 24400 13515 24452 13524
rect 24400 13481 24409 13515
rect 24409 13481 24443 13515
rect 24443 13481 24452 13515
rect 24400 13472 24452 13481
rect 24952 13472 25004 13524
rect 25044 13515 25096 13524
rect 25044 13481 25053 13515
rect 25053 13481 25087 13515
rect 25087 13481 25096 13515
rect 25044 13472 25096 13481
rect 25688 13472 25740 13524
rect 17960 13311 18012 13320
rect 17960 13277 17969 13311
rect 17969 13277 18003 13311
rect 18003 13277 18012 13311
rect 17960 13268 18012 13277
rect 18604 13268 18656 13320
rect 22468 13379 22520 13388
rect 22468 13345 22477 13379
rect 22477 13345 22511 13379
rect 22511 13345 22520 13379
rect 22468 13336 22520 13345
rect 23480 13336 23532 13388
rect 25872 13447 25924 13456
rect 25872 13413 25881 13447
rect 25881 13413 25915 13447
rect 25915 13413 25924 13447
rect 25872 13404 25924 13413
rect 22100 13311 22152 13320
rect 22100 13277 22109 13311
rect 22109 13277 22143 13311
rect 22143 13277 22152 13311
rect 22100 13268 22152 13277
rect 24032 13268 24084 13320
rect 14740 13132 14792 13184
rect 15108 13175 15160 13184
rect 15108 13141 15117 13175
rect 15117 13141 15151 13175
rect 15151 13141 15160 13175
rect 15108 13132 15160 13141
rect 15568 13175 15620 13184
rect 15568 13141 15577 13175
rect 15577 13141 15611 13175
rect 15611 13141 15620 13175
rect 15568 13132 15620 13141
rect 20720 13132 20772 13184
rect 22744 13243 22796 13252
rect 22744 13209 22753 13243
rect 22753 13209 22787 13243
rect 22787 13209 22796 13243
rect 22744 13200 22796 13209
rect 22560 13132 22612 13184
rect 23388 13132 23440 13184
rect 24768 13268 24820 13320
rect 25136 13379 25188 13388
rect 25136 13345 25145 13379
rect 25145 13345 25179 13379
rect 25179 13345 25188 13379
rect 25136 13336 25188 13345
rect 25320 13311 25372 13320
rect 25320 13277 25329 13311
rect 25329 13277 25363 13311
rect 25363 13277 25372 13311
rect 25320 13268 25372 13277
rect 25688 13311 25740 13320
rect 25688 13277 25697 13311
rect 25697 13277 25731 13311
rect 25731 13277 25740 13311
rect 25688 13268 25740 13277
rect 7252 13030 7304 13082
rect 7316 13030 7368 13082
rect 7380 13030 7432 13082
rect 7444 13030 7496 13082
rect 7508 13030 7560 13082
rect 13554 13030 13606 13082
rect 13618 13030 13670 13082
rect 13682 13030 13734 13082
rect 13746 13030 13798 13082
rect 13810 13030 13862 13082
rect 19856 13030 19908 13082
rect 19920 13030 19972 13082
rect 19984 13030 20036 13082
rect 20048 13030 20100 13082
rect 20112 13030 20164 13082
rect 26158 13030 26210 13082
rect 26222 13030 26274 13082
rect 26286 13030 26338 13082
rect 26350 13030 26402 13082
rect 26414 13030 26466 13082
rect 1584 12928 1636 12980
rect 3148 12792 3200 12844
rect 5724 12860 5776 12912
rect 9036 12928 9088 12980
rect 9128 12928 9180 12980
rect 4436 12792 4488 12844
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 5632 12792 5684 12844
rect 4896 12724 4948 12776
rect 5448 12724 5500 12776
rect 6644 12792 6696 12844
rect 7656 12860 7708 12912
rect 6368 12724 6420 12776
rect 6000 12656 6052 12708
rect 5724 12588 5776 12640
rect 5816 12588 5868 12640
rect 6828 12656 6880 12708
rect 7748 12792 7800 12844
rect 8208 12860 8260 12912
rect 9588 12860 9640 12912
rect 8024 12835 8076 12844
rect 8024 12801 8033 12835
rect 8033 12801 8067 12835
rect 8067 12801 8076 12835
rect 8024 12792 8076 12801
rect 12072 12928 12124 12980
rect 12532 12971 12584 12980
rect 12532 12937 12541 12971
rect 12541 12937 12575 12971
rect 12575 12937 12584 12971
rect 12532 12928 12584 12937
rect 13176 12971 13228 12980
rect 13176 12937 13185 12971
rect 13185 12937 13219 12971
rect 13219 12937 13228 12971
rect 13176 12928 13228 12937
rect 10968 12835 11020 12844
rect 10968 12801 10977 12835
rect 10977 12801 11011 12835
rect 11011 12801 11020 12835
rect 10968 12792 11020 12801
rect 6368 12631 6420 12640
rect 6368 12597 6377 12631
rect 6377 12597 6411 12631
rect 6411 12597 6420 12631
rect 6368 12588 6420 12597
rect 7012 12631 7064 12640
rect 7012 12597 7021 12631
rect 7021 12597 7055 12631
rect 7055 12597 7064 12631
rect 7012 12588 7064 12597
rect 8300 12767 8352 12776
rect 8300 12733 8309 12767
rect 8309 12733 8343 12767
rect 8343 12733 8352 12767
rect 8300 12724 8352 12733
rect 9496 12724 9548 12776
rect 11336 12860 11388 12912
rect 12072 12835 12124 12844
rect 12072 12801 12081 12835
rect 12081 12801 12115 12835
rect 12115 12801 12124 12835
rect 12072 12792 12124 12801
rect 12440 12724 12492 12776
rect 12624 12767 12676 12776
rect 12624 12733 12633 12767
rect 12633 12733 12667 12767
rect 12667 12733 12676 12767
rect 12624 12724 12676 12733
rect 13912 12928 13964 12980
rect 14924 12928 14976 12980
rect 15108 12928 15160 12980
rect 15568 12928 15620 12980
rect 13912 12724 13964 12776
rect 9772 12699 9824 12708
rect 9772 12665 9781 12699
rect 9781 12665 9815 12699
rect 9815 12665 9824 12699
rect 9772 12656 9824 12665
rect 8760 12588 8812 12640
rect 10784 12588 10836 12640
rect 11888 12631 11940 12640
rect 11888 12597 11897 12631
rect 11897 12597 11931 12631
rect 11931 12597 11940 12631
rect 11888 12588 11940 12597
rect 13176 12656 13228 12708
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 14556 12792 14608 12844
rect 14924 12835 14976 12844
rect 14924 12801 14933 12835
rect 14933 12801 14967 12835
rect 14967 12801 14976 12835
rect 14924 12792 14976 12801
rect 15660 12860 15712 12912
rect 15752 12860 15804 12912
rect 15476 12835 15528 12844
rect 15476 12801 15485 12835
rect 15485 12801 15519 12835
rect 15519 12801 15528 12835
rect 18512 12860 18564 12912
rect 20260 12860 20312 12912
rect 15476 12792 15528 12801
rect 16396 12835 16448 12844
rect 16396 12801 16405 12835
rect 16405 12801 16439 12835
rect 16439 12801 16448 12835
rect 16396 12792 16448 12801
rect 14464 12656 14516 12708
rect 15936 12699 15988 12708
rect 15936 12665 15945 12699
rect 15945 12665 15979 12699
rect 15979 12665 15988 12699
rect 15936 12656 15988 12665
rect 13820 12588 13872 12640
rect 14280 12588 14332 12640
rect 16304 12588 16356 12640
rect 17224 12767 17276 12776
rect 17224 12733 17233 12767
rect 17233 12733 17267 12767
rect 17267 12733 17276 12767
rect 17224 12724 17276 12733
rect 19616 12724 19668 12776
rect 20536 12792 20588 12844
rect 22744 12928 22796 12980
rect 24676 12928 24728 12980
rect 23756 12903 23808 12912
rect 23756 12869 23765 12903
rect 23765 12869 23799 12903
rect 23799 12869 23808 12903
rect 23756 12860 23808 12869
rect 24032 12860 24084 12912
rect 20352 12724 20404 12776
rect 23480 12835 23532 12844
rect 23480 12801 23489 12835
rect 23489 12801 23523 12835
rect 23523 12801 23532 12835
rect 23480 12792 23532 12801
rect 18420 12588 18472 12640
rect 18788 12631 18840 12640
rect 18788 12597 18797 12631
rect 18797 12597 18831 12631
rect 18831 12597 18840 12631
rect 18788 12588 18840 12597
rect 20996 12588 21048 12640
rect 22100 12588 22152 12640
rect 25228 12724 25280 12776
rect 23296 12588 23348 12640
rect 25136 12588 25188 12640
rect 4101 12486 4153 12538
rect 4165 12486 4217 12538
rect 4229 12486 4281 12538
rect 4293 12486 4345 12538
rect 4357 12486 4409 12538
rect 10403 12486 10455 12538
rect 10467 12486 10519 12538
rect 10531 12486 10583 12538
rect 10595 12486 10647 12538
rect 10659 12486 10711 12538
rect 16705 12486 16757 12538
rect 16769 12486 16821 12538
rect 16833 12486 16885 12538
rect 16897 12486 16949 12538
rect 16961 12486 17013 12538
rect 23007 12486 23059 12538
rect 23071 12486 23123 12538
rect 23135 12486 23187 12538
rect 23199 12486 23251 12538
rect 23263 12486 23315 12538
rect 1676 12384 1728 12436
rect 8300 12384 8352 12436
rect 5724 12316 5776 12368
rect 7840 12316 7892 12368
rect 12440 12384 12492 12436
rect 12716 12384 12768 12436
rect 3700 12248 3752 12300
rect 4712 12291 4764 12300
rect 4712 12257 4721 12291
rect 4721 12257 4755 12291
rect 4755 12257 4764 12291
rect 4712 12248 4764 12257
rect 6092 12248 6144 12300
rect 940 12180 992 12232
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 5908 12180 5960 12232
rect 6736 12248 6788 12300
rect 2044 12155 2096 12164
rect 2044 12121 2053 12155
rect 2053 12121 2087 12155
rect 2087 12121 2096 12155
rect 2044 12112 2096 12121
rect 2780 12112 2832 12164
rect 1400 12044 1452 12096
rect 3976 12112 4028 12164
rect 6368 12155 6420 12164
rect 6368 12121 6377 12155
rect 6377 12121 6411 12155
rect 6411 12121 6420 12155
rect 6368 12112 6420 12121
rect 6644 12180 6696 12232
rect 6920 12223 6972 12232
rect 6920 12189 6929 12223
rect 6929 12189 6963 12223
rect 6963 12189 6972 12223
rect 6920 12180 6972 12189
rect 9772 12248 9824 12300
rect 10232 12248 10284 12300
rect 11152 12248 11204 12300
rect 13176 12291 13228 12300
rect 13176 12257 13185 12291
rect 13185 12257 13219 12291
rect 13219 12257 13228 12291
rect 13176 12248 13228 12257
rect 7104 12180 7156 12232
rect 8392 12180 8444 12232
rect 9404 12180 9456 12232
rect 10140 12180 10192 12232
rect 14096 12316 14148 12368
rect 13820 12248 13872 12300
rect 3608 12044 3660 12096
rect 6920 12044 6972 12096
rect 9128 12087 9180 12096
rect 9128 12053 9137 12087
rect 9137 12053 9171 12087
rect 9171 12053 9180 12087
rect 9128 12044 9180 12053
rect 10784 12155 10836 12164
rect 10784 12121 10793 12155
rect 10793 12121 10827 12155
rect 10827 12121 10836 12155
rect 10784 12112 10836 12121
rect 12992 12112 13044 12164
rect 13912 12223 13964 12232
rect 13912 12189 13921 12223
rect 13921 12189 13955 12223
rect 13955 12189 13964 12223
rect 13912 12180 13964 12189
rect 14464 12248 14516 12300
rect 17224 12384 17276 12436
rect 15292 12248 15344 12300
rect 15660 12248 15712 12300
rect 20904 12384 20956 12436
rect 22100 12384 22152 12436
rect 17684 12248 17736 12300
rect 18052 12291 18104 12300
rect 18052 12257 18061 12291
rect 18061 12257 18095 12291
rect 18095 12257 18104 12291
rect 18052 12248 18104 12257
rect 14556 12112 14608 12164
rect 14832 12223 14884 12232
rect 14832 12189 14841 12223
rect 14841 12189 14875 12223
rect 14875 12189 14884 12223
rect 14832 12180 14884 12189
rect 14924 12223 14976 12232
rect 14924 12189 14933 12223
rect 14933 12189 14967 12223
rect 14967 12189 14976 12223
rect 14924 12180 14976 12189
rect 15016 12112 15068 12164
rect 15384 12112 15436 12164
rect 12348 12044 12400 12096
rect 14924 12044 14976 12096
rect 15568 12087 15620 12096
rect 15568 12053 15577 12087
rect 15577 12053 15611 12087
rect 15611 12053 15620 12087
rect 15568 12044 15620 12053
rect 15752 12087 15804 12096
rect 15752 12053 15761 12087
rect 15761 12053 15795 12087
rect 15795 12053 15804 12087
rect 15752 12044 15804 12053
rect 18788 12180 18840 12232
rect 20168 12223 20220 12232
rect 20168 12189 20177 12223
rect 20177 12189 20211 12223
rect 20211 12189 20220 12223
rect 20168 12180 20220 12189
rect 20260 12180 20312 12232
rect 22468 12248 22520 12300
rect 17960 12044 18012 12096
rect 18972 12044 19024 12096
rect 20352 12112 20404 12164
rect 20720 12155 20772 12164
rect 20720 12121 20729 12155
rect 20729 12121 20763 12155
rect 20763 12121 20772 12155
rect 20720 12112 20772 12121
rect 7252 11942 7304 11994
rect 7316 11942 7368 11994
rect 7380 11942 7432 11994
rect 7444 11942 7496 11994
rect 7508 11942 7560 11994
rect 13554 11942 13606 11994
rect 13618 11942 13670 11994
rect 13682 11942 13734 11994
rect 13746 11942 13798 11994
rect 13810 11942 13862 11994
rect 19856 11942 19908 11994
rect 19920 11942 19972 11994
rect 19984 11942 20036 11994
rect 20048 11942 20100 11994
rect 20112 11942 20164 11994
rect 26158 11942 26210 11994
rect 26222 11942 26274 11994
rect 26286 11942 26338 11994
rect 26350 11942 26402 11994
rect 26414 11942 26466 11994
rect 2044 11840 2096 11892
rect 2780 11704 2832 11756
rect 3608 11840 3660 11892
rect 9772 11840 9824 11892
rect 10324 11840 10376 11892
rect 14004 11840 14056 11892
rect 14188 11840 14240 11892
rect 15016 11840 15068 11892
rect 4896 11772 4948 11824
rect 5540 11772 5592 11824
rect 10784 11772 10836 11824
rect 11152 11815 11204 11824
rect 11152 11781 11161 11815
rect 11161 11781 11195 11815
rect 11195 11781 11204 11815
rect 11152 11772 11204 11781
rect 11888 11815 11940 11824
rect 11888 11781 11897 11815
rect 11897 11781 11931 11815
rect 11931 11781 11940 11815
rect 11888 11772 11940 11781
rect 12348 11772 12400 11824
rect 13176 11772 13228 11824
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 5908 11747 5960 11756
rect 5908 11713 5917 11747
rect 5917 11713 5951 11747
rect 5951 11713 5960 11747
rect 5908 11704 5960 11713
rect 6644 11704 6696 11756
rect 7012 11704 7064 11756
rect 9864 11747 9916 11756
rect 9864 11713 9873 11747
rect 9873 11713 9907 11747
rect 9907 11713 9916 11747
rect 9864 11704 9916 11713
rect 3884 11500 3936 11552
rect 7196 11636 7248 11688
rect 10324 11745 10376 11756
rect 10324 11711 10333 11745
rect 10333 11711 10367 11745
rect 10367 11711 10376 11745
rect 10324 11704 10376 11711
rect 11612 11747 11664 11756
rect 11612 11713 11621 11747
rect 11621 11713 11655 11747
rect 11655 11713 11664 11747
rect 11612 11704 11664 11713
rect 13636 11747 13688 11756
rect 13636 11713 13645 11747
rect 13645 11713 13679 11747
rect 13679 11713 13688 11747
rect 13636 11704 13688 11713
rect 13820 11772 13872 11824
rect 14832 11772 14884 11824
rect 14096 11704 14148 11756
rect 14648 11704 14700 11756
rect 15016 11747 15068 11756
rect 15016 11713 15025 11747
rect 15025 11713 15059 11747
rect 15059 11713 15068 11747
rect 15016 11704 15068 11713
rect 5540 11500 5592 11552
rect 9404 11568 9456 11620
rect 6736 11543 6788 11552
rect 6736 11509 6745 11543
rect 6745 11509 6779 11543
rect 6779 11509 6788 11543
rect 6736 11500 6788 11509
rect 9588 11500 9640 11552
rect 14556 11636 14608 11688
rect 15384 11840 15436 11892
rect 16304 11840 16356 11892
rect 15384 11747 15436 11756
rect 15384 11713 15393 11747
rect 15393 11713 15427 11747
rect 15427 11713 15436 11747
rect 15384 11704 15436 11713
rect 15476 11704 15528 11756
rect 18236 11772 18288 11824
rect 17224 11704 17276 11756
rect 18420 11747 18472 11756
rect 18420 11713 18429 11747
rect 18429 11713 18463 11747
rect 18463 11713 18472 11747
rect 18420 11704 18472 11713
rect 24768 11840 24820 11892
rect 25688 11840 25740 11892
rect 22284 11772 22336 11824
rect 22744 11772 22796 11824
rect 24032 11772 24084 11824
rect 20536 11704 20588 11756
rect 22100 11747 22152 11756
rect 22100 11713 22109 11747
rect 22109 11713 22143 11747
rect 22143 11713 22152 11747
rect 22100 11704 22152 11713
rect 22468 11704 22520 11756
rect 16396 11636 16448 11688
rect 18696 11679 18748 11688
rect 18696 11645 18705 11679
rect 18705 11645 18739 11679
rect 18739 11645 18748 11679
rect 18696 11636 18748 11645
rect 20812 11679 20864 11688
rect 20812 11645 20821 11679
rect 20821 11645 20855 11679
rect 20855 11645 20864 11679
rect 20812 11636 20864 11645
rect 11244 11568 11296 11620
rect 23480 11679 23532 11688
rect 23480 11645 23489 11679
rect 23489 11645 23523 11679
rect 23523 11645 23532 11679
rect 23480 11636 23532 11645
rect 13820 11500 13872 11552
rect 15844 11543 15896 11552
rect 15844 11509 15853 11543
rect 15853 11509 15887 11543
rect 15887 11509 15896 11543
rect 15844 11500 15896 11509
rect 20352 11500 20404 11552
rect 20904 11500 20956 11552
rect 22008 11543 22060 11552
rect 22008 11509 22017 11543
rect 22017 11509 22051 11543
rect 22051 11509 22060 11543
rect 22008 11500 22060 11509
rect 22560 11500 22612 11552
rect 22836 11500 22888 11552
rect 4101 11398 4153 11450
rect 4165 11398 4217 11450
rect 4229 11398 4281 11450
rect 4293 11398 4345 11450
rect 4357 11398 4409 11450
rect 10403 11398 10455 11450
rect 10467 11398 10519 11450
rect 10531 11398 10583 11450
rect 10595 11398 10647 11450
rect 10659 11398 10711 11450
rect 16705 11398 16757 11450
rect 16769 11398 16821 11450
rect 16833 11398 16885 11450
rect 16897 11398 16949 11450
rect 16961 11398 17013 11450
rect 23007 11398 23059 11450
rect 23071 11398 23123 11450
rect 23135 11398 23187 11450
rect 23199 11398 23251 11450
rect 23263 11398 23315 11450
rect 3700 11296 3752 11348
rect 5540 11296 5592 11348
rect 5908 11296 5960 11348
rect 6736 11296 6788 11348
rect 6920 11296 6972 11348
rect 9128 11296 9180 11348
rect 10784 11296 10836 11348
rect 1400 11024 1452 11076
rect 3792 11228 3844 11280
rect 4896 11228 4948 11280
rect 7104 11228 7156 11280
rect 4712 11160 4764 11212
rect 6092 11203 6144 11212
rect 6092 11169 6101 11203
rect 6101 11169 6135 11203
rect 6135 11169 6144 11203
rect 6092 11160 6144 11169
rect 3148 11092 3200 11144
rect 5816 11135 5868 11144
rect 5816 11101 5825 11135
rect 5825 11101 5859 11135
rect 5859 11101 5868 11135
rect 5816 11092 5868 11101
rect 5908 11135 5960 11144
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 5908 11092 5960 11101
rect 6644 11092 6696 11144
rect 7564 11135 7616 11144
rect 7564 11101 7573 11135
rect 7573 11101 7607 11135
rect 7607 11101 7616 11135
rect 7564 11092 7616 11101
rect 3608 10999 3660 11008
rect 3608 10965 3617 10999
rect 3617 10965 3651 10999
rect 3651 10965 3660 10999
rect 3608 10956 3660 10965
rect 6000 10956 6052 11008
rect 6368 10956 6420 11008
rect 7932 11160 7984 11212
rect 8576 11160 8628 11212
rect 8944 11160 8996 11212
rect 10416 11160 10468 11212
rect 9312 11067 9364 11076
rect 9312 11033 9321 11067
rect 9321 11033 9355 11067
rect 9355 11033 9364 11067
rect 9312 11024 9364 11033
rect 8852 10956 8904 11008
rect 9128 10956 9180 11008
rect 9588 11135 9640 11144
rect 9588 11101 9597 11135
rect 9597 11101 9631 11135
rect 9631 11101 9640 11135
rect 9588 11092 9640 11101
rect 11244 11160 11296 11212
rect 11336 11203 11388 11212
rect 11336 11169 11345 11203
rect 11345 11169 11379 11203
rect 11379 11169 11388 11203
rect 11336 11160 11388 11169
rect 11612 11203 11664 11212
rect 11612 11169 11621 11203
rect 11621 11169 11655 11203
rect 11655 11169 11664 11203
rect 11612 11160 11664 11169
rect 18696 11296 18748 11348
rect 23480 11296 23532 11348
rect 25320 11339 25372 11348
rect 25320 11305 25329 11339
rect 25329 11305 25363 11339
rect 25363 11305 25372 11339
rect 25320 11296 25372 11305
rect 14648 11160 14700 11212
rect 17408 11160 17460 11212
rect 18420 11160 18472 11212
rect 21088 11203 21140 11212
rect 21088 11169 21097 11203
rect 21097 11169 21131 11203
rect 21131 11169 21140 11203
rect 21088 11160 21140 11169
rect 21548 11160 21600 11212
rect 22008 11160 22060 11212
rect 22192 11160 22244 11212
rect 22468 11160 22520 11212
rect 11060 11135 11112 11144
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 11060 11092 11112 11101
rect 14464 11135 14516 11144
rect 10048 11067 10100 11076
rect 10048 11033 10057 11067
rect 10057 11033 10091 11067
rect 10091 11033 10100 11067
rect 10048 11024 10100 11033
rect 9680 10956 9732 11008
rect 10784 10956 10836 11008
rect 12348 11024 12400 11076
rect 14464 11101 14473 11135
rect 14473 11101 14507 11135
rect 14507 11101 14516 11135
rect 14464 11092 14516 11101
rect 15752 11092 15804 11144
rect 17500 11092 17552 11144
rect 14188 11024 14240 11076
rect 18972 11135 19024 11144
rect 18972 11101 18981 11135
rect 18981 11101 19015 11135
rect 19015 11101 19024 11135
rect 18972 11092 19024 11101
rect 20812 11092 20864 11144
rect 21456 11092 21508 11144
rect 23388 11092 23440 11144
rect 17040 10999 17092 11008
rect 17040 10965 17049 10999
rect 17049 10965 17083 10999
rect 17083 10965 17092 10999
rect 17040 10956 17092 10965
rect 17316 10999 17368 11008
rect 17316 10965 17325 10999
rect 17325 10965 17359 10999
rect 17359 10965 17368 10999
rect 17316 10956 17368 10965
rect 19248 11024 19300 11076
rect 19524 11067 19576 11076
rect 19524 11033 19533 11067
rect 19533 11033 19567 11067
rect 19567 11033 19576 11067
rect 19524 11024 19576 11033
rect 22284 11024 22336 11076
rect 22652 11024 22704 11076
rect 25688 11135 25740 11144
rect 25688 11101 25697 11135
rect 25697 11101 25731 11135
rect 25731 11101 25740 11135
rect 25688 11092 25740 11101
rect 19708 10956 19760 11008
rect 20904 10956 20956 11008
rect 21272 10956 21324 11008
rect 24400 10956 24452 11008
rect 7252 10854 7304 10906
rect 7316 10854 7368 10906
rect 7380 10854 7432 10906
rect 7444 10854 7496 10906
rect 7508 10854 7560 10906
rect 13554 10854 13606 10906
rect 13618 10854 13670 10906
rect 13682 10854 13734 10906
rect 13746 10854 13798 10906
rect 13810 10854 13862 10906
rect 19856 10854 19908 10906
rect 19920 10854 19972 10906
rect 19984 10854 20036 10906
rect 20048 10854 20100 10906
rect 20112 10854 20164 10906
rect 26158 10854 26210 10906
rect 26222 10854 26274 10906
rect 26286 10854 26338 10906
rect 26350 10854 26402 10906
rect 26414 10854 26466 10906
rect 3148 10752 3200 10804
rect 5908 10752 5960 10804
rect 6736 10795 6788 10804
rect 6736 10761 6745 10795
rect 6745 10761 6779 10795
rect 6779 10761 6788 10795
rect 7104 10795 7156 10804
rect 6736 10752 6788 10761
rect 2780 10684 2832 10736
rect 3792 10616 3844 10668
rect 4712 10616 4764 10668
rect 6000 10684 6052 10736
rect 6092 10684 6144 10736
rect 7104 10761 7131 10795
rect 7131 10761 7156 10795
rect 7104 10752 7156 10761
rect 7564 10752 7616 10804
rect 8668 10752 8720 10804
rect 6460 10616 6512 10668
rect 3608 10591 3660 10600
rect 3608 10557 3617 10591
rect 3617 10557 3651 10591
rect 3651 10557 3660 10591
rect 3608 10548 3660 10557
rect 5632 10591 5684 10600
rect 5632 10557 5641 10591
rect 5641 10557 5675 10591
rect 5675 10557 5684 10591
rect 5632 10548 5684 10557
rect 6184 10548 6236 10600
rect 6368 10548 6420 10600
rect 6920 10616 6972 10668
rect 7196 10616 7248 10668
rect 8944 10795 8996 10804
rect 8944 10761 8953 10795
rect 8953 10761 8987 10795
rect 8987 10761 8996 10795
rect 8944 10752 8996 10761
rect 9864 10752 9916 10804
rect 10140 10684 10192 10736
rect 10968 10752 11020 10804
rect 7564 10659 7616 10668
rect 7564 10625 7573 10659
rect 7573 10625 7607 10659
rect 7607 10625 7616 10659
rect 7564 10616 7616 10625
rect 8484 10616 8536 10668
rect 8668 10616 8720 10668
rect 8852 10659 8904 10668
rect 8852 10625 8861 10659
rect 8861 10625 8895 10659
rect 8895 10625 8904 10659
rect 8852 10616 8904 10625
rect 9036 10616 9088 10668
rect 9312 10616 9364 10668
rect 9956 10659 10008 10668
rect 9956 10625 9965 10659
rect 9965 10625 9999 10659
rect 9999 10625 10008 10659
rect 9956 10616 10008 10625
rect 10232 10616 10284 10668
rect 10416 10659 10468 10668
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 10416 10616 10468 10625
rect 10692 10659 10744 10668
rect 10692 10625 10701 10659
rect 10701 10625 10735 10659
rect 10735 10625 10744 10659
rect 10692 10616 10744 10625
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 6644 10480 6696 10532
rect 3056 10412 3108 10464
rect 3700 10455 3752 10464
rect 3700 10421 3709 10455
rect 3709 10421 3743 10455
rect 3743 10421 3752 10455
rect 3700 10412 3752 10421
rect 5448 10455 5500 10464
rect 5448 10421 5457 10455
rect 5457 10421 5491 10455
rect 5491 10421 5500 10455
rect 5448 10412 5500 10421
rect 7012 10412 7064 10464
rect 7196 10412 7248 10464
rect 8760 10548 8812 10600
rect 9128 10523 9180 10532
rect 9128 10489 9137 10523
rect 9137 10489 9171 10523
rect 9171 10489 9180 10523
rect 9128 10480 9180 10489
rect 7748 10412 7800 10464
rect 9680 10412 9732 10464
rect 9956 10412 10008 10464
rect 10784 10412 10836 10464
rect 15660 10412 15712 10464
rect 16028 10412 16080 10464
rect 16120 10455 16172 10464
rect 16120 10421 16129 10455
rect 16129 10421 16163 10455
rect 16163 10421 16172 10455
rect 16120 10412 16172 10421
rect 17316 10752 17368 10804
rect 17500 10795 17552 10804
rect 17500 10761 17509 10795
rect 17509 10761 17543 10795
rect 17543 10761 17552 10795
rect 17500 10752 17552 10761
rect 18880 10752 18932 10804
rect 19248 10752 19300 10804
rect 19524 10752 19576 10804
rect 20628 10752 20680 10804
rect 22468 10752 22520 10804
rect 19156 10684 19208 10736
rect 17776 10616 17828 10668
rect 17684 10480 17736 10532
rect 19432 10616 19484 10668
rect 19524 10659 19576 10668
rect 19524 10625 19533 10659
rect 19533 10625 19567 10659
rect 19567 10625 19576 10659
rect 19524 10616 19576 10625
rect 20996 10684 21048 10736
rect 20352 10659 20404 10668
rect 20352 10625 20361 10659
rect 20361 10625 20395 10659
rect 20395 10625 20404 10659
rect 20352 10616 20404 10625
rect 21548 10616 21600 10668
rect 23848 10684 23900 10736
rect 24124 10684 24176 10736
rect 20812 10548 20864 10600
rect 22560 10548 22612 10600
rect 24216 10591 24268 10600
rect 20904 10480 20956 10532
rect 21824 10455 21876 10464
rect 21824 10421 21833 10455
rect 21833 10421 21867 10455
rect 21867 10421 21876 10455
rect 21824 10412 21876 10421
rect 24216 10557 24225 10591
rect 24225 10557 24259 10591
rect 24259 10557 24268 10591
rect 24216 10548 24268 10557
rect 24400 10548 24452 10600
rect 24952 10548 25004 10600
rect 25780 10591 25832 10600
rect 25780 10557 25789 10591
rect 25789 10557 25823 10591
rect 25823 10557 25832 10591
rect 25780 10548 25832 10557
rect 25504 10412 25556 10464
rect 4101 10310 4153 10362
rect 4165 10310 4217 10362
rect 4229 10310 4281 10362
rect 4293 10310 4345 10362
rect 4357 10310 4409 10362
rect 10403 10310 10455 10362
rect 10467 10310 10519 10362
rect 10531 10310 10583 10362
rect 10595 10310 10647 10362
rect 10659 10310 10711 10362
rect 16705 10310 16757 10362
rect 16769 10310 16821 10362
rect 16833 10310 16885 10362
rect 16897 10310 16949 10362
rect 16961 10310 17013 10362
rect 23007 10310 23059 10362
rect 23071 10310 23123 10362
rect 23135 10310 23187 10362
rect 23199 10310 23251 10362
rect 23263 10310 23315 10362
rect 5448 10208 5500 10260
rect 5632 10208 5684 10260
rect 6092 10251 6144 10260
rect 6092 10217 6101 10251
rect 6101 10217 6135 10251
rect 6135 10217 6144 10251
rect 6092 10208 6144 10217
rect 6184 10208 6236 10260
rect 7564 10208 7616 10260
rect 8484 10208 8536 10260
rect 9036 10251 9088 10260
rect 9036 10217 9045 10251
rect 9045 10217 9079 10251
rect 9079 10217 9088 10251
rect 9036 10208 9088 10217
rect 9864 10251 9916 10260
rect 9864 10217 9873 10251
rect 9873 10217 9907 10251
rect 9907 10217 9916 10251
rect 9864 10208 9916 10217
rect 10232 10208 10284 10260
rect 16120 10208 16172 10260
rect 19432 10208 19484 10260
rect 21824 10208 21876 10260
rect 22100 10208 22152 10260
rect 23388 10208 23440 10260
rect 24216 10208 24268 10260
rect 25780 10208 25832 10260
rect 2872 10115 2924 10124
rect 2872 10081 2881 10115
rect 2881 10081 2915 10115
rect 2915 10081 2924 10115
rect 2872 10072 2924 10081
rect 3056 10004 3108 10056
rect 3240 9936 3292 9988
rect 3976 10047 4028 10056
rect 3976 10013 3985 10047
rect 3985 10013 4019 10047
rect 4019 10013 4028 10047
rect 3976 10004 4028 10013
rect 4068 10004 4120 10056
rect 5540 10115 5592 10124
rect 5540 10081 5549 10115
rect 5549 10081 5583 10115
rect 5583 10081 5592 10115
rect 5540 10072 5592 10081
rect 6736 10115 6788 10124
rect 6736 10081 6745 10115
rect 6745 10081 6779 10115
rect 6779 10081 6788 10115
rect 6736 10072 6788 10081
rect 4620 9936 4672 9988
rect 5632 10047 5684 10056
rect 5632 10013 5641 10047
rect 5641 10013 5675 10047
rect 5675 10013 5684 10047
rect 5632 10004 5684 10013
rect 6368 10047 6420 10056
rect 6368 10013 6377 10047
rect 6377 10013 6411 10047
rect 6411 10013 6420 10047
rect 6368 10004 6420 10013
rect 6828 10004 6880 10056
rect 7564 10004 7616 10056
rect 7748 10004 7800 10056
rect 7932 10047 7984 10056
rect 7932 10013 7941 10047
rect 7941 10013 7975 10047
rect 7975 10013 7984 10047
rect 7932 10004 7984 10013
rect 7012 9936 7064 9988
rect 8668 10004 8720 10056
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 9680 10115 9732 10124
rect 9680 10081 9689 10115
rect 9689 10081 9723 10115
rect 9723 10081 9732 10115
rect 9680 10072 9732 10081
rect 9956 10004 10008 10056
rect 2412 9911 2464 9920
rect 2412 9877 2421 9911
rect 2421 9877 2455 9911
rect 2455 9877 2464 9911
rect 2412 9868 2464 9877
rect 5540 9868 5592 9920
rect 8576 9911 8628 9920
rect 8576 9877 8585 9911
rect 8585 9877 8619 9911
rect 8619 9877 8628 9911
rect 8576 9868 8628 9877
rect 9864 9936 9916 9988
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 10600 9936 10652 9988
rect 14372 10072 14424 10124
rect 15660 10115 15712 10124
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 18420 10072 18472 10124
rect 20260 10072 20312 10124
rect 14924 10047 14976 10056
rect 14924 10013 14933 10047
rect 14933 10013 14967 10047
rect 14967 10013 14976 10047
rect 14924 10004 14976 10013
rect 17224 10004 17276 10056
rect 23848 10072 23900 10124
rect 21824 10047 21876 10056
rect 21824 10013 21833 10047
rect 21833 10013 21867 10047
rect 21867 10013 21876 10047
rect 21824 10004 21876 10013
rect 22376 10004 22428 10056
rect 24216 10047 24268 10056
rect 24216 10013 24225 10047
rect 24225 10013 24259 10047
rect 24259 10013 24268 10047
rect 25136 10047 25188 10056
rect 24216 10004 24268 10013
rect 25136 10013 25145 10047
rect 25145 10013 25179 10047
rect 25179 10013 25188 10047
rect 25136 10004 25188 10013
rect 25872 10047 25924 10056
rect 25872 10013 25881 10047
rect 25881 10013 25915 10047
rect 25915 10013 25924 10047
rect 25872 10004 25924 10013
rect 10692 9868 10744 9920
rect 14004 9868 14056 9920
rect 14648 9868 14700 9920
rect 15292 9868 15344 9920
rect 21456 9936 21508 9988
rect 23848 9936 23900 9988
rect 23940 9979 23992 9988
rect 23940 9945 23949 9979
rect 23949 9945 23983 9979
rect 23983 9945 23992 9979
rect 23940 9936 23992 9945
rect 17224 9868 17276 9920
rect 17316 9868 17368 9920
rect 21180 9868 21232 9920
rect 22652 9868 22704 9920
rect 25504 9936 25556 9988
rect 7252 9766 7304 9818
rect 7316 9766 7368 9818
rect 7380 9766 7432 9818
rect 7444 9766 7496 9818
rect 7508 9766 7560 9818
rect 13554 9766 13606 9818
rect 13618 9766 13670 9818
rect 13682 9766 13734 9818
rect 13746 9766 13798 9818
rect 13810 9766 13862 9818
rect 19856 9766 19908 9818
rect 19920 9766 19972 9818
rect 19984 9766 20036 9818
rect 20048 9766 20100 9818
rect 20112 9766 20164 9818
rect 26158 9766 26210 9818
rect 26222 9766 26274 9818
rect 26286 9766 26338 9818
rect 26350 9766 26402 9818
rect 26414 9766 26466 9818
rect 3976 9664 4028 9716
rect 2228 9596 2280 9648
rect 2596 9596 2648 9648
rect 2872 9528 2924 9580
rect 3148 9460 3200 9512
rect 1768 9392 1820 9444
rect 3884 9639 3936 9648
rect 3884 9605 3893 9639
rect 3893 9605 3927 9639
rect 3927 9605 3936 9639
rect 3884 9596 3936 9605
rect 3976 9528 4028 9580
rect 4160 9571 4212 9580
rect 4160 9537 4169 9571
rect 4169 9537 4203 9571
rect 4203 9537 4212 9571
rect 4344 9605 4353 9614
rect 4353 9605 4387 9614
rect 4387 9605 4396 9614
rect 4344 9562 4396 9605
rect 4712 9664 4764 9716
rect 6736 9664 6788 9716
rect 6920 9664 6972 9716
rect 7656 9664 7708 9716
rect 8760 9664 8812 9716
rect 8852 9664 8904 9716
rect 9588 9664 9640 9716
rect 9680 9664 9732 9716
rect 10692 9707 10744 9716
rect 10692 9673 10701 9707
rect 10701 9673 10735 9707
rect 10735 9673 10744 9707
rect 10692 9664 10744 9673
rect 10784 9664 10836 9716
rect 14372 9664 14424 9716
rect 14924 9664 14976 9716
rect 17132 9664 17184 9716
rect 17224 9664 17276 9716
rect 22836 9664 22888 9716
rect 24400 9664 24452 9716
rect 25872 9707 25924 9716
rect 25872 9673 25881 9707
rect 25881 9673 25915 9707
rect 25915 9673 25924 9707
rect 25872 9664 25924 9673
rect 4160 9528 4212 9537
rect 3332 9460 3384 9512
rect 2136 9367 2188 9376
rect 2136 9333 2145 9367
rect 2145 9333 2179 9367
rect 2179 9333 2188 9367
rect 2136 9324 2188 9333
rect 2964 9324 3016 9376
rect 3240 9367 3292 9376
rect 3240 9333 3249 9367
rect 3249 9333 3283 9367
rect 3283 9333 3292 9367
rect 3240 9324 3292 9333
rect 3700 9367 3752 9376
rect 3700 9333 3709 9367
rect 3709 9333 3743 9367
rect 3743 9333 3752 9367
rect 3700 9324 3752 9333
rect 3976 9324 4028 9376
rect 4528 9571 4580 9580
rect 4528 9537 4537 9571
rect 4537 9537 4571 9571
rect 4571 9537 4580 9571
rect 4528 9528 4580 9537
rect 4804 9528 4856 9580
rect 6828 9528 6880 9580
rect 8484 9571 8536 9580
rect 8484 9537 8493 9571
rect 8493 9537 8527 9571
rect 8527 9537 8536 9571
rect 8484 9528 8536 9537
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 9864 9528 9916 9580
rect 10048 9596 10100 9648
rect 10968 9596 11020 9648
rect 10140 9528 10192 9580
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 10416 9528 10468 9580
rect 5816 9392 5868 9444
rect 10600 9460 10652 9512
rect 10876 9392 10928 9444
rect 11152 9571 11204 9580
rect 11152 9537 11183 9571
rect 11183 9537 11204 9571
rect 11152 9528 11204 9537
rect 17040 9596 17092 9648
rect 19708 9596 19760 9648
rect 23848 9596 23900 9648
rect 25320 9596 25372 9648
rect 11060 9392 11112 9444
rect 4528 9324 4580 9376
rect 4620 9324 4672 9376
rect 5632 9324 5684 9376
rect 10416 9324 10468 9376
rect 14096 9528 14148 9580
rect 15108 9528 15160 9580
rect 15200 9571 15252 9580
rect 15200 9537 15209 9571
rect 15209 9537 15243 9571
rect 15243 9537 15252 9571
rect 15200 9528 15252 9537
rect 16028 9528 16080 9580
rect 12992 9503 13044 9512
rect 12992 9469 13001 9503
rect 13001 9469 13035 9503
rect 13035 9469 13044 9503
rect 12992 9460 13044 9469
rect 14648 9460 14700 9512
rect 17592 9460 17644 9512
rect 22652 9528 22704 9580
rect 24952 9528 25004 9580
rect 25136 9528 25188 9580
rect 19616 9460 19668 9512
rect 21088 9460 21140 9512
rect 11336 9324 11388 9376
rect 13728 9324 13780 9376
rect 16396 9324 16448 9376
rect 17684 9324 17736 9376
rect 18972 9392 19024 9444
rect 21180 9392 21232 9444
rect 19248 9367 19300 9376
rect 19248 9333 19257 9367
rect 19257 9333 19291 9367
rect 19291 9333 19300 9367
rect 19248 9324 19300 9333
rect 19616 9324 19668 9376
rect 21640 9324 21692 9376
rect 25688 9367 25740 9376
rect 25688 9333 25697 9367
rect 25697 9333 25731 9367
rect 25731 9333 25740 9367
rect 25688 9324 25740 9333
rect 4101 9222 4153 9274
rect 4165 9222 4217 9274
rect 4229 9222 4281 9274
rect 4293 9222 4345 9274
rect 4357 9222 4409 9274
rect 10403 9222 10455 9274
rect 10467 9222 10519 9274
rect 10531 9222 10583 9274
rect 10595 9222 10647 9274
rect 10659 9222 10711 9274
rect 16705 9222 16757 9274
rect 16769 9222 16821 9274
rect 16833 9222 16885 9274
rect 16897 9222 16949 9274
rect 16961 9222 17013 9274
rect 23007 9222 23059 9274
rect 23071 9222 23123 9274
rect 23135 9222 23187 9274
rect 23199 9222 23251 9274
rect 23263 9222 23315 9274
rect 2688 9120 2740 9172
rect 3240 9120 3292 9172
rect 3884 9120 3936 9172
rect 4436 9120 4488 9172
rect 6552 9120 6604 9172
rect 2412 8984 2464 9036
rect 2872 8984 2924 9036
rect 4252 9052 4304 9104
rect 5264 9052 5316 9104
rect 8484 9120 8536 9172
rect 9404 9120 9456 9172
rect 10876 9120 10928 9172
rect 11336 9120 11388 9172
rect 12992 9120 13044 9172
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 2780 8916 2832 8968
rect 3884 8916 3936 8968
rect 4896 8984 4948 9036
rect 7748 9052 7800 9104
rect 8668 9052 8720 9104
rect 8760 9052 8812 9104
rect 15108 9120 15160 9172
rect 17960 9120 18012 9172
rect 19248 9120 19300 9172
rect 14004 9052 14056 9104
rect 14648 9052 14700 9104
rect 16396 9052 16448 9104
rect 4160 8916 4212 8968
rect 4620 8916 4672 8968
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 4068 8848 4120 8900
rect 5264 8959 5316 8968
rect 5264 8925 5273 8959
rect 5273 8925 5307 8959
rect 5307 8925 5316 8959
rect 5264 8916 5316 8925
rect 7104 8891 7156 8900
rect 3792 8780 3844 8832
rect 7104 8857 7113 8891
rect 7113 8857 7147 8891
rect 7147 8857 7156 8891
rect 7104 8848 7156 8857
rect 6736 8780 6788 8832
rect 8392 8916 8444 8968
rect 9956 8916 10008 8968
rect 12072 8984 12124 9036
rect 10324 8848 10376 8900
rect 10876 8848 10928 8900
rect 11612 8823 11664 8832
rect 11612 8789 11621 8823
rect 11621 8789 11655 8823
rect 11655 8789 11664 8823
rect 11612 8780 11664 8789
rect 11796 8780 11848 8832
rect 12348 8780 12400 8832
rect 15200 8984 15252 9036
rect 15292 8984 15344 9036
rect 16028 8984 16080 9036
rect 17684 8984 17736 9036
rect 18420 9027 18472 9036
rect 18420 8993 18429 9027
rect 18429 8993 18463 9027
rect 18463 8993 18472 9027
rect 18420 8984 18472 8993
rect 18512 8984 18564 9036
rect 17040 8916 17092 8968
rect 17132 8848 17184 8900
rect 17592 8848 17644 8900
rect 19248 8916 19300 8968
rect 23848 8916 23900 8968
rect 24216 8916 24268 8968
rect 20720 8848 20772 8900
rect 21456 8848 21508 8900
rect 15016 8780 15068 8832
rect 16580 8780 16632 8832
rect 17224 8823 17276 8832
rect 17224 8789 17233 8823
rect 17233 8789 17267 8823
rect 17267 8789 17276 8823
rect 17224 8780 17276 8789
rect 18604 8780 18656 8832
rect 18696 8823 18748 8832
rect 18696 8789 18705 8823
rect 18705 8789 18739 8823
rect 18739 8789 18748 8823
rect 18696 8780 18748 8789
rect 19340 8780 19392 8832
rect 21916 8823 21968 8832
rect 21916 8789 21925 8823
rect 21925 8789 21959 8823
rect 21959 8789 21968 8823
rect 21916 8780 21968 8789
rect 23572 8780 23624 8832
rect 25320 8848 25372 8900
rect 24952 8780 25004 8832
rect 7252 8678 7304 8730
rect 7316 8678 7368 8730
rect 7380 8678 7432 8730
rect 7444 8678 7496 8730
rect 7508 8678 7560 8730
rect 13554 8678 13606 8730
rect 13618 8678 13670 8730
rect 13682 8678 13734 8730
rect 13746 8678 13798 8730
rect 13810 8678 13862 8730
rect 19856 8678 19908 8730
rect 19920 8678 19972 8730
rect 19984 8678 20036 8730
rect 20048 8678 20100 8730
rect 20112 8678 20164 8730
rect 26158 8678 26210 8730
rect 26222 8678 26274 8730
rect 26286 8678 26338 8730
rect 26350 8678 26402 8730
rect 26414 8678 26466 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 1308 8440 1360 8492
rect 2320 8508 2372 8560
rect 2688 8576 2740 8628
rect 2688 8483 2740 8492
rect 2688 8449 2693 8483
rect 2693 8449 2727 8483
rect 2727 8449 2740 8483
rect 2688 8440 2740 8449
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 3332 8576 3384 8628
rect 4068 8576 4120 8628
rect 4252 8576 4304 8628
rect 2136 8304 2188 8356
rect 2228 8347 2280 8356
rect 2228 8313 2237 8347
rect 2237 8313 2271 8347
rect 2271 8313 2280 8347
rect 2228 8304 2280 8313
rect 3148 8304 3200 8356
rect 3792 8440 3844 8492
rect 4068 8440 4120 8492
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 4712 8440 4764 8492
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 7656 8576 7708 8628
rect 7748 8576 7800 8628
rect 8392 8576 8444 8628
rect 5816 8483 5868 8492
rect 5816 8449 5820 8483
rect 5820 8449 5854 8483
rect 5854 8449 5868 8483
rect 5816 8440 5868 8449
rect 3516 8415 3568 8424
rect 3516 8381 3525 8415
rect 3525 8381 3559 8415
rect 3559 8381 3568 8415
rect 3516 8372 3568 8381
rect 3700 8372 3752 8424
rect 2504 8236 2556 8288
rect 2872 8236 2924 8288
rect 3700 8279 3752 8288
rect 3700 8245 3709 8279
rect 3709 8245 3743 8279
rect 3743 8245 3752 8279
rect 3700 8236 3752 8245
rect 4068 8236 4120 8288
rect 4528 8236 4580 8288
rect 5632 8372 5684 8424
rect 4896 8347 4948 8356
rect 4896 8313 4905 8347
rect 4905 8313 4939 8347
rect 4939 8313 4948 8347
rect 4896 8304 4948 8313
rect 6276 8440 6328 8492
rect 6828 8440 6880 8492
rect 6644 8415 6696 8424
rect 6644 8381 6653 8415
rect 6653 8381 6687 8415
rect 6687 8381 6696 8415
rect 6644 8372 6696 8381
rect 7012 8372 7064 8424
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 7656 8372 7708 8424
rect 6920 8304 6972 8356
rect 8024 8440 8076 8492
rect 11060 8576 11112 8628
rect 13912 8576 13964 8628
rect 14740 8576 14792 8628
rect 15200 8576 15252 8628
rect 16488 8576 16540 8628
rect 17224 8576 17276 8628
rect 8760 8440 8812 8492
rect 9680 8372 9732 8424
rect 6828 8236 6880 8288
rect 15016 8508 15068 8560
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 12072 8483 12124 8492
rect 12072 8449 12081 8483
rect 12081 8449 12115 8483
rect 12115 8449 12124 8483
rect 12072 8440 12124 8449
rect 12348 8483 12400 8492
rect 12348 8449 12357 8483
rect 12357 8449 12391 8483
rect 12391 8449 12400 8483
rect 12348 8440 12400 8449
rect 12992 8440 13044 8492
rect 13176 8483 13228 8492
rect 13176 8449 13185 8483
rect 13185 8449 13219 8483
rect 13219 8449 13228 8483
rect 13176 8440 13228 8449
rect 13820 8440 13872 8492
rect 16580 8440 16632 8492
rect 16028 8415 16080 8424
rect 16028 8381 16037 8415
rect 16037 8381 16071 8415
rect 16071 8381 16080 8415
rect 16028 8372 16080 8381
rect 17132 8372 17184 8424
rect 17592 8508 17644 8560
rect 19064 8576 19116 8628
rect 19708 8508 19760 8560
rect 14740 8304 14792 8356
rect 18328 8372 18380 8424
rect 19248 8372 19300 8424
rect 18604 8304 18656 8356
rect 20812 8576 20864 8628
rect 21088 8576 21140 8628
rect 21824 8619 21876 8628
rect 21824 8585 21833 8619
rect 21833 8585 21867 8619
rect 21867 8585 21876 8619
rect 21824 8576 21876 8585
rect 21916 8576 21968 8628
rect 21272 8508 21324 8560
rect 23940 8576 23992 8628
rect 25688 8576 25740 8628
rect 23664 8440 23716 8492
rect 24216 8508 24268 8560
rect 23388 8372 23440 8424
rect 25136 8372 25188 8424
rect 11244 8279 11296 8288
rect 11244 8245 11253 8279
rect 11253 8245 11287 8279
rect 11287 8245 11296 8279
rect 11244 8236 11296 8245
rect 13268 8279 13320 8288
rect 13268 8245 13277 8279
rect 13277 8245 13311 8279
rect 13311 8245 13320 8279
rect 13268 8236 13320 8245
rect 14556 8236 14608 8288
rect 17224 8236 17276 8288
rect 21180 8279 21232 8288
rect 21180 8245 21189 8279
rect 21189 8245 21223 8279
rect 21223 8245 21232 8279
rect 21180 8236 21232 8245
rect 25228 8236 25280 8288
rect 4101 8134 4153 8186
rect 4165 8134 4217 8186
rect 4229 8134 4281 8186
rect 4293 8134 4345 8186
rect 4357 8134 4409 8186
rect 10403 8134 10455 8186
rect 10467 8134 10519 8186
rect 10531 8134 10583 8186
rect 10595 8134 10647 8186
rect 10659 8134 10711 8186
rect 16705 8134 16757 8186
rect 16769 8134 16821 8186
rect 16833 8134 16885 8186
rect 16897 8134 16949 8186
rect 16961 8134 17013 8186
rect 23007 8134 23059 8186
rect 23071 8134 23123 8186
rect 23135 8134 23187 8186
rect 23199 8134 23251 8186
rect 23263 8134 23315 8186
rect 2872 8075 2924 8084
rect 2872 8041 2881 8075
rect 2881 8041 2915 8075
rect 2915 8041 2924 8075
rect 2872 8032 2924 8041
rect 3148 8032 3200 8084
rect 3792 8032 3844 8084
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 7104 8032 7156 8084
rect 10876 8075 10928 8084
rect 10876 8041 10885 8075
rect 10885 8041 10919 8075
rect 10919 8041 10928 8075
rect 10876 8032 10928 8041
rect 11244 8032 11296 8084
rect 22560 8032 22612 8084
rect 7656 8007 7708 8016
rect 7656 7973 7665 8007
rect 7665 7973 7699 8007
rect 7699 7973 7708 8007
rect 7656 7964 7708 7973
rect 7748 7964 7800 8016
rect 2964 7828 3016 7880
rect 3332 7828 3384 7880
rect 3700 7828 3752 7880
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 5908 7760 5960 7812
rect 6092 7871 6144 7880
rect 6092 7837 6101 7871
rect 6101 7837 6135 7871
rect 6135 7837 6144 7871
rect 6092 7828 6144 7837
rect 6368 7828 6420 7880
rect 6460 7871 6512 7880
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 6552 7828 6604 7880
rect 3976 7735 4028 7744
rect 3976 7701 3985 7735
rect 3985 7701 4019 7735
rect 4019 7701 4028 7735
rect 3976 7692 4028 7701
rect 6276 7692 6328 7744
rect 8024 7828 8076 7880
rect 8760 7828 8812 7880
rect 13268 7964 13320 8016
rect 13820 7964 13872 8016
rect 12532 7896 12584 7948
rect 12900 7939 12952 7948
rect 12900 7905 12909 7939
rect 12909 7905 12943 7939
rect 12943 7905 12952 7939
rect 12900 7896 12952 7905
rect 13912 7896 13964 7948
rect 14556 7896 14608 7948
rect 17040 7939 17092 7948
rect 17040 7905 17049 7939
rect 17049 7905 17083 7939
rect 17083 7905 17092 7939
rect 17040 7896 17092 7905
rect 18512 7896 18564 7948
rect 21640 7939 21692 7948
rect 21640 7905 21649 7939
rect 21649 7905 21683 7939
rect 21683 7905 21692 7939
rect 21640 7896 21692 7905
rect 23664 7896 23716 7948
rect 24952 7939 25004 7948
rect 24952 7905 24961 7939
rect 24961 7905 24995 7939
rect 24995 7905 25004 7939
rect 24952 7896 25004 7905
rect 25320 7896 25372 7948
rect 25964 7939 26016 7948
rect 25964 7905 25973 7939
rect 25973 7905 26007 7939
rect 26007 7905 26016 7939
rect 25964 7896 26016 7905
rect 12072 7828 12124 7880
rect 11796 7760 11848 7812
rect 12716 7828 12768 7880
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 13268 7828 13320 7880
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 15660 7871 15712 7880
rect 15660 7837 15669 7871
rect 15669 7837 15703 7871
rect 15703 7837 15712 7871
rect 15660 7828 15712 7837
rect 16028 7871 16080 7880
rect 16028 7837 16037 7871
rect 16037 7837 16071 7871
rect 16071 7837 16080 7871
rect 16028 7828 16080 7837
rect 16488 7871 16540 7880
rect 16488 7837 16497 7871
rect 16497 7837 16531 7871
rect 16531 7837 16540 7871
rect 16488 7828 16540 7837
rect 8024 7692 8076 7744
rect 16580 7760 16632 7812
rect 19340 7828 19392 7880
rect 22192 7828 22244 7880
rect 14004 7692 14056 7744
rect 17224 7760 17276 7812
rect 17592 7760 17644 7812
rect 18052 7692 18104 7744
rect 19248 7735 19300 7744
rect 19248 7701 19257 7735
rect 19257 7701 19291 7735
rect 19291 7701 19300 7735
rect 19248 7692 19300 7701
rect 21272 7692 21324 7744
rect 21456 7692 21508 7744
rect 21916 7692 21968 7744
rect 22100 7735 22152 7744
rect 22100 7701 22109 7735
rect 22109 7701 22143 7735
rect 22143 7701 22152 7735
rect 22100 7692 22152 7701
rect 22284 7692 22336 7744
rect 24124 7692 24176 7744
rect 7252 7590 7304 7642
rect 7316 7590 7368 7642
rect 7380 7590 7432 7642
rect 7444 7590 7496 7642
rect 7508 7590 7560 7642
rect 13554 7590 13606 7642
rect 13618 7590 13670 7642
rect 13682 7590 13734 7642
rect 13746 7590 13798 7642
rect 13810 7590 13862 7642
rect 19856 7590 19908 7642
rect 19920 7590 19972 7642
rect 19984 7590 20036 7642
rect 20048 7590 20100 7642
rect 20112 7590 20164 7642
rect 26158 7590 26210 7642
rect 26222 7590 26274 7642
rect 26286 7590 26338 7642
rect 26350 7590 26402 7642
rect 26414 7590 26466 7642
rect 6920 7488 6972 7540
rect 7932 7488 7984 7540
rect 11612 7488 11664 7540
rect 14464 7488 14516 7540
rect 15108 7488 15160 7540
rect 16488 7488 16540 7540
rect 18696 7488 18748 7540
rect 6644 7420 6696 7472
rect 8024 7420 8076 7472
rect 6092 7352 6144 7404
rect 6368 7395 6420 7404
rect 6368 7361 6377 7395
rect 6377 7361 6411 7395
rect 6411 7361 6420 7395
rect 6368 7352 6420 7361
rect 6552 7284 6604 7336
rect 6828 7395 6880 7404
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 7748 7352 7800 7404
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8668 7352 8720 7361
rect 13176 7420 13228 7472
rect 9588 7352 9640 7404
rect 11704 7395 11756 7404
rect 11704 7361 11713 7395
rect 11713 7361 11747 7395
rect 11747 7361 11756 7395
rect 11704 7352 11756 7361
rect 11796 7352 11848 7404
rect 12440 7352 12492 7404
rect 12992 7352 13044 7404
rect 14004 7352 14056 7404
rect 14372 7352 14424 7404
rect 9404 7284 9456 7336
rect 12532 7284 12584 7336
rect 15660 7395 15712 7404
rect 15660 7361 15669 7395
rect 15669 7361 15703 7395
rect 15703 7361 15712 7395
rect 15660 7352 15712 7361
rect 17592 7420 17644 7472
rect 19248 7488 19300 7540
rect 20720 7531 20772 7540
rect 20720 7497 20729 7531
rect 20729 7497 20763 7531
rect 20763 7497 20772 7531
rect 20720 7488 20772 7497
rect 21824 7488 21876 7540
rect 21364 7420 21416 7472
rect 21732 7420 21784 7472
rect 23020 7420 23072 7472
rect 24124 7488 24176 7540
rect 25412 7531 25464 7540
rect 25412 7497 25421 7531
rect 25421 7497 25455 7531
rect 25455 7497 25464 7531
rect 25412 7488 25464 7497
rect 25228 7420 25280 7472
rect 17224 7352 17276 7404
rect 17316 7395 17368 7404
rect 17316 7361 17325 7395
rect 17325 7361 17359 7395
rect 17359 7361 17368 7395
rect 17316 7352 17368 7361
rect 16580 7284 16632 7336
rect 21640 7352 21692 7404
rect 16488 7216 16540 7268
rect 11888 7148 11940 7200
rect 14004 7148 14056 7200
rect 15016 7191 15068 7200
rect 15016 7157 15025 7191
rect 15025 7157 15059 7191
rect 15059 7157 15068 7191
rect 15016 7148 15068 7157
rect 15292 7191 15344 7200
rect 15292 7157 15301 7191
rect 15301 7157 15335 7191
rect 15335 7157 15344 7191
rect 15292 7148 15344 7157
rect 17132 7148 17184 7200
rect 18328 7148 18380 7200
rect 22008 7284 22060 7336
rect 23664 7327 23716 7336
rect 23664 7293 23673 7327
rect 23673 7293 23707 7327
rect 23707 7293 23716 7327
rect 23664 7284 23716 7293
rect 22284 7148 22336 7200
rect 4101 7046 4153 7098
rect 4165 7046 4217 7098
rect 4229 7046 4281 7098
rect 4293 7046 4345 7098
rect 4357 7046 4409 7098
rect 10403 7046 10455 7098
rect 10467 7046 10519 7098
rect 10531 7046 10583 7098
rect 10595 7046 10647 7098
rect 10659 7046 10711 7098
rect 16705 7046 16757 7098
rect 16769 7046 16821 7098
rect 16833 7046 16885 7098
rect 16897 7046 16949 7098
rect 16961 7046 17013 7098
rect 23007 7046 23059 7098
rect 23071 7046 23123 7098
rect 23135 7046 23187 7098
rect 23199 7046 23251 7098
rect 23263 7046 23315 7098
rect 5908 6987 5960 6996
rect 5908 6953 5917 6987
rect 5917 6953 5951 6987
rect 5951 6953 5960 6987
rect 5908 6944 5960 6953
rect 6644 6944 6696 6996
rect 11888 6944 11940 6996
rect 12716 6944 12768 6996
rect 13912 6944 13964 6996
rect 3056 6808 3108 6860
rect 12900 6876 12952 6928
rect 10876 6851 10928 6860
rect 10876 6817 10885 6851
rect 10885 6817 10919 6851
rect 10919 6817 10928 6851
rect 10876 6808 10928 6817
rect 3148 6740 3200 6792
rect 5816 6740 5868 6792
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 6460 6740 6512 6792
rect 8300 6783 8352 6792
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 5724 6672 5776 6724
rect 7012 6672 7064 6724
rect 7840 6672 7892 6724
rect 8484 6783 8536 6792
rect 8484 6749 8493 6783
rect 8493 6749 8527 6783
rect 8527 6749 8536 6783
rect 8484 6740 8536 6749
rect 9404 6783 9456 6792
rect 9404 6749 9413 6783
rect 9413 6749 9447 6783
rect 9447 6749 9456 6783
rect 9404 6740 9456 6749
rect 9588 6783 9640 6792
rect 9588 6749 9597 6783
rect 9597 6749 9631 6783
rect 9631 6749 9640 6783
rect 9588 6740 9640 6749
rect 10140 6740 10192 6792
rect 8668 6672 8720 6724
rect 1952 6604 2004 6656
rect 6644 6604 6696 6656
rect 9404 6604 9456 6656
rect 12164 6672 12216 6724
rect 12992 6740 13044 6792
rect 14004 6740 14056 6792
rect 14372 6919 14424 6928
rect 14372 6885 14381 6919
rect 14381 6885 14415 6919
rect 14415 6885 14424 6919
rect 14372 6876 14424 6885
rect 21732 6987 21784 6996
rect 21732 6953 21741 6987
rect 21741 6953 21775 6987
rect 21775 6953 21784 6987
rect 21732 6944 21784 6953
rect 22744 6944 22796 6996
rect 22376 6919 22428 6928
rect 22376 6885 22385 6919
rect 22385 6885 22419 6919
rect 22419 6885 22428 6919
rect 22376 6876 22428 6885
rect 22928 6876 22980 6928
rect 15108 6851 15160 6860
rect 15108 6817 15117 6851
rect 15117 6817 15151 6851
rect 15151 6817 15160 6851
rect 15108 6808 15160 6817
rect 15660 6808 15712 6860
rect 12532 6604 12584 6656
rect 12808 6604 12860 6656
rect 14648 6672 14700 6724
rect 16580 6808 16632 6860
rect 17500 6808 17552 6860
rect 23848 6944 23900 6996
rect 25136 6987 25188 6996
rect 25136 6953 25145 6987
rect 25145 6953 25179 6987
rect 25179 6953 25188 6987
rect 25136 6944 25188 6953
rect 23112 6876 23164 6928
rect 25412 6808 25464 6860
rect 18788 6783 18840 6792
rect 18788 6749 18797 6783
rect 18797 6749 18831 6783
rect 18831 6749 18840 6783
rect 18788 6740 18840 6749
rect 21916 6783 21968 6792
rect 21916 6749 21925 6783
rect 21925 6749 21959 6783
rect 21959 6749 21968 6783
rect 21916 6740 21968 6749
rect 22100 6783 22152 6792
rect 22100 6749 22124 6783
rect 22124 6749 22152 6783
rect 22100 6740 22152 6749
rect 22192 6783 22244 6792
rect 22192 6749 22201 6783
rect 22201 6749 22235 6783
rect 22235 6749 22244 6783
rect 22192 6740 22244 6749
rect 22284 6783 22336 6792
rect 22284 6749 22293 6783
rect 22293 6749 22327 6783
rect 22327 6749 22336 6783
rect 22284 6740 22336 6749
rect 22928 6740 22980 6792
rect 23112 6740 23164 6792
rect 22560 6672 22612 6724
rect 15936 6604 15988 6656
rect 16948 6604 17000 6656
rect 17040 6604 17092 6656
rect 17408 6647 17460 6656
rect 17408 6613 17417 6647
rect 17417 6613 17451 6647
rect 17451 6613 17460 6647
rect 17408 6604 17460 6613
rect 17960 6604 18012 6656
rect 18604 6647 18656 6656
rect 18604 6613 18613 6647
rect 18613 6613 18647 6647
rect 18647 6613 18656 6647
rect 18604 6604 18656 6613
rect 21916 6604 21968 6656
rect 23848 6604 23900 6656
rect 7252 6502 7304 6554
rect 7316 6502 7368 6554
rect 7380 6502 7432 6554
rect 7444 6502 7496 6554
rect 7508 6502 7560 6554
rect 13554 6502 13606 6554
rect 13618 6502 13670 6554
rect 13682 6502 13734 6554
rect 13746 6502 13798 6554
rect 13810 6502 13862 6554
rect 19856 6502 19908 6554
rect 19920 6502 19972 6554
rect 19984 6502 20036 6554
rect 20048 6502 20100 6554
rect 20112 6502 20164 6554
rect 26158 6502 26210 6554
rect 26222 6502 26274 6554
rect 26286 6502 26338 6554
rect 26350 6502 26402 6554
rect 26414 6502 26466 6554
rect 1952 6400 2004 6452
rect 6092 6400 6144 6452
rect 6552 6443 6604 6452
rect 6552 6409 6561 6443
rect 6561 6409 6595 6443
rect 6595 6409 6604 6443
rect 6552 6400 6604 6409
rect 8300 6400 8352 6452
rect 8484 6400 8536 6452
rect 11336 6400 11388 6452
rect 11888 6400 11940 6452
rect 12440 6443 12492 6452
rect 12440 6409 12449 6443
rect 12449 6409 12483 6443
rect 12483 6409 12492 6443
rect 12440 6400 12492 6409
rect 12992 6400 13044 6452
rect 14004 6400 14056 6452
rect 16948 6443 17000 6452
rect 16948 6409 16957 6443
rect 16957 6409 16991 6443
rect 16991 6409 17000 6443
rect 16948 6400 17000 6409
rect 17408 6400 17460 6452
rect 17500 6400 17552 6452
rect 19524 6400 19576 6452
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 2780 6264 2832 6316
rect 3424 6264 3476 6316
rect 5632 6264 5684 6316
rect 5264 6239 5316 6248
rect 5264 6205 5273 6239
rect 5273 6205 5307 6239
rect 5307 6205 5316 6239
rect 5264 6196 5316 6205
rect 6920 6239 6972 6248
rect 6920 6205 6929 6239
rect 6929 6205 6963 6239
rect 6963 6205 6972 6239
rect 6920 6196 6972 6205
rect 5816 6128 5868 6180
rect 3148 6103 3200 6112
rect 3148 6069 3157 6103
rect 3157 6069 3191 6103
rect 3191 6069 3200 6103
rect 3148 6060 3200 6069
rect 6184 6060 6236 6112
rect 8116 6060 8168 6112
rect 9404 6332 9456 6384
rect 12900 6332 12952 6384
rect 10324 6264 10376 6316
rect 10876 6196 10928 6248
rect 11888 6239 11940 6248
rect 11888 6205 11897 6239
rect 11897 6205 11931 6239
rect 11931 6205 11940 6239
rect 11888 6196 11940 6205
rect 14004 6264 14056 6316
rect 16120 6332 16172 6384
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 8852 6128 8904 6180
rect 8944 6060 8996 6112
rect 10324 6060 10376 6112
rect 14464 6239 14516 6248
rect 14464 6205 14473 6239
rect 14473 6205 14507 6239
rect 14507 6205 14516 6239
rect 14464 6196 14516 6205
rect 13912 6128 13964 6180
rect 15292 6307 15344 6316
rect 15292 6273 15301 6307
rect 15301 6273 15335 6307
rect 15335 6273 15344 6307
rect 15292 6264 15344 6273
rect 17040 6264 17092 6316
rect 18052 6375 18104 6384
rect 18052 6341 18061 6375
rect 18061 6341 18095 6375
rect 18095 6341 18104 6375
rect 18052 6332 18104 6341
rect 19064 6332 19116 6384
rect 18328 6307 18380 6316
rect 18328 6273 18337 6307
rect 18337 6273 18371 6307
rect 18371 6273 18380 6307
rect 18328 6264 18380 6273
rect 22376 6400 22428 6452
rect 23664 6400 23716 6452
rect 22836 6332 22888 6384
rect 23664 6264 23716 6316
rect 18604 6239 18656 6248
rect 18604 6205 18613 6239
rect 18613 6205 18647 6239
rect 18647 6205 18656 6239
rect 18604 6196 18656 6205
rect 14096 6060 14148 6112
rect 14280 6103 14332 6112
rect 14280 6069 14289 6103
rect 14289 6069 14323 6103
rect 14323 6069 14332 6103
rect 14280 6060 14332 6069
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 16580 6060 16632 6112
rect 17960 6128 18012 6180
rect 22008 6128 22060 6180
rect 21272 6060 21324 6112
rect 21548 6103 21600 6112
rect 21548 6069 21557 6103
rect 21557 6069 21591 6103
rect 21591 6069 21600 6103
rect 21548 6060 21600 6069
rect 22192 6060 22244 6112
rect 25136 6239 25188 6248
rect 25136 6205 25145 6239
rect 25145 6205 25179 6239
rect 25179 6205 25188 6239
rect 25136 6196 25188 6205
rect 23572 6128 23624 6180
rect 22836 6060 22888 6112
rect 23480 6060 23532 6112
rect 4101 5958 4153 6010
rect 4165 5958 4217 6010
rect 4229 5958 4281 6010
rect 4293 5958 4345 6010
rect 4357 5958 4409 6010
rect 10403 5958 10455 6010
rect 10467 5958 10519 6010
rect 10531 5958 10583 6010
rect 10595 5958 10647 6010
rect 10659 5958 10711 6010
rect 16705 5958 16757 6010
rect 16769 5958 16821 6010
rect 16833 5958 16885 6010
rect 16897 5958 16949 6010
rect 16961 5958 17013 6010
rect 23007 5958 23059 6010
rect 23071 5958 23123 6010
rect 23135 5958 23187 6010
rect 23199 5958 23251 6010
rect 23263 5958 23315 6010
rect 5264 5899 5316 5908
rect 5264 5865 5273 5899
rect 5273 5865 5307 5899
rect 5307 5865 5316 5899
rect 5264 5856 5316 5865
rect 6920 5856 6972 5908
rect 8116 5856 8168 5908
rect 8944 5899 8996 5908
rect 8944 5865 8953 5899
rect 8953 5865 8987 5899
rect 8987 5865 8996 5899
rect 8944 5856 8996 5865
rect 9128 5899 9180 5908
rect 9128 5865 9137 5899
rect 9137 5865 9171 5899
rect 9171 5865 9180 5899
rect 9128 5856 9180 5865
rect 5724 5788 5776 5840
rect 5540 5763 5592 5772
rect 5540 5729 5549 5763
rect 5549 5729 5583 5763
rect 5583 5729 5592 5763
rect 5540 5720 5592 5729
rect 5908 5720 5960 5772
rect 6184 5652 6236 5704
rect 6460 5763 6512 5772
rect 6460 5729 6469 5763
rect 6469 5729 6503 5763
rect 6503 5729 6512 5763
rect 6460 5720 6512 5729
rect 9680 5788 9732 5840
rect 10140 5899 10192 5908
rect 10140 5865 10149 5899
rect 10149 5865 10183 5899
rect 10183 5865 10192 5899
rect 10140 5856 10192 5865
rect 11612 5899 11664 5908
rect 11612 5865 11621 5899
rect 11621 5865 11655 5899
rect 11655 5865 11664 5899
rect 11612 5856 11664 5865
rect 9496 5720 9548 5772
rect 10048 5720 10100 5772
rect 6644 5652 6696 5704
rect 6736 5695 6788 5704
rect 6736 5661 6745 5695
rect 6745 5661 6779 5695
rect 6779 5661 6788 5695
rect 6736 5652 6788 5661
rect 6276 5584 6328 5636
rect 9220 5652 9272 5704
rect 9680 5652 9732 5704
rect 10692 5763 10744 5772
rect 10692 5729 10701 5763
rect 10701 5729 10735 5763
rect 10735 5729 10744 5763
rect 10692 5720 10744 5729
rect 12808 5856 12860 5908
rect 14004 5856 14056 5908
rect 15568 5856 15620 5908
rect 15936 5899 15988 5908
rect 15936 5865 15945 5899
rect 15945 5865 15979 5899
rect 15979 5865 15988 5899
rect 15936 5856 15988 5865
rect 18788 5856 18840 5908
rect 22560 5856 22612 5908
rect 12532 5720 12584 5772
rect 7012 5516 7064 5568
rect 8116 5516 8168 5568
rect 8944 5516 8996 5568
rect 9220 5516 9272 5568
rect 9588 5516 9640 5568
rect 9680 5516 9732 5568
rect 9956 5516 10008 5568
rect 10784 5652 10836 5704
rect 17040 5720 17092 5772
rect 10324 5516 10376 5568
rect 13176 5652 13228 5704
rect 15936 5652 15988 5704
rect 17868 5652 17920 5704
rect 18052 5763 18104 5772
rect 18052 5729 18086 5763
rect 18086 5729 18104 5763
rect 18052 5720 18104 5729
rect 18512 5763 18564 5772
rect 18512 5729 18521 5763
rect 18521 5729 18555 5763
rect 18555 5729 18564 5763
rect 18512 5720 18564 5729
rect 18972 5720 19024 5772
rect 18696 5652 18748 5704
rect 18788 5652 18840 5704
rect 19524 5720 19576 5772
rect 19616 5720 19668 5772
rect 21548 5720 21600 5772
rect 23664 5720 23716 5772
rect 18420 5584 18472 5636
rect 17592 5516 17644 5568
rect 17960 5516 18012 5568
rect 18236 5559 18288 5568
rect 18236 5525 18245 5559
rect 18245 5525 18279 5559
rect 18279 5525 18288 5559
rect 18236 5516 18288 5525
rect 18696 5559 18748 5568
rect 18696 5525 18705 5559
rect 18705 5525 18739 5559
rect 18739 5525 18748 5559
rect 18696 5516 18748 5525
rect 19064 5559 19116 5568
rect 19064 5525 19073 5559
rect 19073 5525 19107 5559
rect 19107 5525 19116 5559
rect 19064 5516 19116 5525
rect 22744 5652 22796 5704
rect 21272 5516 21324 5568
rect 22100 5516 22152 5568
rect 7252 5414 7304 5466
rect 7316 5414 7368 5466
rect 7380 5414 7432 5466
rect 7444 5414 7496 5466
rect 7508 5414 7560 5466
rect 13554 5414 13606 5466
rect 13618 5414 13670 5466
rect 13682 5414 13734 5466
rect 13746 5414 13798 5466
rect 13810 5414 13862 5466
rect 19856 5414 19908 5466
rect 19920 5414 19972 5466
rect 19984 5414 20036 5466
rect 20048 5414 20100 5466
rect 20112 5414 20164 5466
rect 26158 5414 26210 5466
rect 26222 5414 26274 5466
rect 26286 5414 26338 5466
rect 26350 5414 26402 5466
rect 26414 5414 26466 5466
rect 5540 5355 5592 5364
rect 5540 5321 5549 5355
rect 5549 5321 5583 5355
rect 5583 5321 5592 5355
rect 5540 5312 5592 5321
rect 5632 5355 5684 5364
rect 5632 5321 5641 5355
rect 5641 5321 5675 5355
rect 5675 5321 5684 5355
rect 5632 5312 5684 5321
rect 6184 5312 6236 5364
rect 8116 5355 8168 5364
rect 8116 5321 8125 5355
rect 8125 5321 8159 5355
rect 8159 5321 8168 5355
rect 8116 5312 8168 5321
rect 3976 5108 4028 5160
rect 5632 5176 5684 5228
rect 6736 5287 6788 5296
rect 6736 5253 6745 5287
rect 6745 5253 6779 5287
rect 6779 5253 6788 5287
rect 6736 5244 6788 5253
rect 6092 5219 6144 5228
rect 6092 5185 6101 5219
rect 6101 5185 6135 5219
rect 6135 5185 6144 5219
rect 6092 5176 6144 5185
rect 7012 5176 7064 5228
rect 8852 5244 8904 5296
rect 9220 5312 9272 5364
rect 9496 5312 9548 5364
rect 9680 5312 9732 5364
rect 11612 5312 11664 5364
rect 13268 5312 13320 5364
rect 6276 5108 6328 5160
rect 9036 5176 9088 5228
rect 9772 5244 9824 5296
rect 10692 5244 10744 5296
rect 9312 5219 9364 5228
rect 9312 5185 9321 5219
rect 9321 5185 9355 5219
rect 9355 5185 9364 5219
rect 9312 5176 9364 5185
rect 9680 5217 9732 5228
rect 9680 5183 9689 5217
rect 9689 5183 9723 5217
rect 9723 5183 9732 5217
rect 9680 5176 9732 5183
rect 9956 5176 10008 5228
rect 9864 5108 9916 5160
rect 12992 5176 13044 5228
rect 13268 5219 13320 5228
rect 13268 5185 13277 5219
rect 13277 5185 13311 5219
rect 13311 5185 13320 5219
rect 13268 5176 13320 5185
rect 14280 5244 14332 5296
rect 16580 5312 16632 5364
rect 17592 5355 17644 5364
rect 17592 5321 17601 5355
rect 17601 5321 17635 5355
rect 17635 5321 17644 5355
rect 17592 5312 17644 5321
rect 18696 5312 18748 5364
rect 23480 5355 23532 5364
rect 23480 5321 23489 5355
rect 23489 5321 23523 5355
rect 23523 5321 23532 5355
rect 23480 5312 23532 5321
rect 11428 5040 11480 5092
rect 8852 5015 8904 5024
rect 8852 4981 8861 5015
rect 8861 4981 8895 5015
rect 8895 4981 8904 5015
rect 8852 4972 8904 4981
rect 8944 4972 8996 5024
rect 12624 4972 12676 5024
rect 12716 4972 12768 5024
rect 17040 5219 17092 5228
rect 17040 5185 17049 5219
rect 17049 5185 17083 5219
rect 17083 5185 17092 5219
rect 17040 5176 17092 5185
rect 17868 5176 17920 5228
rect 18420 5287 18472 5296
rect 18420 5253 18429 5287
rect 18429 5253 18463 5287
rect 18463 5253 18472 5287
rect 18420 5244 18472 5253
rect 21272 5244 21324 5296
rect 18144 5219 18196 5228
rect 18144 5185 18153 5219
rect 18153 5185 18187 5219
rect 18187 5185 18196 5219
rect 18144 5176 18196 5185
rect 18328 5108 18380 5160
rect 18144 5040 18196 5092
rect 18236 5040 18288 5092
rect 13084 4972 13136 5024
rect 13360 5015 13412 5024
rect 13360 4981 13369 5015
rect 13369 4981 13403 5015
rect 13403 4981 13412 5015
rect 13360 4972 13412 4981
rect 17040 4972 17092 5024
rect 18972 5108 19024 5160
rect 22560 5108 22612 5160
rect 18880 4972 18932 5024
rect 4101 4870 4153 4922
rect 4165 4870 4217 4922
rect 4229 4870 4281 4922
rect 4293 4870 4345 4922
rect 4357 4870 4409 4922
rect 10403 4870 10455 4922
rect 10467 4870 10519 4922
rect 10531 4870 10583 4922
rect 10595 4870 10647 4922
rect 10659 4870 10711 4922
rect 16705 4870 16757 4922
rect 16769 4870 16821 4922
rect 16833 4870 16885 4922
rect 16897 4870 16949 4922
rect 16961 4870 17013 4922
rect 23007 4870 23059 4922
rect 23071 4870 23123 4922
rect 23135 4870 23187 4922
rect 23199 4870 23251 4922
rect 23263 4870 23315 4922
rect 5816 4811 5868 4820
rect 5816 4777 5825 4811
rect 5825 4777 5859 4811
rect 5859 4777 5868 4811
rect 5816 4768 5868 4777
rect 6092 4811 6144 4820
rect 6092 4777 6101 4811
rect 6101 4777 6135 4811
rect 6135 4777 6144 4811
rect 6092 4768 6144 4777
rect 7012 4811 7064 4820
rect 7012 4777 7021 4811
rect 7021 4777 7055 4811
rect 7055 4777 7064 4811
rect 7012 4768 7064 4777
rect 8944 4768 8996 4820
rect 9128 4768 9180 4820
rect 9312 4768 9364 4820
rect 9496 4811 9548 4820
rect 9496 4777 9505 4811
rect 9505 4777 9539 4811
rect 9539 4777 9548 4811
rect 9496 4768 9548 4777
rect 10048 4768 10100 4820
rect 5632 4700 5684 4752
rect 3148 4564 3200 4616
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 5908 4607 5960 4616
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 6276 4632 6328 4684
rect 8852 4632 8904 4684
rect 9772 4675 9824 4684
rect 9772 4641 9781 4675
rect 9781 4641 9815 4675
rect 9815 4641 9824 4675
rect 9772 4632 9824 4641
rect 11336 4768 11388 4820
rect 11428 4768 11480 4820
rect 12900 4768 12952 4820
rect 13544 4768 13596 4820
rect 13912 4768 13964 4820
rect 14004 4768 14056 4820
rect 16764 4700 16816 4752
rect 10876 4632 10928 4684
rect 12992 4632 13044 4684
rect 13544 4632 13596 4684
rect 940 4496 992 4548
rect 7104 4607 7156 4616
rect 7104 4573 7113 4607
rect 7113 4573 7147 4607
rect 7147 4573 7156 4607
rect 7104 4564 7156 4573
rect 9404 4564 9456 4616
rect 12164 4564 12216 4616
rect 13360 4564 13412 4616
rect 7656 4428 7708 4480
rect 9680 4428 9732 4480
rect 10416 4471 10468 4480
rect 10416 4437 10425 4471
rect 10425 4437 10459 4471
rect 10459 4437 10468 4471
rect 10416 4428 10468 4437
rect 11152 4496 11204 4548
rect 12348 4471 12400 4480
rect 12348 4437 12357 4471
rect 12357 4437 12391 4471
rect 12391 4437 12400 4471
rect 12348 4428 12400 4437
rect 16028 4632 16080 4684
rect 18788 4768 18840 4820
rect 18972 4768 19024 4820
rect 17040 4632 17092 4684
rect 18052 4564 18104 4616
rect 19064 4607 19116 4616
rect 19064 4573 19073 4607
rect 19073 4573 19107 4607
rect 19107 4573 19116 4607
rect 19064 4564 19116 4573
rect 17776 4496 17828 4548
rect 15200 4428 15252 4480
rect 15936 4471 15988 4480
rect 15936 4437 15945 4471
rect 15945 4437 15979 4471
rect 15979 4437 15988 4471
rect 15936 4428 15988 4437
rect 16764 4428 16816 4480
rect 25964 4428 26016 4480
rect 7252 4326 7304 4378
rect 7316 4326 7368 4378
rect 7380 4326 7432 4378
rect 7444 4326 7496 4378
rect 7508 4326 7560 4378
rect 13554 4326 13606 4378
rect 13618 4326 13670 4378
rect 13682 4326 13734 4378
rect 13746 4326 13798 4378
rect 13810 4326 13862 4378
rect 19856 4326 19908 4378
rect 19920 4326 19972 4378
rect 19984 4326 20036 4378
rect 20048 4326 20100 4378
rect 20112 4326 20164 4378
rect 26158 4326 26210 4378
rect 26222 4326 26274 4378
rect 26286 4326 26338 4378
rect 26350 4326 26402 4378
rect 26414 4326 26466 4378
rect 6276 4224 6328 4276
rect 7656 4224 7708 4276
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 9312 4156 9364 4208
rect 10416 4224 10468 4276
rect 10784 4224 10836 4276
rect 11152 4224 11204 4276
rect 13084 4224 13136 4276
rect 13636 4267 13688 4276
rect 13636 4233 13645 4267
rect 13645 4233 13679 4267
rect 13679 4233 13688 4267
rect 13636 4224 13688 4233
rect 9680 4199 9732 4208
rect 9680 4165 9689 4199
rect 9689 4165 9723 4199
rect 9723 4165 9732 4199
rect 9680 4156 9732 4165
rect 10232 4156 10284 4208
rect 10048 4131 10100 4140
rect 10048 4097 10057 4131
rect 10057 4097 10091 4131
rect 10091 4097 10100 4131
rect 10048 4088 10100 4097
rect 7932 4063 7984 4072
rect 7932 4029 7941 4063
rect 7941 4029 7975 4063
rect 7975 4029 7984 4063
rect 7932 4020 7984 4029
rect 10232 4020 10284 4072
rect 9404 3995 9456 4004
rect 9404 3961 9413 3995
rect 9413 3961 9447 3995
rect 9447 3961 9456 3995
rect 9404 3952 9456 3961
rect 10140 3927 10192 3936
rect 10140 3893 10149 3927
rect 10149 3893 10183 3927
rect 10183 3893 10192 3927
rect 10140 3884 10192 3893
rect 13176 4199 13228 4208
rect 13176 4165 13185 4199
rect 13185 4165 13219 4199
rect 13219 4165 13228 4199
rect 13176 4156 13228 4165
rect 16120 4156 16172 4208
rect 21272 4156 21324 4208
rect 11980 4131 12032 4140
rect 11980 4097 11989 4131
rect 11989 4097 12023 4131
rect 12023 4097 12032 4131
rect 11980 4088 12032 4097
rect 12716 4088 12768 4140
rect 13452 4088 13504 4140
rect 12348 4063 12400 4072
rect 12348 4029 12357 4063
rect 12357 4029 12391 4063
rect 12391 4029 12400 4063
rect 12348 4020 12400 4029
rect 11888 3952 11940 4004
rect 17132 4131 17184 4140
rect 17132 4097 17141 4131
rect 17141 4097 17175 4131
rect 17175 4097 17184 4131
rect 17132 4088 17184 4097
rect 17776 4131 17828 4140
rect 17776 4097 17785 4131
rect 17785 4097 17819 4131
rect 17819 4097 17828 4131
rect 17776 4088 17828 4097
rect 17868 4131 17920 4140
rect 17868 4097 17877 4131
rect 17877 4097 17911 4131
rect 17911 4097 17920 4131
rect 17868 4088 17920 4097
rect 18052 4088 18104 4140
rect 23664 4088 23716 4140
rect 16028 4063 16080 4072
rect 16028 4029 16037 4063
rect 16037 4029 16071 4063
rect 16071 4029 16080 4063
rect 16028 4020 16080 4029
rect 11796 3927 11848 3936
rect 11796 3893 11805 3927
rect 11805 3893 11839 3927
rect 11839 3893 11848 3927
rect 11796 3884 11848 3893
rect 13268 3927 13320 3936
rect 13268 3893 13277 3927
rect 13277 3893 13311 3927
rect 13311 3893 13320 3927
rect 13268 3884 13320 3893
rect 15016 3927 15068 3936
rect 15016 3893 15025 3927
rect 15025 3893 15059 3927
rect 15059 3893 15068 3927
rect 15016 3884 15068 3893
rect 18512 4020 18564 4072
rect 22560 4020 22612 4072
rect 22836 4020 22888 4072
rect 16396 3884 16448 3936
rect 18236 3927 18288 3936
rect 18236 3893 18245 3927
rect 18245 3893 18279 3927
rect 18279 3893 18288 3927
rect 18236 3884 18288 3893
rect 4101 3782 4153 3834
rect 4165 3782 4217 3834
rect 4229 3782 4281 3834
rect 4293 3782 4345 3834
rect 4357 3782 4409 3834
rect 10403 3782 10455 3834
rect 10467 3782 10519 3834
rect 10531 3782 10583 3834
rect 10595 3782 10647 3834
rect 10659 3782 10711 3834
rect 16705 3782 16757 3834
rect 16769 3782 16821 3834
rect 16833 3782 16885 3834
rect 16897 3782 16949 3834
rect 16961 3782 17013 3834
rect 23007 3782 23059 3834
rect 23071 3782 23123 3834
rect 23135 3782 23187 3834
rect 23199 3782 23251 3834
rect 23263 3782 23315 3834
rect 7104 3680 7156 3732
rect 1400 3544 1452 3596
rect 7932 3680 7984 3732
rect 11796 3680 11848 3732
rect 12440 3680 12492 3732
rect 12992 3680 13044 3732
rect 13452 3680 13504 3732
rect 13636 3680 13688 3732
rect 11520 3612 11572 3664
rect 8024 3544 8076 3596
rect 9772 3544 9824 3596
rect 10232 3587 10284 3596
rect 10232 3553 10241 3587
rect 10241 3553 10275 3587
rect 10275 3553 10284 3587
rect 10232 3544 10284 3553
rect 10876 3544 10928 3596
rect 5908 3451 5960 3460
rect 5908 3417 5917 3451
rect 5917 3417 5951 3451
rect 5951 3417 5960 3451
rect 5908 3408 5960 3417
rect 3424 3340 3476 3392
rect 7656 3340 7708 3392
rect 9404 3476 9456 3528
rect 15200 3680 15252 3732
rect 15936 3680 15988 3732
rect 18052 3723 18104 3732
rect 18052 3689 18061 3723
rect 18061 3689 18095 3723
rect 18095 3689 18104 3723
rect 18052 3680 18104 3689
rect 22836 3680 22888 3732
rect 14372 3476 14424 3528
rect 18880 3544 18932 3596
rect 18236 3476 18288 3528
rect 11520 3340 11572 3392
rect 12348 3451 12400 3460
rect 12348 3417 12357 3451
rect 12357 3417 12391 3451
rect 12391 3417 12400 3451
rect 12348 3408 12400 3417
rect 12164 3340 12216 3392
rect 15200 3408 15252 3460
rect 16580 3451 16632 3460
rect 16580 3417 16589 3451
rect 16589 3417 16623 3451
rect 16623 3417 16632 3451
rect 16580 3408 16632 3417
rect 17040 3408 17092 3460
rect 20260 3408 20312 3460
rect 21272 3408 21324 3460
rect 18328 3383 18380 3392
rect 18328 3349 18337 3383
rect 18337 3349 18371 3383
rect 18371 3349 18380 3383
rect 18328 3340 18380 3349
rect 7252 3238 7304 3290
rect 7316 3238 7368 3290
rect 7380 3238 7432 3290
rect 7444 3238 7496 3290
rect 7508 3238 7560 3290
rect 13554 3238 13606 3290
rect 13618 3238 13670 3290
rect 13682 3238 13734 3290
rect 13746 3238 13798 3290
rect 13810 3238 13862 3290
rect 19856 3238 19908 3290
rect 19920 3238 19972 3290
rect 19984 3238 20036 3290
rect 20048 3238 20100 3290
rect 20112 3238 20164 3290
rect 26158 3238 26210 3290
rect 26222 3238 26274 3290
rect 26286 3238 26338 3290
rect 26350 3238 26402 3290
rect 26414 3238 26466 3290
rect 5908 3136 5960 3188
rect 7656 3136 7708 3188
rect 9680 3136 9732 3188
rect 9312 3068 9364 3120
rect 10140 3136 10192 3188
rect 11980 3136 12032 3188
rect 12348 3136 12400 3188
rect 13268 3136 13320 3188
rect 15016 3136 15068 3188
rect 16120 3179 16172 3188
rect 16120 3145 16129 3179
rect 16129 3145 16163 3179
rect 16163 3145 16172 3179
rect 16120 3136 16172 3145
rect 16396 3136 16448 3188
rect 16580 3136 16632 3188
rect 17868 3136 17920 3188
rect 18328 3136 18380 3188
rect 10232 3000 10284 3052
rect 8024 2932 8076 2984
rect 12440 3068 12492 3120
rect 15292 3068 15344 3120
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 17040 3068 17092 3120
rect 11888 2932 11940 2984
rect 18880 2975 18932 2984
rect 18880 2941 18889 2975
rect 18889 2941 18923 2975
rect 18923 2941 18932 2975
rect 18880 2932 18932 2941
rect 4101 2694 4153 2746
rect 4165 2694 4217 2746
rect 4229 2694 4281 2746
rect 4293 2694 4345 2746
rect 4357 2694 4409 2746
rect 10403 2694 10455 2746
rect 10467 2694 10519 2746
rect 10531 2694 10583 2746
rect 10595 2694 10647 2746
rect 10659 2694 10711 2746
rect 16705 2694 16757 2746
rect 16769 2694 16821 2746
rect 16833 2694 16885 2746
rect 16897 2694 16949 2746
rect 16961 2694 17013 2746
rect 23007 2694 23059 2746
rect 23071 2694 23123 2746
rect 23135 2694 23187 2746
rect 23199 2694 23251 2746
rect 23263 2694 23315 2746
rect 20260 2592 20312 2644
rect 25136 2592 25188 2644
rect 3516 2456 3568 2508
rect 2228 2388 2280 2440
rect 4896 2388 4948 2440
rect 14188 2388 14240 2440
rect 15936 2431 15988 2440
rect 15936 2397 15945 2431
rect 15945 2397 15979 2431
rect 15979 2397 15988 2431
rect 15936 2388 15988 2397
rect 20260 2431 20312 2440
rect 20260 2397 20269 2431
rect 20269 2397 20303 2431
rect 20303 2397 20312 2431
rect 20260 2388 20312 2397
rect 20 2320 72 2372
rect 3976 2363 4028 2372
rect 3976 2329 3985 2363
rect 3985 2329 4019 2363
rect 4019 2329 4028 2363
rect 3976 2320 4028 2329
rect 11704 2363 11756 2372
rect 11704 2329 11713 2363
rect 11713 2329 11747 2363
rect 11747 2329 11756 2363
rect 11704 2320 11756 2329
rect 15568 2363 15620 2372
rect 15568 2329 15577 2363
rect 15577 2329 15611 2363
rect 15611 2329 15620 2363
rect 15568 2320 15620 2329
rect 16396 2320 16448 2372
rect 7748 2252 7800 2304
rect 23848 2252 23900 2304
rect 24768 2252 24820 2304
rect 7252 2150 7304 2202
rect 7316 2150 7368 2202
rect 7380 2150 7432 2202
rect 7444 2150 7496 2202
rect 7508 2150 7560 2202
rect 13554 2150 13606 2202
rect 13618 2150 13670 2202
rect 13682 2150 13734 2202
rect 13746 2150 13798 2202
rect 13810 2150 13862 2202
rect 19856 2150 19908 2202
rect 19920 2150 19972 2202
rect 19984 2150 20036 2202
rect 20048 2150 20100 2202
rect 20112 2150 20164 2202
rect 26158 2150 26210 2202
rect 26222 2150 26274 2202
rect 26286 2150 26338 2202
rect 26350 2150 26402 2202
rect 26414 2150 26466 2202
<< metal2 >>
rect 2778 29336 2834 29345
rect 2778 29271 2834 29280
rect 2792 27130 2820 29271
rect 3238 28809 3294 29609
rect 7102 28809 7158 29609
rect 11610 28809 11666 29609
rect 15474 28914 15530 29609
rect 15474 28886 15792 28914
rect 15474 28809 15530 28886
rect 3252 27130 3280 28809
rect 7116 27130 7144 28809
rect 7252 27228 7560 27237
rect 7252 27226 7258 27228
rect 7314 27226 7338 27228
rect 7394 27226 7418 27228
rect 7474 27226 7498 27228
rect 7554 27226 7560 27228
rect 7314 27174 7316 27226
rect 7496 27174 7498 27226
rect 7252 27172 7258 27174
rect 7314 27172 7338 27174
rect 7394 27172 7418 27174
rect 7474 27172 7498 27174
rect 7554 27172 7560 27174
rect 7252 27163 7560 27172
rect 11624 27130 11652 28809
rect 13554 27228 13862 27237
rect 13554 27226 13560 27228
rect 13616 27226 13640 27228
rect 13696 27226 13720 27228
rect 13776 27226 13800 27228
rect 13856 27226 13862 27228
rect 13616 27174 13618 27226
rect 13798 27174 13800 27226
rect 13554 27172 13560 27174
rect 13616 27172 13640 27174
rect 13696 27172 13720 27174
rect 13776 27172 13800 27174
rect 13856 27172 13862 27174
rect 13554 27163 13862 27172
rect 15764 27130 15792 28886
rect 19338 28809 19394 29609
rect 23202 28914 23258 29609
rect 23202 28886 23428 28914
rect 23202 28809 23258 28886
rect 19352 27130 19380 28809
rect 23400 27554 23428 28886
rect 27066 28809 27122 29609
rect 23400 27526 23520 27554
rect 19856 27228 20164 27237
rect 19856 27226 19862 27228
rect 19918 27226 19942 27228
rect 19998 27226 20022 27228
rect 20078 27226 20102 27228
rect 20158 27226 20164 27228
rect 19918 27174 19920 27226
rect 20100 27174 20102 27226
rect 19856 27172 19862 27174
rect 19918 27172 19942 27174
rect 19998 27172 20022 27174
rect 20078 27172 20102 27174
rect 20158 27172 20164 27174
rect 19856 27163 20164 27172
rect 23492 27130 23520 27526
rect 26158 27228 26466 27237
rect 26158 27226 26164 27228
rect 26220 27226 26244 27228
rect 26300 27226 26324 27228
rect 26380 27226 26404 27228
rect 26460 27226 26466 27228
rect 26220 27174 26222 27226
rect 26402 27174 26404 27226
rect 26158 27172 26164 27174
rect 26220 27172 26244 27174
rect 26300 27172 26324 27174
rect 26380 27172 26404 27174
rect 26460 27172 26466 27174
rect 26158 27163 26466 27172
rect 2780 27124 2832 27130
rect 2780 27066 2832 27072
rect 3240 27124 3292 27130
rect 3240 27066 3292 27072
rect 7104 27124 7156 27130
rect 7104 27066 7156 27072
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 15200 27124 15252 27130
rect 15200 27066 15252 27072
rect 15752 27124 15804 27130
rect 15752 27066 15804 27072
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 23480 27124 23532 27130
rect 23480 27066 23532 27072
rect 13452 27056 13504 27062
rect 13452 26998 13504 27004
rect 1768 26988 1820 26994
rect 1768 26930 1820 26936
rect 5080 26988 5132 26994
rect 5080 26930 5132 26936
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 11336 26988 11388 26994
rect 11336 26930 11388 26936
rect 940 25288 992 25294
rect 938 25256 940 25265
rect 992 25256 994 25265
rect 938 25191 994 25200
rect 940 21344 992 21350
rect 940 21286 992 21292
rect 952 21185 980 21286
rect 938 21176 994 21185
rect 938 21111 994 21120
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 1596 19378 1624 19790
rect 1584 19372 1636 19378
rect 1584 19314 1636 19320
rect 1596 18834 1624 19314
rect 1584 18828 1636 18834
rect 1584 18770 1636 18776
rect 1584 17128 1636 17134
rect 1584 17070 1636 17076
rect 1492 16652 1544 16658
rect 1492 16594 1544 16600
rect 1504 16561 1532 16594
rect 1490 16552 1546 16561
rect 1490 16487 1546 16496
rect 1596 15570 1624 17070
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1596 15026 1624 15506
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1596 13258 1624 14962
rect 1584 13252 1636 13258
rect 1584 13194 1636 13200
rect 1676 13252 1728 13258
rect 1676 13194 1728 13200
rect 1596 12986 1624 13194
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1688 12866 1716 13194
rect 1596 12838 1716 12866
rect 938 12336 994 12345
rect 938 12271 994 12280
rect 952 12238 980 12271
rect 940 12232 992 12238
rect 940 12174 992 12180
rect 1400 12096 1452 12102
rect 1400 12038 1452 12044
rect 1412 11082 1440 12038
rect 1400 11076 1452 11082
rect 1400 11018 1452 11024
rect 1412 8974 1440 11018
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1308 8492 1360 8498
rect 1308 8434 1360 8440
rect 1320 8265 1348 8434
rect 1306 8256 1362 8265
rect 1306 8191 1362 8200
rect 1412 6322 1440 8910
rect 1596 8634 1624 12838
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1688 12442 1716 12718
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1780 9450 1808 26930
rect 4101 26684 4409 26693
rect 4101 26682 4107 26684
rect 4163 26682 4187 26684
rect 4243 26682 4267 26684
rect 4323 26682 4347 26684
rect 4403 26682 4409 26684
rect 4163 26630 4165 26682
rect 4345 26630 4347 26682
rect 4101 26628 4107 26630
rect 4163 26628 4187 26630
rect 4243 26628 4267 26630
rect 4323 26628 4347 26630
rect 4403 26628 4409 26630
rect 4101 26619 4409 26628
rect 4988 26240 5040 26246
rect 4988 26182 5040 26188
rect 4101 25596 4409 25605
rect 4101 25594 4107 25596
rect 4163 25594 4187 25596
rect 4243 25594 4267 25596
rect 4323 25594 4347 25596
rect 4403 25594 4409 25596
rect 4163 25542 4165 25594
rect 4345 25542 4347 25594
rect 4101 25540 4107 25542
rect 4163 25540 4187 25542
rect 4243 25540 4267 25542
rect 4323 25540 4347 25542
rect 4403 25540 4409 25542
rect 4101 25531 4409 25540
rect 5000 25294 5028 26182
rect 4436 25288 4488 25294
rect 4436 25230 4488 25236
rect 4988 25288 5040 25294
rect 4988 25230 5040 25236
rect 4448 24750 4476 25230
rect 4436 24744 4488 24750
rect 4436 24686 4488 24692
rect 4712 24744 4764 24750
rect 4712 24686 4764 24692
rect 4101 24508 4409 24517
rect 4101 24506 4107 24508
rect 4163 24506 4187 24508
rect 4243 24506 4267 24508
rect 4323 24506 4347 24508
rect 4403 24506 4409 24508
rect 4163 24454 4165 24506
rect 4345 24454 4347 24506
rect 4101 24452 4107 24454
rect 4163 24452 4187 24454
rect 4243 24452 4267 24454
rect 4323 24452 4347 24454
rect 4403 24452 4409 24454
rect 4101 24443 4409 24452
rect 4448 24070 4476 24686
rect 4436 24064 4488 24070
rect 4436 24006 4488 24012
rect 4101 23420 4409 23429
rect 4101 23418 4107 23420
rect 4163 23418 4187 23420
rect 4243 23418 4267 23420
rect 4323 23418 4347 23420
rect 4403 23418 4409 23420
rect 4163 23366 4165 23418
rect 4345 23366 4347 23418
rect 4101 23364 4107 23366
rect 4163 23364 4187 23366
rect 4243 23364 4267 23366
rect 4323 23364 4347 23366
rect 4403 23364 4409 23366
rect 4101 23355 4409 23364
rect 4448 23186 4476 24006
rect 4724 23866 4752 24686
rect 4712 23860 4764 23866
rect 4712 23802 4764 23808
rect 4712 23656 4764 23662
rect 4712 23598 4764 23604
rect 4988 23656 5040 23662
rect 4988 23598 5040 23604
rect 4528 23520 4580 23526
rect 4528 23462 4580 23468
rect 4436 23180 4488 23186
rect 4436 23122 4488 23128
rect 4540 22982 4568 23462
rect 4528 22976 4580 22982
rect 4528 22918 4580 22924
rect 3148 22772 3200 22778
rect 3148 22714 3200 22720
rect 2688 22568 2740 22574
rect 2688 22510 2740 22516
rect 2700 21622 2728 22510
rect 3160 21622 3188 22714
rect 4724 22574 4752 23598
rect 5000 22642 5028 23598
rect 4988 22636 5040 22642
rect 4988 22578 5040 22584
rect 3516 22568 3568 22574
rect 3516 22510 3568 22516
rect 4712 22568 4764 22574
rect 4712 22510 4764 22516
rect 2688 21616 2740 21622
rect 2688 21558 2740 21564
rect 3148 21616 3200 21622
rect 3148 21558 3200 21564
rect 1952 21548 2004 21554
rect 1952 21490 2004 21496
rect 1860 18692 1912 18698
rect 1860 18634 1912 18640
rect 1872 18426 1900 18634
rect 1860 18420 1912 18426
rect 1860 18362 1912 18368
rect 1964 18154 1992 21490
rect 2136 20256 2188 20262
rect 2136 20198 2188 20204
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 2148 19446 2176 20198
rect 2424 19922 2452 20198
rect 2412 19916 2464 19922
rect 2412 19858 2464 19864
rect 2700 19514 2728 21558
rect 3056 21480 3108 21486
rect 3056 21422 3108 21428
rect 3068 21146 3096 21422
rect 3056 21140 3108 21146
rect 3056 21082 3108 21088
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2792 19514 2820 20334
rect 3160 19786 3188 21558
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 3148 19780 3200 19786
rect 3148 19722 3200 19728
rect 2688 19508 2740 19514
rect 2688 19450 2740 19456
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 2136 19440 2188 19446
rect 2136 19382 2188 19388
rect 3160 19378 3188 19722
rect 3344 19446 3372 20334
rect 3332 19440 3384 19446
rect 3332 19382 3384 19388
rect 3148 19372 3200 19378
rect 3200 19320 3280 19334
rect 3148 19314 3280 19320
rect 3160 19306 3280 19314
rect 3252 18698 3280 19306
rect 3240 18692 3292 18698
rect 3240 18634 3292 18640
rect 1952 18148 2004 18154
rect 1952 18090 2004 18096
rect 3252 17202 3280 18634
rect 3528 18426 3556 22510
rect 4101 22332 4409 22341
rect 4101 22330 4107 22332
rect 4163 22330 4187 22332
rect 4243 22330 4267 22332
rect 4323 22330 4347 22332
rect 4403 22330 4409 22332
rect 4163 22278 4165 22330
rect 4345 22278 4347 22330
rect 4101 22276 4107 22278
rect 4163 22276 4187 22278
rect 4243 22276 4267 22278
rect 4323 22276 4347 22278
rect 4403 22276 4409 22278
rect 4101 22267 4409 22276
rect 5000 22001 5028 22578
rect 4986 21992 5042 22001
rect 4986 21927 5042 21936
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 4101 21244 4409 21253
rect 4101 21242 4107 21244
rect 4163 21242 4187 21244
rect 4243 21242 4267 21244
rect 4323 21242 4347 21244
rect 4403 21242 4409 21244
rect 4163 21190 4165 21242
rect 4345 21190 4347 21242
rect 4101 21188 4107 21190
rect 4163 21188 4187 21190
rect 4243 21188 4267 21190
rect 4323 21188 4347 21190
rect 4403 21188 4409 21190
rect 4101 21179 4409 21188
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 4172 20398 4200 20946
rect 4816 20942 4844 21422
rect 4804 20936 4856 20942
rect 4804 20878 4856 20884
rect 4804 20800 4856 20806
rect 4804 20742 4856 20748
rect 4816 20466 4844 20742
rect 4896 20528 4948 20534
rect 4896 20470 4948 20476
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 3976 20392 4028 20398
rect 3976 20334 4028 20340
rect 4160 20392 4212 20398
rect 4160 20334 4212 20340
rect 4436 20392 4488 20398
rect 4436 20334 4488 20340
rect 3988 19446 4016 20334
rect 4101 20156 4409 20165
rect 4101 20154 4107 20156
rect 4163 20154 4187 20156
rect 4243 20154 4267 20156
rect 4323 20154 4347 20156
rect 4403 20154 4409 20156
rect 4163 20102 4165 20154
rect 4345 20102 4347 20154
rect 4101 20100 4107 20102
rect 4163 20100 4187 20102
rect 4243 20100 4267 20102
rect 4323 20100 4347 20102
rect 4403 20100 4409 20102
rect 4101 20091 4409 20100
rect 4448 20058 4476 20334
rect 4436 20052 4488 20058
rect 4436 19994 4488 20000
rect 4620 19916 4672 19922
rect 4620 19858 4672 19864
rect 4632 19514 4660 19858
rect 4816 19718 4844 20402
rect 4908 20058 4936 20470
rect 4896 20052 4948 20058
rect 4896 19994 4948 20000
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 4620 19508 4672 19514
rect 4620 19450 4672 19456
rect 3976 19440 4028 19446
rect 3976 19382 4028 19388
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 3332 18216 3384 18222
rect 3332 18158 3384 18164
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 1872 16794 1900 17070
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 2228 16516 2280 16522
rect 2228 16458 2280 16464
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 2056 15162 2084 15846
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 2044 12164 2096 12170
rect 2044 12106 2096 12112
rect 2056 11898 2084 12106
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 2240 9654 2268 16458
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 3068 16114 3096 16390
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 3056 16108 3108 16114
rect 3056 16050 3108 16056
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2332 15706 2360 15846
rect 2516 15706 2544 16050
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2608 13938 2636 15506
rect 3252 15502 3280 17138
rect 3344 16658 3372 18158
rect 3528 17678 3556 18226
rect 3988 18222 4016 19382
rect 4632 19334 4660 19450
rect 4632 19306 4752 19334
rect 4101 19068 4409 19077
rect 4101 19066 4107 19068
rect 4163 19066 4187 19068
rect 4243 19066 4267 19068
rect 4323 19066 4347 19068
rect 4403 19066 4409 19068
rect 4163 19014 4165 19066
rect 4345 19014 4347 19066
rect 4101 19012 4107 19014
rect 4163 19012 4187 19014
rect 4243 19012 4267 19014
rect 4323 19012 4347 19014
rect 4403 19012 4409 19014
rect 4101 19003 4409 19012
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 4172 18426 4200 18702
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 4436 18216 4488 18222
rect 4436 18158 4488 18164
rect 4101 17980 4409 17989
rect 4101 17978 4107 17980
rect 4163 17978 4187 17980
rect 4243 17978 4267 17980
rect 4323 17978 4347 17980
rect 4403 17978 4409 17980
rect 4163 17926 4165 17978
rect 4345 17926 4347 17978
rect 4101 17924 4107 17926
rect 4163 17924 4187 17926
rect 4243 17924 4267 17926
rect 4323 17924 4347 17926
rect 4403 17924 4409 17926
rect 4101 17915 4409 17924
rect 3516 17672 3568 17678
rect 3516 17614 3568 17620
rect 3332 16652 3384 16658
rect 3332 16594 3384 16600
rect 3344 16046 3372 16594
rect 3528 16182 3556 17614
rect 4101 16892 4409 16901
rect 4101 16890 4107 16892
rect 4163 16890 4187 16892
rect 4243 16890 4267 16892
rect 4323 16890 4347 16892
rect 4403 16890 4409 16892
rect 4163 16838 4165 16890
rect 4345 16838 4347 16890
rect 4101 16836 4107 16838
rect 4163 16836 4187 16838
rect 4243 16836 4267 16838
rect 4323 16836 4347 16838
rect 4403 16836 4409 16838
rect 4101 16827 4409 16836
rect 3608 16448 3660 16454
rect 3608 16390 3660 16396
rect 3516 16176 3568 16182
rect 3516 16118 3568 16124
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3344 15502 3372 15982
rect 3240 15496 3292 15502
rect 3238 15464 3240 15473
rect 3332 15496 3384 15502
rect 3292 15464 3294 15473
rect 3332 15438 3384 15444
rect 3238 15399 3294 15408
rect 3252 15094 3280 15399
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 3528 15026 3556 16118
rect 3620 15434 3648 16390
rect 4101 15804 4409 15813
rect 4101 15802 4107 15804
rect 4163 15802 4187 15804
rect 4243 15802 4267 15804
rect 4323 15802 4347 15804
rect 4403 15802 4409 15804
rect 4163 15750 4165 15802
rect 4345 15750 4347 15802
rect 4101 15748 4107 15750
rect 4163 15748 4187 15750
rect 4243 15748 4267 15750
rect 4323 15748 4347 15750
rect 4403 15748 4409 15750
rect 4101 15739 4409 15748
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 3608 15428 3660 15434
rect 3608 15370 3660 15376
rect 4080 15162 4108 15438
rect 4172 15162 4200 15642
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 3146 14920 3202 14929
rect 3146 14855 3202 14864
rect 3160 14414 3188 14855
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3712 14618 3740 14758
rect 3700 14612 3752 14618
rect 3700 14554 3752 14560
rect 3988 14482 4016 14962
rect 4356 14890 4384 15302
rect 4344 14884 4396 14890
rect 4344 14826 4396 14832
rect 4101 14716 4409 14725
rect 4101 14714 4107 14716
rect 4163 14714 4187 14716
rect 4243 14714 4267 14716
rect 4323 14714 4347 14716
rect 4403 14714 4409 14716
rect 4163 14662 4165 14714
rect 4345 14662 4347 14714
rect 4101 14660 4107 14662
rect 4163 14660 4187 14662
rect 4243 14660 4267 14662
rect 4323 14660 4347 14662
rect 4403 14660 4409 14662
rect 4101 14651 4409 14660
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3148 14272 3200 14278
rect 3148 14214 3200 14220
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 3160 13870 3188 14214
rect 3344 14006 3372 14214
rect 3332 14000 3384 14006
rect 3332 13942 3384 13948
rect 3148 13864 3200 13870
rect 3148 13806 3200 13812
rect 3160 13326 3188 13806
rect 4101 13628 4409 13637
rect 4101 13626 4107 13628
rect 4163 13626 4187 13628
rect 4243 13626 4267 13628
rect 4323 13626 4347 13628
rect 4403 13626 4409 13628
rect 4163 13574 4165 13626
rect 4345 13574 4347 13626
rect 4101 13572 4107 13574
rect 4163 13572 4187 13574
rect 4243 13572 4267 13574
rect 4323 13572 4347 13574
rect 4403 13572 4409 13574
rect 4101 13563 4409 13572
rect 4344 13456 4396 13462
rect 4448 13410 4476 18158
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 4396 13404 4476 13410
rect 4344 13398 4476 13404
rect 4356 13382 4476 13398
rect 3148 13320 3200 13326
rect 4540 13308 4568 17614
rect 4632 16522 4660 18226
rect 4724 17134 4752 19306
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4816 17066 4844 19654
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 5000 17678 5028 18702
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 4804 17060 4856 17066
rect 4804 17002 4856 17008
rect 5000 16998 5028 17138
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 4724 16522 4752 16662
rect 4620 16516 4672 16522
rect 4620 16458 4672 16464
rect 4712 16516 4764 16522
rect 4712 16458 4764 16464
rect 4632 15366 4660 16458
rect 4724 15706 4752 16458
rect 5000 16182 5028 16934
rect 4988 16176 5040 16182
rect 4988 16118 5040 16124
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 3148 13262 3200 13268
rect 4448 13280 4568 13308
rect 3160 12850 3188 13262
rect 4448 12850 4476 13280
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 3160 12434 3188 12786
rect 4101 12540 4409 12549
rect 4101 12538 4107 12540
rect 4163 12538 4187 12540
rect 4243 12538 4267 12540
rect 4323 12538 4347 12540
rect 4403 12538 4409 12540
rect 4163 12486 4165 12538
rect 4345 12486 4347 12538
rect 4101 12484 4107 12486
rect 4163 12484 4187 12486
rect 4243 12484 4267 12486
rect 4323 12484 4347 12486
rect 4403 12484 4409 12486
rect 4101 12475 4409 12484
rect 2792 12406 3188 12434
rect 2792 12170 2820 12406
rect 4724 12306 4752 15506
rect 5000 15502 5028 16118
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 4816 13870 4844 14826
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4908 13938 4936 14758
rect 5092 13938 5120 26930
rect 7196 26784 7248 26790
rect 7196 26726 7248 26732
rect 9772 26784 9824 26790
rect 9772 26726 9824 26732
rect 10784 26784 10836 26790
rect 10784 26726 10836 26732
rect 7208 26586 7236 26726
rect 7196 26580 7248 26586
rect 7196 26522 7248 26528
rect 8484 26376 8536 26382
rect 8484 26318 8536 26324
rect 7656 26308 7708 26314
rect 7656 26250 7708 26256
rect 7252 26140 7560 26149
rect 7252 26138 7258 26140
rect 7314 26138 7338 26140
rect 7394 26138 7418 26140
rect 7474 26138 7498 26140
rect 7554 26138 7560 26140
rect 7314 26086 7316 26138
rect 7496 26086 7498 26138
rect 7252 26084 7258 26086
rect 7314 26084 7338 26086
rect 7394 26084 7418 26086
rect 7474 26084 7498 26086
rect 7554 26084 7560 26086
rect 7252 26075 7560 26084
rect 7472 25968 7524 25974
rect 7668 25956 7696 26250
rect 8024 26240 8076 26246
rect 8024 26182 8076 26188
rect 8208 26240 8260 26246
rect 8208 26182 8260 26188
rect 8036 25974 8064 26182
rect 7524 25928 7696 25956
rect 7472 25910 7524 25916
rect 5908 25832 5960 25838
rect 6920 25832 6972 25838
rect 5908 25774 5960 25780
rect 6840 25792 6920 25820
rect 5356 25696 5408 25702
rect 5356 25638 5408 25644
rect 5368 25362 5396 25638
rect 5356 25356 5408 25362
rect 5356 25298 5408 25304
rect 5920 24698 5948 25774
rect 6276 25220 6328 25226
rect 6276 25162 6328 25168
rect 6288 24886 6316 25162
rect 6000 24880 6052 24886
rect 6000 24822 6052 24828
rect 6276 24880 6328 24886
rect 6276 24822 6328 24828
rect 5828 24670 5948 24698
rect 5828 24206 5856 24670
rect 5448 24200 5500 24206
rect 5448 24142 5500 24148
rect 5816 24200 5868 24206
rect 5816 24142 5868 24148
rect 5356 23724 5408 23730
rect 5356 23666 5408 23672
rect 5368 22778 5396 23666
rect 5460 23662 5488 24142
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 5356 22772 5408 22778
rect 5356 22714 5408 22720
rect 5368 22094 5396 22714
rect 5460 22710 5488 23054
rect 5448 22704 5500 22710
rect 5448 22646 5500 22652
rect 5828 22642 5856 24142
rect 6012 23118 6040 24822
rect 6460 24812 6512 24818
rect 6460 24754 6512 24760
rect 6472 24721 6500 24754
rect 6458 24712 6514 24721
rect 6458 24647 6514 24656
rect 6840 24070 6868 25792
rect 6920 25774 6972 25780
rect 7484 25702 7512 25910
rect 7472 25696 7524 25702
rect 7472 25638 7524 25644
rect 6920 25220 6972 25226
rect 6920 25162 6972 25168
rect 6932 24818 6960 25162
rect 7104 25152 7156 25158
rect 7104 25094 7156 25100
rect 7116 24818 7144 25094
rect 7252 25052 7560 25061
rect 7252 25050 7258 25052
rect 7314 25050 7338 25052
rect 7394 25050 7418 25052
rect 7474 25050 7498 25052
rect 7554 25050 7560 25052
rect 7314 24998 7316 25050
rect 7496 24998 7498 25050
rect 7252 24996 7258 24998
rect 7314 24996 7338 24998
rect 7394 24996 7418 24998
rect 7474 24996 7498 24998
rect 7554 24996 7560 24998
rect 7252 24987 7560 24996
rect 7668 24886 7696 25928
rect 8024 25968 8076 25974
rect 8024 25910 8076 25916
rect 8220 25362 8248 26182
rect 8496 25838 8524 26318
rect 8852 26308 8904 26314
rect 8852 26250 8904 26256
rect 8484 25832 8536 25838
rect 8484 25774 8536 25780
rect 8760 25832 8812 25838
rect 8760 25774 8812 25780
rect 8208 25356 8260 25362
rect 8208 25298 8260 25304
rect 7656 24880 7708 24886
rect 7656 24822 7708 24828
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 7104 24812 7156 24818
rect 7104 24754 7156 24760
rect 7196 24812 7248 24818
rect 7196 24754 7248 24760
rect 7208 24410 7236 24754
rect 7562 24712 7618 24721
rect 7562 24647 7564 24656
rect 7616 24647 7618 24656
rect 7564 24618 7616 24624
rect 7196 24404 7248 24410
rect 7196 24346 7248 24352
rect 6460 24064 6512 24070
rect 6460 24006 6512 24012
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 7104 24064 7156 24070
rect 7104 24006 7156 24012
rect 6472 23730 6500 24006
rect 6460 23724 6512 23730
rect 6460 23666 6512 23672
rect 6276 23520 6328 23526
rect 6276 23462 6328 23468
rect 6000 23112 6052 23118
rect 6000 23054 6052 23060
rect 6288 23050 6316 23462
rect 6472 23322 6500 23666
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 6460 23316 6512 23322
rect 6460 23258 6512 23264
rect 6932 23254 6960 23598
rect 6920 23248 6972 23254
rect 6920 23190 6972 23196
rect 6920 23112 6972 23118
rect 6920 23054 6972 23060
rect 7116 23066 7144 24006
rect 7252 23964 7560 23973
rect 7252 23962 7258 23964
rect 7314 23962 7338 23964
rect 7394 23962 7418 23964
rect 7474 23962 7498 23964
rect 7554 23962 7560 23964
rect 7314 23910 7316 23962
rect 7496 23910 7498 23962
rect 7252 23908 7258 23910
rect 7314 23908 7338 23910
rect 7394 23908 7418 23910
rect 7474 23908 7498 23910
rect 7554 23908 7560 23910
rect 7252 23899 7560 23908
rect 7668 23866 7696 24822
rect 8496 24818 8524 25774
rect 8772 25498 8800 25774
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 8864 25294 8892 26250
rect 9588 25356 9640 25362
rect 9588 25298 9640 25304
rect 8576 25288 8628 25294
rect 8576 25230 8628 25236
rect 8852 25288 8904 25294
rect 8852 25230 8904 25236
rect 8588 24954 8616 25230
rect 9496 25152 9548 25158
rect 9496 25094 9548 25100
rect 8576 24948 8628 24954
rect 8576 24890 8628 24896
rect 8484 24812 8536 24818
rect 8484 24754 8536 24760
rect 9508 24750 9536 25094
rect 9404 24744 9456 24750
rect 9404 24686 9456 24692
rect 9496 24744 9548 24750
rect 9496 24686 9548 24692
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 8312 23866 8340 24210
rect 7656 23860 7708 23866
rect 7656 23802 7708 23808
rect 8300 23860 8352 23866
rect 8300 23802 8352 23808
rect 6276 23044 6328 23050
rect 6276 22986 6328 22992
rect 6552 23044 6604 23050
rect 6552 22986 6604 22992
rect 6184 22704 6236 22710
rect 6184 22646 6236 22652
rect 5816 22636 5868 22642
rect 5816 22578 5868 22584
rect 5908 22432 5960 22438
rect 5908 22374 5960 22380
rect 5276 22066 5396 22094
rect 5276 21010 5304 22066
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5552 21690 5580 21966
rect 5816 21956 5868 21962
rect 5816 21898 5868 21904
rect 5540 21684 5592 21690
rect 5540 21626 5592 21632
rect 5828 21146 5856 21898
rect 5816 21140 5868 21146
rect 5816 21082 5868 21088
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 5264 20868 5316 20874
rect 5264 20810 5316 20816
rect 5276 19854 5304 20810
rect 5356 20596 5408 20602
rect 5356 20538 5408 20544
rect 5368 19854 5396 20538
rect 5448 20460 5500 20466
rect 5448 20402 5500 20408
rect 5644 20420 5856 20448
rect 5460 20058 5488 20402
rect 5644 20330 5672 20420
rect 5828 20330 5856 20420
rect 5632 20324 5684 20330
rect 5632 20266 5684 20272
rect 5724 20324 5776 20330
rect 5724 20266 5776 20272
rect 5816 20324 5868 20330
rect 5816 20266 5868 20272
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 5644 19854 5672 20266
rect 5736 19854 5764 20266
rect 5264 19848 5316 19854
rect 5262 19816 5264 19825
rect 5356 19848 5408 19854
rect 5316 19816 5318 19825
rect 5356 19790 5408 19796
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5262 19751 5318 19760
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 5184 19378 5212 19654
rect 5368 19514 5396 19790
rect 5816 19780 5868 19786
rect 5816 19722 5868 19728
rect 5828 19514 5856 19722
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5816 19508 5868 19514
rect 5816 19450 5868 19456
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5184 18970 5212 19314
rect 5644 18970 5672 19314
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 5632 18964 5684 18970
rect 5632 18906 5684 18912
rect 5632 18760 5684 18766
rect 5816 18760 5868 18766
rect 5684 18720 5816 18748
rect 5632 18702 5684 18708
rect 5816 18702 5868 18708
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5264 17672 5316 17678
rect 5264 17614 5316 17620
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5172 17536 5224 17542
rect 5172 17478 5224 17484
rect 5184 17202 5212 17478
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 5184 16590 5212 17138
rect 5276 16794 5304 17614
rect 5368 17338 5396 17614
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5552 17202 5580 18022
rect 5644 17746 5672 18702
rect 5920 18290 5948 22374
rect 6000 21344 6052 21350
rect 6000 21286 6052 21292
rect 6012 20466 6040 21286
rect 6196 20942 6224 22646
rect 6288 22438 6316 22986
rect 6276 22432 6328 22438
rect 6276 22374 6328 22380
rect 6276 21548 6328 21554
rect 6276 21490 6328 21496
rect 6184 20936 6236 20942
rect 6104 20896 6184 20924
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 6012 20058 6040 20402
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 6104 19514 6132 20896
rect 6184 20878 6236 20884
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 6196 20466 6224 20742
rect 6184 20460 6236 20466
rect 6184 20402 6236 20408
rect 6184 20052 6236 20058
rect 6184 19994 6236 20000
rect 6196 19922 6224 19994
rect 6288 19922 6316 21490
rect 6368 21480 6420 21486
rect 6368 21422 6420 21428
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 6276 19916 6328 19922
rect 6276 19858 6328 19864
rect 6182 19816 6238 19825
rect 6182 19751 6238 19760
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 6012 18834 6040 19110
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5632 17740 5684 17746
rect 5632 17682 5684 17688
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 5184 16114 5212 16526
rect 5276 16114 5304 16730
rect 5368 16658 5396 17138
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5368 15978 5396 16594
rect 5460 16402 5488 17138
rect 5552 16590 5580 17138
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5632 16448 5684 16454
rect 5460 16374 5580 16402
rect 5632 16390 5684 16396
rect 5356 15972 5408 15978
rect 5356 15914 5408 15920
rect 5552 15042 5580 16374
rect 5644 16250 5672 16390
rect 5632 16244 5684 16250
rect 5632 16186 5684 16192
rect 5736 16114 5764 17614
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5736 15162 5764 16050
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5552 15014 5764 15042
rect 4896 13932 4948 13938
rect 5080 13932 5132 13938
rect 4896 13874 4948 13880
rect 5000 13892 5080 13920
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4908 13258 4936 13874
rect 5000 13530 5028 13892
rect 5080 13874 5132 13880
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5644 13530 5672 13670
rect 5736 13530 5764 15014
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 4896 13252 4948 13258
rect 4896 13194 4948 13200
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5460 12782 5488 13126
rect 5736 12918 5764 13262
rect 5724 12912 5776 12918
rect 5724 12854 5776 12860
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2792 11762 2820 12106
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3620 11898 3648 12038
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2792 10742 2820 11698
rect 3712 11354 3740 12242
rect 3976 12164 4028 12170
rect 3976 12106 4028 12112
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3160 10810 3188 11086
rect 3608 11008 3660 11014
rect 3608 10950 3660 10956
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 3160 10690 3188 10746
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 1768 9444 1820 9450
rect 1768 9386 1820 9392
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 2148 8362 2176 9318
rect 2424 9042 2452 9862
rect 2596 9648 2648 9654
rect 2596 9590 2648 9596
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 2608 8514 2636 9590
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2700 8634 2728 9114
rect 2792 8974 2820 10678
rect 3160 10662 3280 10690
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2884 9586 2912 10066
rect 3068 10062 3096 10406
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2884 9042 2912 9522
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1964 6458 1992 6598
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 940 4548 992 4554
rect 940 4490 992 4496
rect 952 4185 980 4490
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 1412 3602 1440 6258
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 2240 2446 2268 8298
rect 2332 8276 2360 8502
rect 2608 8498 2728 8514
rect 2608 8492 2740 8498
rect 2608 8486 2688 8492
rect 2688 8434 2740 8440
rect 2504 8288 2556 8294
rect 2332 8248 2504 8276
rect 2504 8230 2556 8236
rect 2792 6322 2820 8910
rect 2884 8498 2912 8978
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2884 8090 2912 8230
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2976 7886 3004 9318
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 3068 6866 3096 9998
rect 3252 9994 3280 10662
rect 3620 10606 3648 10950
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3712 10470 3740 11290
rect 3792 11280 3844 11286
rect 3792 11222 3844 11228
rect 3804 10674 3832 11222
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3240 9988 3292 9994
rect 3240 9930 3292 9936
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3160 8362 3188 9454
rect 3252 9382 3280 9930
rect 3896 9654 3924 11494
rect 3988 10062 4016 12106
rect 4908 11830 4936 12718
rect 5644 12594 5672 12786
rect 5828 12646 5856 17070
rect 5920 16726 5948 18226
rect 6104 17882 6132 19450
rect 6196 19378 6224 19751
rect 6380 19378 6408 21422
rect 6564 21146 6592 22986
rect 6828 22976 6880 22982
rect 6828 22918 6880 22924
rect 6840 22642 6868 22918
rect 6828 22636 6880 22642
rect 6932 22624 6960 23054
rect 7116 23050 7236 23066
rect 7116 23044 7248 23050
rect 7116 23038 7196 23044
rect 7196 22986 7248 22992
rect 7668 22982 7696 23802
rect 9036 23724 9088 23730
rect 9036 23666 9088 23672
rect 9312 23724 9364 23730
rect 9312 23666 9364 23672
rect 8484 23520 8536 23526
rect 8484 23462 8536 23468
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 7104 22976 7156 22982
rect 7104 22918 7156 22924
rect 7656 22976 7708 22982
rect 7656 22918 7708 22924
rect 7116 22778 7144 22918
rect 7252 22876 7560 22885
rect 7252 22874 7258 22876
rect 7314 22874 7338 22876
rect 7394 22874 7418 22876
rect 7474 22874 7498 22876
rect 7554 22874 7560 22876
rect 7314 22822 7316 22874
rect 7496 22822 7498 22874
rect 7252 22820 7258 22822
rect 7314 22820 7338 22822
rect 7394 22820 7418 22822
rect 7474 22820 7498 22822
rect 7554 22820 7560 22822
rect 7252 22811 7560 22820
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 7104 22636 7156 22642
rect 6932 22596 7104 22624
rect 6828 22578 6880 22584
rect 7104 22578 7156 22584
rect 6840 22098 6868 22578
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 6828 22092 6880 22098
rect 6656 22052 6828 22080
rect 6552 21140 6604 21146
rect 6552 21082 6604 21088
rect 6656 21010 6684 22052
rect 6828 22034 6880 22040
rect 6932 22030 6960 22170
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 6932 21298 6960 21966
rect 6932 21270 7052 21298
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6644 21004 6696 21010
rect 6472 20964 6644 20992
rect 6472 19904 6500 20964
rect 6644 20946 6696 20952
rect 6552 20800 6604 20806
rect 6748 20754 6776 21082
rect 6918 20904 6974 20913
rect 6918 20839 6974 20848
rect 6604 20748 6776 20754
rect 6552 20742 6776 20748
rect 6564 20726 6776 20742
rect 6748 20602 6776 20726
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 6736 20596 6788 20602
rect 6736 20538 6788 20544
rect 6656 20466 6684 20538
rect 6644 20460 6696 20466
rect 6644 20402 6696 20408
rect 6932 20058 6960 20839
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6552 19916 6604 19922
rect 6472 19876 6552 19904
rect 6552 19858 6604 19864
rect 6460 19780 6512 19786
rect 6460 19722 6512 19728
rect 6472 19514 6500 19722
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6184 19372 6236 19378
rect 6368 19372 6420 19378
rect 6236 19320 6316 19334
rect 6184 19314 6316 19320
rect 6368 19314 6420 19320
rect 6196 19306 6316 19314
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6196 18222 6224 18566
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6092 17876 6144 17882
rect 6092 17818 6144 17824
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 6012 16674 6040 17614
rect 6196 16998 6224 18158
rect 6288 17678 6316 19306
rect 6380 18290 6408 19314
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6380 17814 6408 18226
rect 6460 18216 6512 18222
rect 6460 18158 6512 18164
rect 6472 17882 6500 18158
rect 6460 17876 6512 17882
rect 6460 17818 6512 17824
rect 6564 17814 6592 19858
rect 7024 19786 7052 21270
rect 7116 21128 7144 22578
rect 7668 22234 7696 22918
rect 8312 22778 8340 23122
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8496 22574 8524 23462
rect 9048 23322 9076 23666
rect 9128 23520 9180 23526
rect 9128 23462 9180 23468
rect 9036 23316 9088 23322
rect 9036 23258 9088 23264
rect 9140 22778 9168 23462
rect 9128 22772 9180 22778
rect 9128 22714 9180 22720
rect 8484 22568 8536 22574
rect 8484 22510 8536 22516
rect 7656 22228 7708 22234
rect 7656 22170 7708 22176
rect 8024 21888 8076 21894
rect 8024 21830 8076 21836
rect 8576 21888 8628 21894
rect 8576 21830 8628 21836
rect 7252 21788 7560 21797
rect 7252 21786 7258 21788
rect 7314 21786 7338 21788
rect 7394 21786 7418 21788
rect 7474 21786 7498 21788
rect 7554 21786 7560 21788
rect 7314 21734 7316 21786
rect 7496 21734 7498 21786
rect 7252 21732 7258 21734
rect 7314 21732 7338 21734
rect 7394 21732 7418 21734
rect 7474 21732 7498 21734
rect 7554 21732 7560 21734
rect 7252 21723 7560 21732
rect 8036 21486 8064 21830
rect 8588 21622 8616 21830
rect 8576 21616 8628 21622
rect 8576 21558 8628 21564
rect 8300 21548 8352 21554
rect 8300 21490 8352 21496
rect 7472 21480 7524 21486
rect 7472 21422 7524 21428
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 7116 21100 7236 21128
rect 7104 20936 7156 20942
rect 7208 20913 7236 21100
rect 7104 20878 7156 20884
rect 7194 20904 7250 20913
rect 7116 20602 7144 20878
rect 7300 20874 7328 21286
rect 7392 21010 7420 21286
rect 7380 21004 7432 21010
rect 7380 20946 7432 20952
rect 7484 20874 7512 21422
rect 7194 20839 7196 20848
rect 7248 20839 7250 20848
rect 7288 20868 7340 20874
rect 7196 20810 7248 20816
rect 7288 20810 7340 20816
rect 7472 20868 7524 20874
rect 7472 20810 7524 20816
rect 8116 20868 8168 20874
rect 8116 20810 8168 20816
rect 7252 20700 7560 20709
rect 7252 20698 7258 20700
rect 7314 20698 7338 20700
rect 7394 20698 7418 20700
rect 7474 20698 7498 20700
rect 7554 20698 7560 20700
rect 7314 20646 7316 20698
rect 7496 20646 7498 20698
rect 7252 20644 7258 20646
rect 7314 20644 7338 20646
rect 7394 20644 7418 20646
rect 7474 20644 7498 20646
rect 7554 20644 7560 20646
rect 7252 20635 7560 20644
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 7012 19780 7064 19786
rect 7012 19722 7064 19728
rect 7252 19612 7560 19621
rect 7252 19610 7258 19612
rect 7314 19610 7338 19612
rect 7394 19610 7418 19612
rect 7474 19610 7498 19612
rect 7554 19610 7560 19612
rect 7314 19558 7316 19610
rect 7496 19558 7498 19610
rect 7252 19556 7258 19558
rect 7314 19556 7338 19558
rect 7394 19556 7418 19558
rect 7474 19556 7498 19558
rect 7554 19556 7560 19558
rect 7252 19547 7560 19556
rect 8036 19378 8064 19994
rect 8128 19854 8156 20810
rect 8312 19922 8340 21490
rect 9324 21146 9352 23666
rect 9312 21140 9364 21146
rect 9312 21082 9364 21088
rect 9416 21010 9444 24686
rect 9508 24342 9536 24686
rect 9496 24336 9548 24342
rect 9496 24278 9548 24284
rect 9600 22386 9628 25298
rect 9784 24954 9812 26726
rect 10403 26684 10711 26693
rect 10403 26682 10409 26684
rect 10465 26682 10489 26684
rect 10545 26682 10569 26684
rect 10625 26682 10649 26684
rect 10705 26682 10711 26684
rect 10465 26630 10467 26682
rect 10647 26630 10649 26682
rect 10403 26628 10409 26630
rect 10465 26628 10489 26630
rect 10545 26628 10569 26630
rect 10625 26628 10649 26630
rect 10705 26628 10711 26630
rect 10403 26619 10711 26628
rect 10796 26586 10824 26726
rect 10784 26580 10836 26586
rect 10784 26522 10836 26528
rect 10980 26489 11008 26930
rect 10966 26480 11022 26489
rect 10966 26415 11022 26424
rect 11348 26382 11376 26930
rect 11428 26784 11480 26790
rect 11428 26726 11480 26732
rect 12256 26784 12308 26790
rect 12256 26726 12308 26732
rect 12440 26784 12492 26790
rect 12440 26726 12492 26732
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 9956 26240 10008 26246
rect 9956 26182 10008 26188
rect 9968 25362 9996 26182
rect 11348 26042 11376 26318
rect 11336 26036 11388 26042
rect 11336 25978 11388 25984
rect 11336 25900 11388 25906
rect 11336 25842 11388 25848
rect 10876 25832 10928 25838
rect 10876 25774 10928 25780
rect 10784 25696 10836 25702
rect 10784 25638 10836 25644
rect 10403 25596 10711 25605
rect 10403 25594 10409 25596
rect 10465 25594 10489 25596
rect 10545 25594 10569 25596
rect 10625 25594 10649 25596
rect 10705 25594 10711 25596
rect 10465 25542 10467 25594
rect 10647 25542 10649 25594
rect 10403 25540 10409 25542
rect 10465 25540 10489 25542
rect 10545 25540 10569 25542
rect 10625 25540 10649 25542
rect 10705 25540 10711 25542
rect 10403 25531 10711 25540
rect 10796 25498 10824 25638
rect 10784 25492 10836 25498
rect 10784 25434 10836 25440
rect 9956 25356 10008 25362
rect 9956 25298 10008 25304
rect 10888 25226 10916 25774
rect 10876 25220 10928 25226
rect 10876 25162 10928 25168
rect 9772 24948 9824 24954
rect 9772 24890 9824 24896
rect 10888 24818 10916 25162
rect 11348 24954 11376 25842
rect 11336 24948 11388 24954
rect 11336 24890 11388 24896
rect 10876 24812 10928 24818
rect 10876 24754 10928 24760
rect 9864 24744 9916 24750
rect 9864 24686 9916 24692
rect 9876 24410 9904 24686
rect 10403 24508 10711 24517
rect 10403 24506 10409 24508
rect 10465 24506 10489 24508
rect 10545 24506 10569 24508
rect 10625 24506 10649 24508
rect 10705 24506 10711 24508
rect 10465 24454 10467 24506
rect 10647 24454 10649 24506
rect 10403 24452 10409 24454
rect 10465 24452 10489 24454
rect 10545 24452 10569 24454
rect 10625 24452 10649 24454
rect 10705 24452 10711 24454
rect 10403 24443 10711 24452
rect 9864 24404 9916 24410
rect 9864 24346 9916 24352
rect 10324 23520 10376 23526
rect 10324 23462 10376 23468
rect 10336 23322 10364 23462
rect 10403 23420 10711 23429
rect 10403 23418 10409 23420
rect 10465 23418 10489 23420
rect 10545 23418 10569 23420
rect 10625 23418 10649 23420
rect 10705 23418 10711 23420
rect 10465 23366 10467 23418
rect 10647 23366 10649 23418
rect 10403 23364 10409 23366
rect 10465 23364 10489 23366
rect 10545 23364 10569 23366
rect 10625 23364 10649 23366
rect 10705 23364 10711 23366
rect 10403 23355 10711 23364
rect 10324 23316 10376 23322
rect 10324 23258 10376 23264
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 10140 23044 10192 23050
rect 10140 22986 10192 22992
rect 9864 22704 9916 22710
rect 9864 22646 9916 22652
rect 9772 22568 9824 22574
rect 9772 22510 9824 22516
rect 9600 22358 9720 22386
rect 9600 22234 9628 22358
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 9588 21888 9640 21894
rect 9588 21830 9640 21836
rect 9600 21554 9628 21830
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 9220 20256 9272 20262
rect 9220 20198 9272 20204
rect 9232 19922 9260 20198
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 9220 19916 9272 19922
rect 9220 19858 9272 19864
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 6918 19272 6974 19281
rect 6918 19207 6974 19216
rect 6932 18426 6960 19207
rect 7252 18524 7560 18533
rect 7252 18522 7258 18524
rect 7314 18522 7338 18524
rect 7394 18522 7418 18524
rect 7474 18522 7498 18524
rect 7554 18522 7560 18524
rect 7314 18470 7316 18522
rect 7496 18470 7498 18522
rect 7252 18468 7258 18470
rect 7314 18468 7338 18470
rect 7394 18468 7418 18470
rect 7474 18468 7498 18470
rect 7554 18468 7560 18470
rect 7252 18459 7560 18468
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 6828 18284 6880 18290
rect 6828 18226 6880 18232
rect 6368 17808 6420 17814
rect 6368 17750 6420 17756
rect 6552 17808 6604 17814
rect 6552 17750 6604 17756
rect 6736 17808 6788 17814
rect 6736 17750 6788 17756
rect 6276 17672 6328 17678
rect 6276 17614 6328 17620
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6380 17338 6408 17614
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6564 17270 6592 17614
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6552 17264 6604 17270
rect 6552 17206 6604 17212
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6288 17066 6316 17138
rect 6276 17060 6328 17066
rect 6276 17002 6328 17008
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 6104 16794 6132 16934
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 6012 16646 6132 16674
rect 5906 15464 5962 15473
rect 5906 15399 5908 15408
rect 5960 15399 5962 15408
rect 5908 15370 5960 15376
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 5552 12566 5672 12594
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5552 12238 5580 12566
rect 5736 12434 5764 12582
rect 5736 12406 5856 12434
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 11830 5580 12174
rect 4896 11824 4948 11830
rect 4896 11766 4948 11772
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 4101 11452 4409 11461
rect 4101 11450 4107 11452
rect 4163 11450 4187 11452
rect 4243 11450 4267 11452
rect 4323 11450 4347 11452
rect 4403 11450 4409 11452
rect 4163 11398 4165 11450
rect 4345 11398 4347 11450
rect 4101 11396 4107 11398
rect 4163 11396 4187 11398
rect 4243 11396 4267 11398
rect 4323 11396 4347 11398
rect 4403 11396 4409 11398
rect 4101 11387 4409 11396
rect 4908 11286 4936 11766
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 11354 5580 11494
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 4896 11280 4948 11286
rect 4896 11222 4948 11228
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4724 10674 4752 11154
rect 5630 10704 5686 10713
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 5552 10662 5630 10690
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 4101 10364 4409 10373
rect 4101 10362 4107 10364
rect 4163 10362 4187 10364
rect 4243 10362 4267 10364
rect 4323 10362 4347 10364
rect 4403 10362 4409 10364
rect 4163 10310 4165 10362
rect 4345 10310 4347 10362
rect 4101 10308 4107 10310
rect 4163 10308 4187 10310
rect 4243 10308 4267 10310
rect 4323 10308 4347 10310
rect 4403 10308 4409 10310
rect 4101 10299 4409 10308
rect 5460 10266 5488 10406
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5552 10130 5580 10662
rect 5630 10639 5686 10648
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5644 10266 5672 10542
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 3988 9722 4016 9998
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 4080 9674 4108 9998
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 3884 9648 3936 9654
rect 3882 9616 3884 9625
rect 3936 9616 3938 9625
rect 3988 9586 4016 9658
rect 4080 9646 4200 9674
rect 4172 9586 4200 9646
rect 4344 9614 4396 9620
rect 3882 9551 3938 9560
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 4160 9580 4212 9586
rect 4528 9580 4580 9586
rect 4396 9562 4476 9568
rect 4344 9556 4476 9562
rect 4356 9540 4476 9556
rect 4160 9522 4212 9528
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 9178 3280 9318
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3344 8634 3372 9454
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 3160 8090 3188 8298
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3344 7886 3372 8570
rect 3712 8430 3740 9318
rect 3884 9172 3936 9178
rect 3988 9160 4016 9318
rect 4101 9276 4409 9285
rect 4101 9274 4107 9276
rect 4163 9274 4187 9276
rect 4243 9274 4267 9276
rect 4323 9274 4347 9276
rect 4403 9274 4409 9276
rect 4163 9222 4165 9274
rect 4345 9222 4347 9274
rect 4101 9220 4107 9222
rect 4163 9220 4187 9222
rect 4243 9220 4267 9222
rect 4323 9220 4347 9222
rect 4403 9220 4409 9222
rect 4101 9211 4409 9220
rect 4448 9178 4476 9540
rect 4528 9522 4580 9528
rect 4540 9382 4568 9522
rect 4632 9382 4660 9930
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4436 9172 4488 9178
rect 3988 9132 4108 9160
rect 3884 9114 3936 9120
rect 3896 8974 3924 9114
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 4080 8906 4108 9132
rect 4436 9114 4488 9120
rect 4252 9104 4304 9110
rect 4252 9046 4304 9052
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3804 8498 3832 8774
rect 4080 8634 4108 8842
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4172 8498 4200 8910
rect 4264 8634 4292 9046
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 3160 6118 3188 6734
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3160 4622 3188 6054
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3436 3398 3464 6258
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3528 2514 3556 8366
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3712 7886 3740 8230
rect 3804 8090 3832 8434
rect 4080 8294 4108 8434
rect 4540 8294 4568 9318
rect 4632 8974 4660 9318
rect 4724 8974 4752 9658
rect 4802 9616 4858 9625
rect 4802 9551 4804 9560
rect 4856 9551 4858 9560
rect 4804 9522 4856 9528
rect 4816 8974 4844 9522
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4724 8498 4752 8910
rect 4908 8498 4936 8978
rect 5276 8974 5304 9046
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4896 8356 4948 8362
rect 4896 8298 4948 8304
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4101 8188 4409 8197
rect 4101 8186 4107 8188
rect 4163 8186 4187 8188
rect 4243 8186 4267 8188
rect 4323 8186 4347 8188
rect 4403 8186 4409 8188
rect 4163 8134 4165 8186
rect 4345 8134 4347 8186
rect 4101 8132 4107 8134
rect 4163 8132 4187 8134
rect 4243 8132 4267 8134
rect 4323 8132 4347 8134
rect 4403 8132 4409 8134
rect 4101 8123 4409 8132
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3988 5166 4016 7686
rect 4101 7100 4409 7109
rect 4101 7098 4107 7100
rect 4163 7098 4187 7100
rect 4243 7098 4267 7100
rect 4323 7098 4347 7100
rect 4403 7098 4409 7100
rect 4163 7046 4165 7098
rect 4345 7046 4347 7098
rect 4101 7044 4107 7046
rect 4163 7044 4187 7046
rect 4243 7044 4267 7046
rect 4323 7044 4347 7046
rect 4403 7044 4409 7046
rect 4101 7035 4409 7044
rect 4101 6012 4409 6021
rect 4101 6010 4107 6012
rect 4163 6010 4187 6012
rect 4243 6010 4267 6012
rect 4323 6010 4347 6012
rect 4403 6010 4409 6012
rect 4163 5958 4165 6010
rect 4345 5958 4347 6010
rect 4101 5956 4107 5958
rect 4163 5956 4187 5958
rect 4243 5956 4267 5958
rect 4323 5956 4347 5958
rect 4403 5956 4409 5958
rect 4101 5947 4409 5956
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 4101 4924 4409 4933
rect 4101 4922 4107 4924
rect 4163 4922 4187 4924
rect 4243 4922 4267 4924
rect 4323 4922 4347 4924
rect 4403 4922 4409 4924
rect 4163 4870 4165 4922
rect 4345 4870 4347 4922
rect 4101 4868 4107 4870
rect 4163 4868 4187 4870
rect 4243 4868 4267 4870
rect 4323 4868 4347 4870
rect 4403 4868 4409 4870
rect 4101 4859 4409 4868
rect 4101 3836 4409 3845
rect 4101 3834 4107 3836
rect 4163 3834 4187 3836
rect 4243 3834 4267 3836
rect 4323 3834 4347 3836
rect 4403 3834 4409 3836
rect 4163 3782 4165 3834
rect 4345 3782 4347 3834
rect 4101 3780 4107 3782
rect 4163 3780 4187 3782
rect 4243 3780 4267 3782
rect 4323 3780 4347 3782
rect 4403 3780 4409 3782
rect 4101 3771 4409 3780
rect 4101 2748 4409 2757
rect 4101 2746 4107 2748
rect 4163 2746 4187 2748
rect 4243 2746 4267 2748
rect 4323 2746 4347 2748
rect 4403 2746 4409 2748
rect 4163 2694 4165 2746
rect 4345 2694 4347 2746
rect 4101 2692 4107 2694
rect 4163 2692 4187 2694
rect 4243 2692 4267 2694
rect 4323 2692 4347 2694
rect 4403 2692 4409 2694
rect 4101 2683 4409 2692
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 4908 2446 4936 8298
rect 5552 8090 5580 9862
rect 5644 9382 5672 9998
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5644 8430 5672 9318
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5736 6730 5764 12310
rect 5828 11762 5856 12406
rect 5920 12238 5948 14350
rect 6000 13796 6052 13802
rect 6000 13738 6052 13744
rect 6012 13326 6040 13738
rect 6104 13530 6132 16646
rect 6196 15026 6224 16934
rect 6288 16454 6316 17002
rect 6380 16590 6408 17138
rect 6656 17134 6684 17478
rect 6644 17128 6696 17134
rect 6644 17070 6696 17076
rect 6460 16992 6512 16998
rect 6460 16934 6512 16940
rect 6472 16658 6500 16934
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 6748 16590 6776 17750
rect 6840 17066 6868 18226
rect 8024 18216 8076 18222
rect 8024 18158 8076 18164
rect 8036 17882 8064 18158
rect 8024 17876 8076 17882
rect 8024 17818 8076 17824
rect 8128 17746 8156 19790
rect 8312 19394 8340 19858
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8588 19446 8616 19654
rect 8220 19378 8340 19394
rect 8576 19440 8628 19446
rect 8576 19382 8628 19388
rect 8220 19372 8352 19378
rect 8220 19366 8300 19372
rect 8220 18426 8248 19366
rect 8300 19314 8352 19320
rect 8772 18970 8800 19790
rect 9416 19310 9444 20946
rect 9692 20398 9720 22358
rect 9784 21962 9812 22510
rect 9772 21956 9824 21962
rect 9772 21898 9824 21904
rect 9876 21554 9904 22646
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9968 22012 9996 22374
rect 10048 22024 10100 22030
rect 9968 21984 10048 22012
rect 10048 21966 10100 21972
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 9680 20392 9732 20398
rect 9732 20352 9812 20380
rect 9680 20334 9732 20340
rect 9680 19440 9732 19446
rect 9680 19382 9732 19388
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 9416 18834 9444 19246
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 6828 17060 6880 17066
rect 6828 17002 6880 17008
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6276 16108 6328 16114
rect 6276 16050 6328 16056
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6196 13462 6224 13874
rect 6184 13456 6236 13462
rect 6184 13398 6236 13404
rect 6288 13326 6316 16050
rect 6380 15366 6408 16390
rect 6564 16250 6592 16526
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6748 16114 6776 16526
rect 6920 16516 6972 16522
rect 6920 16458 6972 16464
rect 6932 16250 6960 16458
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 6828 15972 6880 15978
rect 6828 15914 6880 15920
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6472 14618 6500 15098
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6564 14482 6592 14962
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6748 14482 6776 14894
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6840 13530 6868 15914
rect 6932 15706 6960 16050
rect 7024 16046 7052 17138
rect 7116 17134 7144 17614
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7252 17436 7560 17445
rect 7252 17434 7258 17436
rect 7314 17434 7338 17436
rect 7394 17434 7418 17436
rect 7474 17434 7498 17436
rect 7554 17434 7560 17436
rect 7314 17382 7316 17434
rect 7496 17382 7498 17434
rect 7252 17380 7258 17382
rect 7314 17380 7338 17382
rect 7394 17380 7418 17382
rect 7474 17380 7498 17382
rect 7554 17380 7560 17382
rect 7252 17371 7560 17380
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7116 16046 7144 17070
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7252 16348 7560 16357
rect 7252 16346 7258 16348
rect 7314 16346 7338 16348
rect 7394 16346 7418 16348
rect 7474 16346 7498 16348
rect 7554 16346 7560 16348
rect 7314 16294 7316 16346
rect 7496 16294 7498 16346
rect 7252 16292 7258 16294
rect 7314 16292 7338 16294
rect 7394 16292 7418 16294
rect 7474 16292 7498 16294
rect 7554 16292 7560 16294
rect 7252 16283 7560 16292
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7024 15706 7052 15982
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 6932 13870 6960 14350
rect 7024 13870 7052 15642
rect 7196 15428 7248 15434
rect 7116 15388 7196 15416
rect 7116 15162 7144 15388
rect 7196 15370 7248 15376
rect 7252 15260 7560 15269
rect 7252 15258 7258 15260
rect 7314 15258 7338 15260
rect 7394 15258 7418 15260
rect 7474 15258 7498 15260
rect 7554 15258 7560 15260
rect 7314 15206 7316 15258
rect 7496 15206 7498 15258
rect 7252 15204 7258 15206
rect 7314 15204 7338 15206
rect 7394 15204 7418 15206
rect 7474 15204 7498 15206
rect 7554 15204 7560 15206
rect 7252 15195 7560 15204
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 7668 15094 7696 16594
rect 7944 16028 7972 17478
rect 8128 16658 8156 17682
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8024 16040 8076 16046
rect 7944 16000 8024 16028
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7852 15570 7880 15846
rect 7840 15564 7892 15570
rect 7840 15506 7892 15512
rect 7380 15088 7432 15094
rect 7380 15030 7432 15036
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7208 14618 7236 14962
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 7392 14362 7420 15030
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 7116 14334 7420 14362
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6000 13320 6052 13326
rect 6276 13320 6328 13326
rect 6000 13262 6052 13268
rect 6104 13280 6276 13308
rect 6012 12714 6040 13262
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 6104 12306 6132 13280
rect 6276 13262 6328 13268
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6288 12434 6316 13126
rect 6380 12782 6408 13466
rect 6460 13456 6512 13462
rect 6512 13416 6592 13444
rect 6460 13398 6512 13404
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6196 12406 6316 12434
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 6196 12050 6224 12406
rect 6380 12322 6408 12582
rect 6380 12294 6500 12322
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6104 12022 6224 12050
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5920 11354 5948 11698
rect 5908 11348 5960 11354
rect 5908 11290 5960 11296
rect 6104 11218 6132 12022
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5828 9450 5856 11086
rect 5920 10810 5948 11086
rect 6380 11014 6408 12106
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 6012 10742 6040 10950
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 6092 10736 6144 10742
rect 6092 10678 6144 10684
rect 6104 10266 6132 10678
rect 6472 10674 6500 12294
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6196 10266 6224 10542
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6380 10062 6408 10542
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 6564 9178 6592 13416
rect 6932 13394 6960 13806
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6656 12238 6684 12786
rect 6840 12714 6868 13262
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 7012 12640 7064 12646
rect 6932 12588 7012 12594
rect 6932 12582 7064 12588
rect 6932 12566 7052 12582
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6644 11756 6696 11762
rect 6748 11744 6776 12242
rect 6932 12238 6960 12566
rect 7116 12238 7144 14334
rect 7252 14172 7560 14181
rect 7252 14170 7258 14172
rect 7314 14170 7338 14172
rect 7394 14170 7418 14172
rect 7474 14170 7498 14172
rect 7554 14170 7560 14172
rect 7314 14118 7316 14170
rect 7496 14118 7498 14170
rect 7252 14116 7258 14118
rect 7314 14116 7338 14118
rect 7394 14116 7418 14118
rect 7474 14116 7498 14118
rect 7554 14116 7560 14118
rect 7252 14107 7560 14116
rect 7760 14006 7788 14486
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7392 13462 7420 13670
rect 7380 13456 7432 13462
rect 7380 13398 7432 13404
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7252 13084 7560 13093
rect 7252 13082 7258 13084
rect 7314 13082 7338 13084
rect 7394 13082 7418 13084
rect 7474 13082 7498 13084
rect 7554 13082 7560 13084
rect 7314 13030 7316 13082
rect 7496 13030 7498 13082
rect 7252 13028 7258 13030
rect 7314 13028 7338 13030
rect 7394 13028 7418 13030
rect 7474 13028 7498 13030
rect 7554 13028 7560 13030
rect 7252 13019 7560 13028
rect 7668 12918 7696 13330
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7760 12850 7788 13262
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7852 12374 7880 15506
rect 7944 13734 7972 16000
rect 8024 15982 8076 15988
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 8036 15706 8064 15846
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 8036 12850 8064 15302
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 7840 12368 7892 12374
rect 7840 12310 7892 12316
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6696 11716 6776 11744
rect 6644 11698 6696 11704
rect 6656 11234 6684 11698
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6748 11354 6776 11494
rect 6932 11354 6960 12038
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6656 11206 6776 11234
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6656 10538 6684 11086
rect 6748 10810 6776 11206
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6748 10713 6776 10746
rect 6734 10704 6790 10713
rect 6734 10639 6790 10648
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6644 10532 6696 10538
rect 6644 10474 6696 10480
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6748 9722 6776 10066
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6840 9586 6868 9998
rect 6932 9722 6960 10610
rect 7024 10470 7052 11698
rect 7116 11286 7144 12174
rect 7252 11996 7560 12005
rect 7252 11994 7258 11996
rect 7314 11994 7338 11996
rect 7394 11994 7418 11996
rect 7474 11994 7498 11996
rect 7554 11994 7560 11996
rect 7314 11942 7316 11994
rect 7496 11942 7498 11994
rect 7252 11940 7258 11942
rect 7314 11940 7338 11942
rect 7394 11940 7418 11942
rect 7474 11940 7498 11942
rect 7554 11940 7560 11942
rect 7252 11931 7560 11940
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 7208 10996 7236 11630
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 7564 11144 7616 11150
rect 7616 11092 7880 11098
rect 7564 11086 7880 11092
rect 7576 11070 7880 11086
rect 7116 10968 7236 10996
rect 7116 10810 7144 10968
rect 7252 10908 7560 10917
rect 7252 10906 7258 10908
rect 7314 10906 7338 10908
rect 7394 10906 7418 10908
rect 7474 10906 7498 10908
rect 7554 10906 7560 10908
rect 7314 10854 7316 10906
rect 7496 10854 7498 10906
rect 7252 10852 7258 10854
rect 7314 10852 7338 10854
rect 7394 10852 7418 10854
rect 7474 10852 7498 10854
rect 7554 10852 7560 10854
rect 7252 10843 7560 10852
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7576 10674 7604 10746
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7208 10470 7236 10610
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7024 9994 7052 10406
rect 7576 10266 7604 10610
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7576 10062 7604 10202
rect 7760 10062 7788 10406
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6458 8528 6514 8537
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 6276 8492 6328 8498
rect 6748 8514 6776 8774
rect 6748 8498 6868 8514
rect 6748 8492 6880 8498
rect 6748 8486 6828 8492
rect 6458 8463 6514 8472
rect 6276 8434 6328 8440
rect 5828 7886 5856 8434
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 5920 7002 5948 7754
rect 6104 7410 6132 7822
rect 6288 7750 6316 8434
rect 6472 7886 6500 8463
rect 6828 8434 6880 8440
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5276 5914 5304 6190
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5552 5370 5580 5714
rect 5644 5370 5672 6258
rect 5828 6186 5856 6734
rect 6104 6458 6132 7346
rect 6288 6798 6316 7686
rect 6380 7410 6408 7822
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6564 7342 6592 7822
rect 6656 7478 6684 8366
rect 6840 8294 6868 8434
rect 7024 8430 7052 9930
rect 7252 9820 7560 9829
rect 7252 9818 7258 9820
rect 7314 9818 7338 9820
rect 7394 9818 7418 9820
rect 7474 9818 7498 9820
rect 7554 9818 7560 9820
rect 7314 9766 7316 9818
rect 7496 9766 7498 9818
rect 7252 9764 7258 9766
rect 7314 9764 7338 9766
rect 7394 9764 7418 9766
rect 7474 9764 7498 9766
rect 7554 9764 7560 9766
rect 7252 9755 7560 9764
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 5816 6180 5868 6186
rect 5816 6122 5868 6128
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5644 4758 5672 5170
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5736 4622 5764 5782
rect 5828 4826 5856 6122
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5920 4622 5948 5714
rect 6196 5710 6224 6054
rect 6472 5778 6500 6734
rect 6564 6458 6592 7278
rect 6656 7002 6684 7414
rect 6840 7410 6868 8230
rect 6932 7546 6960 8298
rect 7116 8090 7144 8842
rect 7252 8732 7560 8741
rect 7252 8730 7258 8732
rect 7314 8730 7338 8732
rect 7394 8730 7418 8732
rect 7474 8730 7498 8732
rect 7554 8730 7560 8732
rect 7314 8678 7316 8730
rect 7496 8678 7498 8730
rect 7252 8676 7258 8678
rect 7314 8676 7338 8678
rect 7394 8676 7418 8678
rect 7474 8676 7498 8678
rect 7554 8676 7560 8678
rect 7252 8667 7560 8676
rect 7668 8634 7696 9658
rect 7748 9104 7800 9110
rect 7748 9046 7800 9052
rect 7760 8634 7788 9046
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7668 8022 7696 8366
rect 7760 8022 7788 8434
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7252 7644 7560 7653
rect 7252 7642 7258 7644
rect 7314 7642 7338 7644
rect 7394 7642 7418 7644
rect 7474 7642 7498 7644
rect 7554 7642 7560 7644
rect 7314 7590 7316 7642
rect 7496 7590 7498 7642
rect 7252 7588 7258 7590
rect 7314 7588 7338 7590
rect 7394 7588 7418 7590
rect 7474 7588 7498 7590
rect 7554 7588 7560 7590
rect 7252 7579 7560 7588
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 7760 7410 7788 7958
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 7852 6730 7880 11070
rect 7944 10062 7972 11154
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7944 7546 7972 9998
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 8036 7886 8064 8434
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 8036 7478 8064 7686
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6656 5710 6684 6598
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6932 5914 6960 6190
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6196 5370 6224 5646
rect 6276 5636 6328 5642
rect 6276 5578 6328 5584
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6104 4826 6132 5170
rect 6288 5166 6316 5578
rect 6748 5302 6776 5646
rect 7024 5574 7052 6666
rect 7252 6556 7560 6565
rect 7252 6554 7258 6556
rect 7314 6554 7338 6556
rect 7394 6554 7418 6556
rect 7474 6554 7498 6556
rect 7554 6554 7560 6556
rect 7314 6502 7316 6554
rect 7496 6502 7498 6554
rect 7252 6500 7258 6502
rect 7314 6500 7338 6502
rect 7394 6500 7418 6502
rect 7474 6500 7498 6502
rect 7554 6500 7560 6502
rect 7252 6491 7560 6500
rect 8128 6202 8156 14486
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 8220 13870 8248 14214
rect 8312 14074 8340 14214
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8220 13326 8248 13806
rect 8496 13462 8524 18022
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 8760 17060 8812 17066
rect 8760 17002 8812 17008
rect 8772 16590 8800 17002
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 8864 15910 8892 16934
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8956 16182 8984 16526
rect 8944 16176 8996 16182
rect 8944 16118 8996 16124
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8864 15026 8892 15302
rect 8852 15020 8904 15026
rect 8852 14962 8904 14968
rect 8956 14074 8984 16118
rect 9048 15706 9076 17138
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9416 15570 9444 18770
rect 9692 18358 9720 19382
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 9508 16522 9536 18226
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9692 17678 9720 18022
rect 9784 17882 9812 20352
rect 9876 20330 9904 21490
rect 9968 20806 9996 21830
rect 10060 21622 10088 21966
rect 10152 21690 10180 22986
rect 10244 22098 10272 23054
rect 10888 22982 10916 24754
rect 11060 24744 11112 24750
rect 11060 24686 11112 24692
rect 11072 24410 11100 24686
rect 11060 24404 11112 24410
rect 11060 24346 11112 24352
rect 11244 24268 11296 24274
rect 11244 24210 11296 24216
rect 10876 22976 10928 22982
rect 10876 22918 10928 22924
rect 11256 22710 11284 24210
rect 11440 24206 11468 26726
rect 11796 26376 11848 26382
rect 11796 26318 11848 26324
rect 11808 25498 11836 26318
rect 11888 26240 11940 26246
rect 11888 26182 11940 26188
rect 11796 25492 11848 25498
rect 11796 25434 11848 25440
rect 11520 24608 11572 24614
rect 11520 24550 11572 24556
rect 11532 24342 11560 24550
rect 11704 24404 11756 24410
rect 11704 24346 11756 24352
rect 11520 24336 11572 24342
rect 11520 24278 11572 24284
rect 11532 24206 11560 24278
rect 11428 24200 11480 24206
rect 11428 24142 11480 24148
rect 11520 24200 11572 24206
rect 11520 24142 11572 24148
rect 11520 23724 11572 23730
rect 11520 23666 11572 23672
rect 11428 22976 11480 22982
rect 11428 22918 11480 22924
rect 11244 22704 11296 22710
rect 11244 22646 11296 22652
rect 11152 22636 11204 22642
rect 11152 22578 11204 22584
rect 10324 22568 10376 22574
rect 10324 22510 10376 22516
rect 10232 22092 10284 22098
rect 10232 22034 10284 22040
rect 10336 21962 10364 22510
rect 10968 22432 11020 22438
rect 10968 22374 11020 22380
rect 10403 22332 10711 22341
rect 10403 22330 10409 22332
rect 10465 22330 10489 22332
rect 10545 22330 10569 22332
rect 10625 22330 10649 22332
rect 10705 22330 10711 22332
rect 10465 22278 10467 22330
rect 10647 22278 10649 22330
rect 10403 22276 10409 22278
rect 10465 22276 10489 22278
rect 10545 22276 10569 22278
rect 10625 22276 10649 22278
rect 10705 22276 10711 22278
rect 10403 22267 10711 22276
rect 10600 22024 10652 22030
rect 10652 21972 10732 21978
rect 10600 21966 10732 21972
rect 10232 21956 10284 21962
rect 10232 21898 10284 21904
rect 10324 21956 10376 21962
rect 10612 21950 10732 21966
rect 10980 21962 11008 22374
rect 10324 21898 10376 21904
rect 10140 21684 10192 21690
rect 10140 21626 10192 21632
rect 10048 21616 10100 21622
rect 10048 21558 10100 21564
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 10152 21146 10180 21286
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 9864 20324 9916 20330
rect 9864 20266 9916 20272
rect 9968 20058 9996 20470
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9968 18698 9996 19994
rect 10244 19334 10272 21898
rect 10336 21486 10364 21898
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 10612 21622 10640 21830
rect 10600 21616 10652 21622
rect 10600 21558 10652 21564
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 10704 21332 10732 21950
rect 10968 21956 11020 21962
rect 10968 21898 11020 21904
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 10796 21554 10824 21830
rect 11072 21690 11100 21830
rect 11164 21690 11192 22578
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 11440 21486 11468 22918
rect 11532 22778 11560 23666
rect 11520 22772 11572 22778
rect 11520 22714 11572 22720
rect 11428 21480 11480 21486
rect 11428 21422 11480 21428
rect 10704 21304 10916 21332
rect 10403 21244 10711 21253
rect 10403 21242 10409 21244
rect 10465 21242 10489 21244
rect 10545 21242 10569 21244
rect 10625 21242 10649 21244
rect 10705 21242 10711 21244
rect 10465 21190 10467 21242
rect 10647 21190 10649 21242
rect 10403 21188 10409 21190
rect 10465 21188 10489 21190
rect 10545 21188 10569 21190
rect 10625 21188 10649 21190
rect 10705 21188 10711 21190
rect 10403 21179 10711 21188
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10403 20156 10711 20165
rect 10403 20154 10409 20156
rect 10465 20154 10489 20156
rect 10545 20154 10569 20156
rect 10625 20154 10649 20156
rect 10705 20154 10711 20156
rect 10465 20102 10467 20154
rect 10647 20102 10649 20154
rect 10403 20100 10409 20102
rect 10465 20100 10489 20102
rect 10545 20100 10569 20102
rect 10625 20100 10649 20102
rect 10705 20100 10711 20102
rect 10403 20091 10711 20100
rect 10796 20058 10824 20334
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10152 19306 10272 19334
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 10152 18612 10180 19306
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10232 19168 10284 19174
rect 10232 19110 10284 19116
rect 10244 18766 10272 19110
rect 10336 18766 10364 19246
rect 10403 19068 10711 19077
rect 10403 19066 10409 19068
rect 10465 19066 10489 19068
rect 10545 19066 10569 19068
rect 10625 19066 10649 19068
rect 10705 19066 10711 19068
rect 10465 19014 10467 19066
rect 10647 19014 10649 19066
rect 10403 19012 10409 19014
rect 10465 19012 10489 19014
rect 10545 19012 10569 19014
rect 10625 19012 10649 19014
rect 10705 19012 10711 19014
rect 10403 19003 10711 19012
rect 10796 18970 10824 19994
rect 10888 18970 10916 21304
rect 10968 20324 11020 20330
rect 10968 20266 11020 20272
rect 10980 19854 11008 20266
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11624 20058 11652 20198
rect 11612 20052 11664 20058
rect 11612 19994 11664 20000
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11164 19378 11192 19654
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 10232 18624 10284 18630
rect 10152 18584 10232 18612
rect 10232 18566 10284 18572
rect 10600 18624 10652 18630
rect 10600 18566 10652 18572
rect 10612 18358 10640 18566
rect 10600 18352 10652 18358
rect 10600 18294 10652 18300
rect 10796 18290 10824 18702
rect 10784 18284 10836 18290
rect 10784 18226 10836 18232
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9588 17264 9640 17270
rect 9588 17206 9640 17212
rect 9496 16516 9548 16522
rect 9496 16458 9548 16464
rect 9508 16250 9536 16458
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9508 15502 9536 16186
rect 9496 15496 9548 15502
rect 9496 15438 9548 15444
rect 9600 15366 9628 17206
rect 9784 17134 9812 17818
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 10152 16250 10180 18158
rect 10403 17980 10711 17989
rect 10403 17978 10409 17980
rect 10465 17978 10489 17980
rect 10545 17978 10569 17980
rect 10625 17978 10649 17980
rect 10705 17978 10711 17980
rect 10465 17926 10467 17978
rect 10647 17926 10649 17978
rect 10403 17924 10409 17926
rect 10465 17924 10489 17926
rect 10545 17924 10569 17926
rect 10625 17924 10649 17926
rect 10705 17924 10711 17926
rect 10403 17915 10711 17924
rect 10888 17678 10916 18226
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 10244 17338 10272 17478
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10336 16794 10364 16934
rect 10403 16892 10711 16901
rect 10403 16890 10409 16892
rect 10465 16890 10489 16892
rect 10545 16890 10569 16892
rect 10625 16890 10649 16892
rect 10705 16890 10711 16892
rect 10465 16838 10467 16890
rect 10647 16838 10649 16890
rect 10403 16836 10409 16838
rect 10465 16836 10489 16838
rect 10545 16836 10569 16838
rect 10625 16836 10649 16838
rect 10705 16836 10711 16838
rect 10403 16827 10711 16836
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10796 16658 10824 16934
rect 10888 16794 10916 17614
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11532 17338 11560 17478
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11152 17196 11204 17202
rect 11152 17138 11204 17144
rect 11164 16794 11192 17138
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 10244 15706 10272 15846
rect 10403 15804 10711 15813
rect 10403 15802 10409 15804
rect 10465 15802 10489 15804
rect 10545 15802 10569 15804
rect 10625 15802 10649 15804
rect 10705 15802 10711 15804
rect 10465 15750 10467 15802
rect 10647 15750 10649 15802
rect 10403 15748 10409 15750
rect 10465 15748 10489 15750
rect 10545 15748 10569 15750
rect 10625 15748 10649 15750
rect 10705 15748 10711 15750
rect 10403 15739 10711 15748
rect 11716 15706 11744 24346
rect 11808 24206 11836 25434
rect 11900 24954 11928 26182
rect 11980 25832 12032 25838
rect 11980 25774 12032 25780
rect 11992 25498 12020 25774
rect 12164 25696 12216 25702
rect 12164 25638 12216 25644
rect 12176 25498 12204 25638
rect 12268 25498 12296 26726
rect 12348 25968 12400 25974
rect 12452 25956 12480 26726
rect 12898 26480 12954 26489
rect 12898 26415 12954 26424
rect 12532 26240 12584 26246
rect 12532 26182 12584 26188
rect 12544 25974 12572 26182
rect 12400 25928 12480 25956
rect 12532 25968 12584 25974
rect 12348 25910 12400 25916
rect 12532 25910 12584 25916
rect 12624 25696 12676 25702
rect 12624 25638 12676 25644
rect 11980 25492 12032 25498
rect 11980 25434 12032 25440
rect 12164 25492 12216 25498
rect 12164 25434 12216 25440
rect 12256 25492 12308 25498
rect 12256 25434 12308 25440
rect 12636 25226 12664 25638
rect 12624 25220 12676 25226
rect 12624 25162 12676 25168
rect 11888 24948 11940 24954
rect 11888 24890 11940 24896
rect 12348 24744 12400 24750
rect 12348 24686 12400 24692
rect 12360 24206 12388 24686
rect 11796 24200 11848 24206
rect 11796 24142 11848 24148
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 11980 23520 12032 23526
rect 11980 23462 12032 23468
rect 11992 22778 12020 23462
rect 12084 23322 12112 24142
rect 12360 23746 12388 24142
rect 12532 24064 12584 24070
rect 12532 24006 12584 24012
rect 12268 23718 12388 23746
rect 12072 23316 12124 23322
rect 12072 23258 12124 23264
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 11980 22568 12032 22574
rect 11980 22510 12032 22516
rect 11992 21554 12020 22510
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 12084 21486 12112 21966
rect 12268 21486 12296 23718
rect 12544 23662 12572 24006
rect 12532 23656 12584 23662
rect 12532 23598 12584 23604
rect 12624 23656 12676 23662
rect 12624 23598 12676 23604
rect 12636 23186 12664 23598
rect 12808 23316 12860 23322
rect 12808 23258 12860 23264
rect 12624 23180 12676 23186
rect 12624 23122 12676 23128
rect 12820 23118 12848 23258
rect 12912 23118 12940 26415
rect 13464 26246 13492 26998
rect 14004 26988 14056 26994
rect 14004 26930 14056 26936
rect 13912 26376 13964 26382
rect 13912 26318 13964 26324
rect 13452 26240 13504 26246
rect 13452 26182 13504 26188
rect 13176 24948 13228 24954
rect 13176 24890 13228 24896
rect 13084 24608 13136 24614
rect 13084 24550 13136 24556
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 13004 23526 13032 24074
rect 13096 23730 13124 24550
rect 13188 23730 13216 24890
rect 13268 24744 13320 24750
rect 13268 24686 13320 24692
rect 13280 24410 13308 24686
rect 13268 24404 13320 24410
rect 13268 24346 13320 24352
rect 13464 24070 13492 26182
rect 13554 26140 13862 26149
rect 13554 26138 13560 26140
rect 13616 26138 13640 26140
rect 13696 26138 13720 26140
rect 13776 26138 13800 26140
rect 13856 26138 13862 26140
rect 13616 26086 13618 26138
rect 13798 26086 13800 26138
rect 13554 26084 13560 26086
rect 13616 26084 13640 26086
rect 13696 26084 13720 26086
rect 13776 26084 13800 26086
rect 13856 26084 13862 26086
rect 13554 26075 13862 26084
rect 13924 26042 13952 26318
rect 14016 26042 14044 26930
rect 14924 26920 14976 26926
rect 14924 26862 14976 26868
rect 14936 26586 14964 26862
rect 14924 26580 14976 26586
rect 14924 26522 14976 26528
rect 14830 26480 14886 26489
rect 14556 26444 14608 26450
rect 14608 26404 14688 26432
rect 14830 26415 14886 26424
rect 14556 26386 14608 26392
rect 14556 26240 14608 26246
rect 14556 26182 14608 26188
rect 13912 26036 13964 26042
rect 13912 25978 13964 25984
rect 14004 26036 14056 26042
rect 14004 25978 14056 25984
rect 14464 25900 14516 25906
rect 14464 25842 14516 25848
rect 14476 25362 14504 25842
rect 14568 25838 14596 26182
rect 14660 25974 14688 26404
rect 14844 26246 14872 26415
rect 14832 26240 14884 26246
rect 14832 26182 14884 26188
rect 14648 25968 14700 25974
rect 14648 25910 14700 25916
rect 14556 25832 14608 25838
rect 14556 25774 14608 25780
rect 14568 25498 14596 25774
rect 14556 25492 14608 25498
rect 14556 25434 14608 25440
rect 14464 25356 14516 25362
rect 14292 25316 14464 25344
rect 13554 25052 13862 25061
rect 13554 25050 13560 25052
rect 13616 25050 13640 25052
rect 13696 25050 13720 25052
rect 13776 25050 13800 25052
rect 13856 25050 13862 25052
rect 13616 24998 13618 25050
rect 13798 24998 13800 25050
rect 13554 24996 13560 24998
rect 13616 24996 13640 24998
rect 13696 24996 13720 24998
rect 13776 24996 13800 24998
rect 13856 24996 13862 24998
rect 13554 24987 13862 24996
rect 14292 24954 14320 25316
rect 14464 25298 14516 25304
rect 14280 24948 14332 24954
rect 14280 24890 14332 24896
rect 14556 24812 14608 24818
rect 14660 24800 14688 25910
rect 14936 24834 14964 26522
rect 15212 26382 15240 27066
rect 15660 26988 15712 26994
rect 15660 26930 15712 26936
rect 17132 26988 17184 26994
rect 17132 26930 17184 26936
rect 20996 26988 21048 26994
rect 20996 26930 21048 26936
rect 15384 26920 15436 26926
rect 15384 26862 15436 26868
rect 15292 26512 15344 26518
rect 15292 26454 15344 26460
rect 15200 26376 15252 26382
rect 15200 26318 15252 26324
rect 15212 25362 15240 26318
rect 15304 25498 15332 26454
rect 15396 26042 15424 26862
rect 15476 26512 15528 26518
rect 15476 26454 15528 26460
rect 15384 26036 15436 26042
rect 15384 25978 15436 25984
rect 15292 25492 15344 25498
rect 15292 25434 15344 25440
rect 15200 25356 15252 25362
rect 15200 25298 15252 25304
rect 15108 25152 15160 25158
rect 15108 25094 15160 25100
rect 14936 24806 15056 24834
rect 14608 24772 14688 24800
rect 14556 24754 14608 24760
rect 13820 24744 13872 24750
rect 13820 24686 13872 24692
rect 13832 24206 13860 24686
rect 13820 24200 13872 24206
rect 13820 24142 13872 24148
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 14464 24200 14516 24206
rect 14568 24154 14596 24754
rect 14924 24744 14976 24750
rect 14924 24686 14976 24692
rect 14516 24148 14596 24154
rect 14464 24142 14596 24148
rect 13924 24070 13952 24142
rect 14476 24126 14596 24142
rect 13452 24064 13504 24070
rect 13452 24006 13504 24012
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 14096 24064 14148 24070
rect 14096 24006 14148 24012
rect 13554 23964 13862 23973
rect 13554 23962 13560 23964
rect 13616 23962 13640 23964
rect 13696 23962 13720 23964
rect 13776 23962 13800 23964
rect 13856 23962 13862 23964
rect 13616 23910 13618 23962
rect 13798 23910 13800 23962
rect 13554 23908 13560 23910
rect 13616 23908 13640 23910
rect 13696 23908 13720 23910
rect 13776 23908 13800 23910
rect 13856 23908 13862 23910
rect 13554 23899 13862 23908
rect 14108 23866 14136 24006
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 13176 23724 13228 23730
rect 13176 23666 13228 23672
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 13096 23118 13124 23666
rect 12808 23112 12860 23118
rect 12808 23054 12860 23060
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 13084 23112 13136 23118
rect 13084 23054 13136 23060
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 12360 21690 12388 22374
rect 12452 21894 12480 22510
rect 12532 21956 12584 21962
rect 12532 21898 12584 21904
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12452 21690 12480 21830
rect 12348 21684 12400 21690
rect 12348 21626 12400 21632
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 12072 21480 12124 21486
rect 12072 21422 12124 21428
rect 12256 21480 12308 21486
rect 12256 21422 12308 21428
rect 12084 20330 12112 21422
rect 12268 20398 12296 21422
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12452 20602 12480 21286
rect 12544 20942 12572 21898
rect 12820 21622 12848 23054
rect 12992 22228 13044 22234
rect 12992 22170 13044 22176
rect 12808 21616 12860 21622
rect 12728 21576 12808 21604
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 12072 20324 12124 20330
rect 12072 20266 12124 20272
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12176 19174 12204 19246
rect 12268 19174 12296 20334
rect 12452 19922 12480 20334
rect 12532 20324 12584 20330
rect 12532 20266 12584 20272
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 12452 19514 12480 19858
rect 12544 19854 12572 20266
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12164 18692 12216 18698
rect 12164 18634 12216 18640
rect 12176 18358 12204 18634
rect 12164 18352 12216 18358
rect 12164 18294 12216 18300
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11808 17134 11836 17750
rect 12268 17746 12296 19110
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 11888 17264 11940 17270
rect 11888 17206 11940 17212
rect 11900 17134 11928 17206
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 12452 16794 12480 18022
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9954 15056 10010 15065
rect 9954 14991 10010 15000
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 9324 14006 9352 14214
rect 9128 14000 9180 14006
rect 9312 14000 9364 14006
rect 9180 13948 9260 13954
rect 9128 13942 9260 13948
rect 9312 13942 9364 13948
rect 9140 13926 9260 13942
rect 9232 13818 9260 13926
rect 9600 13818 9628 14758
rect 9968 14346 9996 14991
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9876 14006 9904 14214
rect 10152 14006 10180 14758
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10336 14362 10364 15642
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 10403 14716 10711 14725
rect 10403 14714 10409 14716
rect 10465 14714 10489 14716
rect 10545 14714 10569 14716
rect 10625 14714 10649 14716
rect 10705 14714 10711 14716
rect 10465 14662 10467 14714
rect 10647 14662 10649 14714
rect 10403 14660 10409 14662
rect 10465 14660 10489 14662
rect 10545 14660 10569 14662
rect 10625 14660 10649 14662
rect 10705 14660 10711 14662
rect 10403 14651 10711 14660
rect 11072 14618 11100 14894
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 10692 14544 10744 14550
rect 10744 14504 11008 14532
rect 10692 14486 10744 14492
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 9232 13790 9628 13818
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 8484 13456 8536 13462
rect 8484 13398 8536 13404
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8220 12918 8248 13262
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8208 12912 8260 12918
rect 8208 12854 8260 12860
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8312 12442 8340 12718
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8404 12238 8432 13126
rect 8772 12646 8800 13262
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 9048 12986 9076 13194
rect 9140 12986 9168 13670
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9416 12764 9444 13194
rect 9600 12918 9628 13790
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9496 12776 9548 12782
rect 9416 12736 9496 12764
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8772 12434 8800 12582
rect 8680 12406 8800 12434
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8496 10266 8524 10610
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8496 9586 8524 10202
rect 8588 9926 8616 11154
rect 8680 10810 8708 12406
rect 9416 12238 9444 12736
rect 9496 12718 9548 12724
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9784 12306 9812 12650
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 10152 12238 10180 13942
rect 10244 13870 10272 14350
rect 10336 14346 10456 14362
rect 10336 14340 10468 14346
rect 10336 14334 10416 14340
rect 10416 14282 10468 14288
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 10336 13870 10364 14214
rect 10612 14074 10640 14418
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10980 13988 11008 14504
rect 11256 14346 11284 14894
rect 11348 14482 11376 15302
rect 11440 15162 11468 15438
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11716 15094 11744 15302
rect 12084 15094 12112 16390
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 12072 15088 12124 15094
rect 12072 15030 12124 15036
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11440 14498 11468 14962
rect 11440 14482 11652 14498
rect 11336 14476 11388 14482
rect 11440 14476 11664 14482
rect 11440 14470 11612 14476
rect 11336 14418 11388 14424
rect 11612 14418 11664 14424
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 11152 14000 11204 14006
rect 10980 13960 11152 13988
rect 11152 13942 11204 13948
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10244 12306 10272 13806
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9140 11354 9168 12038
rect 9416 11626 9444 12174
rect 10336 11898 10364 13806
rect 10403 13628 10711 13637
rect 10403 13626 10409 13628
rect 10465 13626 10489 13628
rect 10545 13626 10569 13628
rect 10625 13626 10649 13628
rect 10705 13626 10711 13628
rect 10465 13574 10467 13626
rect 10647 13574 10649 13626
rect 10403 13572 10409 13574
rect 10465 13572 10489 13574
rect 10545 13572 10569 13574
rect 10625 13572 10649 13574
rect 10705 13572 10711 13574
rect 10403 13563 10711 13572
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10403 12540 10711 12549
rect 10403 12538 10409 12540
rect 10465 12538 10489 12540
rect 10545 12538 10569 12540
rect 10625 12538 10649 12540
rect 10705 12538 10711 12540
rect 10465 12486 10467 12538
rect 10647 12486 10649 12538
rect 10403 12484 10409 12486
rect 10465 12484 10489 12486
rect 10545 12484 10569 12486
rect 10625 12484 10649 12486
rect 10705 12484 10711 12486
rect 10403 12475 10711 12484
rect 10796 12170 10824 12582
rect 10784 12164 10836 12170
rect 10784 12106 10836 12112
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8864 10674 8892 10950
rect 8956 10810 8984 11154
rect 9600 11150 9628 11494
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8680 10062 8708 10610
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8680 9586 8708 9998
rect 8772 9722 8800 10542
rect 8864 9722 8892 10610
rect 9048 10266 9076 10610
rect 9140 10538 9168 10950
rect 9324 10674 9352 11018
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 9692 10470 9720 10950
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9692 10282 9720 10406
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9600 10254 9720 10282
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8496 9178 8524 9522
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8680 9110 8708 9522
rect 9416 9178 9444 9998
rect 9600 9722 9628 10254
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9692 9722 9720 10066
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8404 8634 8432 8910
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8404 8537 8432 8570
rect 8390 8528 8446 8537
rect 8772 8498 8800 9046
rect 8390 8463 8446 8472
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8772 7886 8800 8434
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8312 6458 8340 6734
rect 8496 6458 8524 6734
rect 8680 6730 8708 7346
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9416 6798 9444 7278
rect 9600 6798 9628 7346
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 9416 6390 9444 6598
rect 9404 6384 9456 6390
rect 9404 6326 9456 6332
rect 8036 6174 8156 6202
rect 8852 6180 8904 6186
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7252 5468 7560 5477
rect 7252 5466 7258 5468
rect 7314 5466 7338 5468
rect 7394 5466 7418 5468
rect 7474 5466 7498 5468
rect 7554 5466 7560 5468
rect 7314 5414 7316 5466
rect 7496 5414 7498 5466
rect 7252 5412 7258 5414
rect 7314 5412 7338 5414
rect 7394 5412 7418 5414
rect 7474 5412 7498 5414
rect 7554 5412 7560 5414
rect 7252 5403 7560 5412
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6276 5160 6328 5166
rect 6276 5102 6328 5108
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6288 4690 6316 5102
rect 7024 4826 7052 5170
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 6288 4282 6316 4626
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 7116 4146 7144 4558
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7252 4380 7560 4389
rect 7252 4378 7258 4380
rect 7314 4378 7338 4380
rect 7394 4378 7418 4380
rect 7474 4378 7498 4380
rect 7554 4378 7560 4380
rect 7314 4326 7316 4378
rect 7496 4326 7498 4378
rect 7252 4324 7258 4326
rect 7314 4324 7338 4326
rect 7394 4324 7418 4326
rect 7474 4324 7498 4326
rect 7554 4324 7560 4326
rect 7252 4315 7560 4324
rect 7668 4282 7696 4422
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7116 3738 7144 4082
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7944 3738 7972 4014
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 8036 3602 8064 6174
rect 8852 6122 8904 6128
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8128 5914 8156 6054
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8128 5370 8156 5510
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8864 5302 8892 6122
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8956 5914 8984 6054
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8956 5250 8984 5510
rect 9140 5250 9168 5850
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9232 5574 9260 5646
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9232 5370 9260 5510
rect 9508 5370 9536 5714
rect 9600 5574 9628 6734
rect 9692 5846 9720 8366
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9784 5760 9812 11834
rect 10784 11824 10836 11830
rect 10784 11766 10836 11772
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 9876 10810 9904 11698
rect 10336 11200 10364 11698
rect 10403 11452 10711 11461
rect 10403 11450 10409 11452
rect 10465 11450 10489 11452
rect 10545 11450 10569 11452
rect 10625 11450 10649 11452
rect 10705 11450 10711 11452
rect 10465 11398 10467 11450
rect 10647 11398 10649 11450
rect 10403 11396 10409 11398
rect 10465 11396 10489 11398
rect 10545 11396 10569 11398
rect 10625 11396 10649 11398
rect 10705 11396 10711 11398
rect 10403 11387 10711 11396
rect 10796 11354 10824 11766
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10416 11212 10468 11218
rect 10336 11172 10416 11200
rect 10416 11154 10468 11160
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9862 10568 9918 10577
rect 9862 10503 9918 10512
rect 9876 10266 9904 10503
rect 9968 10470 9996 10610
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9968 10062 9996 10406
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 9864 9988 9916 9994
rect 9864 9930 9916 9936
rect 9876 9586 9904 9930
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9968 8974 9996 9998
rect 10060 9654 10088 11018
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 10152 9586 10180 10678
rect 10428 10674 10456 11154
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10796 10674 10824 10950
rect 10980 10810 11008 12786
rect 11072 11150 11100 13466
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 11164 11830 11192 12242
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11256 11218 11284 11562
rect 11348 11218 11376 12854
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11900 11830 11928 12582
rect 11888 11824 11940 11830
rect 11888 11766 11940 11772
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11624 11218 11652 11698
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10244 10266 10272 10610
rect 10704 10577 10732 10610
rect 10690 10568 10746 10577
rect 10690 10503 10746 10512
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10403 10364 10711 10373
rect 10403 10362 10409 10364
rect 10465 10362 10489 10364
rect 10545 10362 10569 10364
rect 10625 10362 10649 10364
rect 10705 10362 10711 10364
rect 10465 10310 10467 10362
rect 10647 10310 10649 10362
rect 10403 10308 10409 10310
rect 10465 10308 10489 10310
rect 10545 10308 10569 10310
rect 10625 10308 10649 10310
rect 10705 10308 10711 10310
rect 10403 10299 10711 10308
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10796 10146 10824 10406
rect 10704 10118 10824 10146
rect 10704 10062 10732 10118
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10336 9586 10364 9998
rect 10428 9586 10456 9998
rect 10600 9988 10652 9994
rect 10600 9930 10652 9936
rect 10612 9602 10640 9930
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10704 9722 10732 9862
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10796 9602 10824 9658
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10612 9574 10824 9602
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 10336 8906 10364 9522
rect 10428 9382 10456 9522
rect 10612 9518 10640 9574
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10403 9276 10711 9285
rect 10403 9274 10409 9276
rect 10465 9274 10489 9276
rect 10545 9274 10569 9276
rect 10625 9274 10649 9276
rect 10705 9274 10711 9276
rect 10465 9222 10467 9274
rect 10647 9222 10649 9274
rect 10403 9220 10409 9222
rect 10465 9220 10489 9222
rect 10545 9220 10569 9222
rect 10625 9220 10649 9222
rect 10705 9220 10711 9222
rect 10403 9211 10711 9220
rect 10888 9178 10916 9386
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10876 8900 10928 8906
rect 10876 8842 10928 8848
rect 10403 8188 10711 8197
rect 10403 8186 10409 8188
rect 10465 8186 10489 8188
rect 10545 8186 10569 8188
rect 10625 8186 10649 8188
rect 10705 8186 10711 8188
rect 10465 8134 10467 8186
rect 10647 8134 10649 8186
rect 10403 8132 10409 8134
rect 10465 8132 10489 8134
rect 10545 8132 10569 8134
rect 10625 8132 10649 8134
rect 10705 8132 10711 8134
rect 10403 8123 10711 8132
rect 10888 8090 10916 8842
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10403 7100 10711 7109
rect 10403 7098 10409 7100
rect 10465 7098 10489 7100
rect 10545 7098 10569 7100
rect 10625 7098 10649 7100
rect 10705 7098 10711 7100
rect 10465 7046 10467 7098
rect 10647 7046 10649 7098
rect 10403 7044 10409 7046
rect 10465 7044 10489 7046
rect 10545 7044 10569 7046
rect 10625 7044 10649 7046
rect 10705 7044 10711 7046
rect 10403 7035 10711 7044
rect 10980 6882 11008 9590
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 11060 9444 11112 9450
rect 11164 9432 11192 9522
rect 11112 9404 11192 9432
rect 11060 9386 11112 9392
rect 11060 8628 11112 8634
rect 11164 8616 11192 9404
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11348 9178 11376 9318
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11112 8588 11192 8616
rect 11060 8570 11112 8576
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11256 8090 11284 8230
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11624 7546 11652 8774
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11716 7410 11744 8434
rect 11808 7818 11836 8774
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 11808 7410 11836 7754
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11900 7002 11928 7142
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 10888 6866 11008 6882
rect 10876 6860 11008 6866
rect 10928 6854 11008 6860
rect 10876 6802 10928 6808
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10152 5914 10180 6734
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10336 6202 10364 6258
rect 10888 6254 10916 6802
rect 11992 6746 12020 14418
rect 12268 14414 12296 15030
rect 12360 14550 12388 15506
rect 12544 15434 12572 18838
rect 12728 18766 12756 21576
rect 12808 21558 12860 21564
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 12820 19718 12848 21422
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12912 20058 12940 20402
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12728 18290 12756 18702
rect 12820 18698 12848 19654
rect 12912 19378 12940 19790
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12636 17746 12664 18226
rect 12728 17785 12756 18226
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12714 17776 12770 17785
rect 12624 17740 12676 17746
rect 12714 17711 12770 17720
rect 12624 17682 12676 17688
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12728 16522 12756 17274
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12820 14958 12848 18022
rect 12912 17202 12940 19314
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12900 17060 12952 17066
rect 12900 17002 12952 17008
rect 12912 16794 12940 17002
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12360 13802 12388 14486
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12544 12986 12572 13262
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12084 12850 12112 12922
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12452 12442 12480 12718
rect 12440 12436 12492 12442
rect 12636 12424 12664 12718
rect 12716 12436 12768 12442
rect 12636 12396 12716 12424
rect 12440 12378 12492 12384
rect 12716 12378 12768 12384
rect 13004 12170 13032 22170
rect 13188 22098 13216 23666
rect 13452 23520 13504 23526
rect 13452 23462 13504 23468
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 13176 22092 13228 22098
rect 13176 22034 13228 22040
rect 13188 21486 13216 22034
rect 13372 21554 13400 23122
rect 13464 21570 13492 23462
rect 13554 22876 13862 22885
rect 13554 22874 13560 22876
rect 13616 22874 13640 22876
rect 13696 22874 13720 22876
rect 13776 22874 13800 22876
rect 13856 22874 13862 22876
rect 13616 22822 13618 22874
rect 13798 22822 13800 22874
rect 13554 22820 13560 22822
rect 13616 22820 13640 22822
rect 13696 22820 13720 22822
rect 13776 22820 13800 22822
rect 13856 22820 13862 22822
rect 13554 22811 13862 22820
rect 14004 22432 14056 22438
rect 14004 22374 14056 22380
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 13554 21788 13862 21797
rect 13554 21786 13560 21788
rect 13616 21786 13640 21788
rect 13696 21786 13720 21788
rect 13776 21786 13800 21788
rect 13856 21786 13862 21788
rect 13616 21734 13618 21786
rect 13798 21734 13800 21786
rect 13554 21732 13560 21734
rect 13616 21732 13640 21734
rect 13696 21732 13720 21734
rect 13776 21732 13800 21734
rect 13856 21732 13862 21734
rect 13554 21723 13862 21732
rect 13924 21622 13952 21830
rect 13544 21616 13596 21622
rect 13464 21564 13544 21570
rect 13464 21558 13596 21564
rect 13912 21616 13964 21622
rect 13912 21558 13964 21564
rect 13360 21548 13412 21554
rect 13360 21490 13412 21496
rect 13464 21542 13584 21558
rect 13176 21480 13228 21486
rect 13176 21422 13228 21428
rect 13084 20868 13136 20874
rect 13084 20810 13136 20816
rect 13096 20398 13124 20810
rect 13084 20392 13136 20398
rect 13084 20334 13136 20340
rect 13360 19984 13412 19990
rect 13360 19926 13412 19932
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13280 19242 13308 19790
rect 13268 19236 13320 19242
rect 13268 19178 13320 19184
rect 13280 18834 13308 19178
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 13372 18714 13400 19926
rect 13280 18686 13400 18714
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 13188 17338 13216 17682
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 13280 16998 13308 18686
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13372 17746 13400 18158
rect 13464 18086 13492 21542
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 13554 20700 13862 20709
rect 13554 20698 13560 20700
rect 13616 20698 13640 20700
rect 13696 20698 13720 20700
rect 13776 20698 13800 20700
rect 13856 20698 13862 20700
rect 13616 20646 13618 20698
rect 13798 20646 13800 20698
rect 13554 20644 13560 20646
rect 13616 20644 13640 20646
rect 13696 20644 13720 20646
rect 13776 20644 13800 20646
rect 13856 20644 13862 20646
rect 13554 20635 13862 20644
rect 13554 19612 13862 19621
rect 13554 19610 13560 19612
rect 13616 19610 13640 19612
rect 13696 19610 13720 19612
rect 13776 19610 13800 19612
rect 13856 19610 13862 19612
rect 13616 19558 13618 19610
rect 13798 19558 13800 19610
rect 13554 19556 13560 19558
rect 13616 19556 13640 19558
rect 13696 19556 13720 19558
rect 13776 19556 13800 19558
rect 13856 19556 13862 19558
rect 13554 19547 13862 19556
rect 13554 18524 13862 18533
rect 13554 18522 13560 18524
rect 13616 18522 13640 18524
rect 13696 18522 13720 18524
rect 13776 18522 13800 18524
rect 13856 18522 13862 18524
rect 13616 18470 13618 18522
rect 13798 18470 13800 18522
rect 13554 18468 13560 18470
rect 13616 18468 13640 18470
rect 13696 18468 13720 18470
rect 13776 18468 13800 18470
rect 13856 18468 13862 18470
rect 13554 18459 13862 18468
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13648 17882 13676 18158
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 13372 17134 13400 17682
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13464 17134 13492 17478
rect 13554 17436 13862 17445
rect 13554 17434 13560 17436
rect 13616 17434 13640 17436
rect 13696 17434 13720 17436
rect 13776 17434 13800 17436
rect 13856 17434 13862 17436
rect 13616 17382 13618 17434
rect 13798 17382 13800 17434
rect 13554 17380 13560 17382
rect 13616 17380 13640 17382
rect 13696 17380 13720 17382
rect 13776 17380 13800 17382
rect 13856 17380 13862 17382
rect 13554 17371 13862 17380
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 13280 16794 13308 16934
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13554 16348 13862 16357
rect 13554 16346 13560 16348
rect 13616 16346 13640 16348
rect 13696 16346 13720 16348
rect 13776 16346 13800 16348
rect 13856 16346 13862 16348
rect 13616 16294 13618 16346
rect 13798 16294 13800 16346
rect 13554 16292 13560 16294
rect 13616 16292 13640 16294
rect 13696 16292 13720 16294
rect 13776 16292 13800 16294
rect 13856 16292 13862 16294
rect 13554 16283 13862 16292
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13464 14822 13492 15302
rect 13554 15260 13862 15269
rect 13554 15258 13560 15260
rect 13616 15258 13640 15260
rect 13696 15258 13720 15260
rect 13776 15258 13800 15260
rect 13856 15258 13862 15260
rect 13616 15206 13618 15258
rect 13798 15206 13800 15258
rect 13554 15204 13560 15206
rect 13616 15204 13640 15206
rect 13696 15204 13720 15206
rect 13776 15204 13800 15206
rect 13856 15204 13862 15206
rect 13554 15195 13862 15204
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 13188 12986 13216 13262
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 13188 12306 13216 12650
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12360 11830 12388 12038
rect 13188 11830 13216 12242
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 12360 11082 12388 11766
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12360 9674 12388 11018
rect 12176 9646 12388 9674
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 12084 8498 12112 8978
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 12084 7886 12112 8434
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 11900 6718 12020 6746
rect 12176 6730 12204 9646
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 13004 9178 13032 9454
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12360 8498 12388 8774
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12164 6724 12216 6730
rect 11900 6458 11928 6718
rect 12164 6666 12216 6672
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 10244 6174 10364 6202
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10048 5772 10100 5778
rect 9784 5732 10048 5760
rect 10048 5714 10100 5720
rect 9680 5704 9732 5710
rect 9732 5664 9904 5692
rect 9680 5646 9732 5652
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9692 5370 9720 5510
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 8956 5228 9168 5250
rect 8956 5222 9036 5228
rect 9088 5222 9168 5228
rect 9036 5170 9088 5176
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8864 4690 8892 4966
rect 8956 4826 8984 4966
rect 9140 4826 9168 5222
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9324 4826 9352 5170
rect 9508 4826 9536 5306
rect 9772 5296 9824 5302
rect 9772 5238 9824 5244
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 5908 3460 5960 3466
rect 5908 3402 5960 3408
rect 5920 3194 5948 3402
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7252 3292 7560 3301
rect 7252 3290 7258 3292
rect 7314 3290 7338 3292
rect 7394 3290 7418 3292
rect 7474 3290 7498 3292
rect 7554 3290 7560 3292
rect 7314 3238 7316 3290
rect 7496 3238 7498 3290
rect 7252 3236 7258 3238
rect 7314 3236 7338 3238
rect 7394 3236 7418 3238
rect 7474 3236 7498 3238
rect 7554 3236 7560 3238
rect 7252 3227 7560 3236
rect 7668 3194 7696 3334
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 8036 2990 8064 3538
rect 9324 3126 9352 4150
rect 9416 4010 9444 4558
rect 9692 4486 9720 5170
rect 9784 4690 9812 5238
rect 9876 5166 9904 5664
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9968 5234 9996 5510
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9692 4214 9720 4422
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9416 3534 9444 3946
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9692 3194 9720 4150
rect 9784 3602 9812 4626
rect 10060 4146 10088 4762
rect 10244 4214 10272 6174
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10336 5574 10364 6054
rect 10403 6012 10711 6021
rect 10403 6010 10409 6012
rect 10465 6010 10489 6012
rect 10545 6010 10569 6012
rect 10625 6010 10649 6012
rect 10705 6010 10711 6012
rect 10465 5958 10467 6010
rect 10647 5958 10649 6010
rect 10403 5956 10409 5958
rect 10465 5956 10489 5958
rect 10545 5956 10569 5958
rect 10625 5956 10649 5958
rect 10705 5956 10711 5958
rect 10403 5947 10711 5956
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10704 5302 10732 5714
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 10403 4924 10711 4933
rect 10403 4922 10409 4924
rect 10465 4922 10489 4924
rect 10545 4922 10569 4924
rect 10625 4922 10649 4924
rect 10705 4922 10711 4924
rect 10465 4870 10467 4922
rect 10647 4870 10649 4922
rect 10403 4868 10409 4870
rect 10465 4868 10489 4870
rect 10545 4868 10569 4870
rect 10625 4868 10649 4870
rect 10705 4868 10711 4870
rect 10403 4859 10711 4868
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10428 4282 10456 4422
rect 10796 4282 10824 5646
rect 10888 4690 10916 6190
rect 11348 4826 11376 6394
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11624 5370 11652 5850
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 11428 5092 11480 5098
rect 11428 5034 11480 5040
rect 11440 4826 11468 5034
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 10152 3194 10180 3878
rect 10244 3602 10272 4014
rect 10403 3836 10711 3845
rect 10403 3834 10409 3836
rect 10465 3834 10489 3836
rect 10545 3834 10569 3836
rect 10625 3834 10649 3836
rect 10705 3834 10711 3836
rect 10465 3782 10467 3834
rect 10647 3782 10649 3834
rect 10403 3780 10409 3782
rect 10465 3780 10489 3782
rect 10545 3780 10569 3782
rect 10625 3780 10649 3782
rect 10705 3780 10711 3782
rect 10403 3771 10711 3780
rect 10888 3602 10916 4626
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11164 4282 11192 4490
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11900 4010 11928 6190
rect 12176 4622 12204 6666
rect 12452 6458 12480 7346
rect 12544 7342 12572 7890
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12728 7002 12756 7822
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12912 6934 12940 7890
rect 13004 7886 13032 8434
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13188 7478 13216 8434
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13280 8022 13308 8230
rect 13268 8016 13320 8022
rect 13268 7958 13320 7964
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12544 5778 12572 6598
rect 12820 5914 12848 6598
rect 12912 6390 12940 6870
rect 13004 6798 13032 7346
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 13004 6458 13032 6734
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 12636 5086 12940 5114
rect 12636 5030 12664 5086
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11808 3738 11836 3878
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 9312 3120 9364 3126
rect 9312 3062 9364 3068
rect 10244 3058 10272 3538
rect 11532 3398 11560 3606
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 11900 2990 11928 3946
rect 11992 3194 12020 4082
rect 12176 3398 12204 4558
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12360 4078 12388 4422
rect 12728 4146 12756 4966
rect 12912 4826 12940 5086
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 13004 4690 13032 5170
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 13004 3738 13032 4626
rect 13096 4282 13124 4966
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 13188 4214 13216 5646
rect 13280 5370 13308 7822
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 13280 5234 13308 5306
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13372 4622 13400 4966
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13176 4208 13228 4214
rect 13176 4150 13228 4156
rect 13464 4146 13492 14758
rect 13554 14172 13862 14181
rect 13554 14170 13560 14172
rect 13616 14170 13640 14172
rect 13696 14170 13720 14172
rect 13776 14170 13800 14172
rect 13856 14170 13862 14172
rect 13616 14118 13618 14170
rect 13798 14118 13800 14170
rect 13554 14116 13560 14118
rect 13616 14116 13640 14118
rect 13696 14116 13720 14118
rect 13776 14116 13800 14118
rect 13856 14116 13862 14118
rect 13554 14107 13862 14116
rect 13924 14006 13952 21286
rect 14016 20942 14044 22374
rect 14372 21956 14424 21962
rect 14372 21898 14424 21904
rect 14464 21956 14516 21962
rect 14464 21898 14516 21904
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 14004 20936 14056 20942
rect 14004 20878 14056 20884
rect 14108 20398 14136 21830
rect 14384 21690 14412 21898
rect 14372 21684 14424 21690
rect 14372 21626 14424 21632
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 14476 19281 14504 21898
rect 14568 20806 14596 24126
rect 14936 23866 14964 24686
rect 14924 23860 14976 23866
rect 14924 23802 14976 23808
rect 14924 23724 14976 23730
rect 14924 23666 14976 23672
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 14740 22568 14792 22574
rect 14740 22510 14792 22516
rect 14752 22030 14780 22510
rect 14844 22234 14872 22714
rect 14832 22228 14884 22234
rect 14832 22170 14884 22176
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 14752 21486 14780 21966
rect 14936 21622 14964 23666
rect 15028 22574 15056 24806
rect 15120 24274 15148 25094
rect 15212 24834 15240 25298
rect 15212 24806 15424 24834
rect 15488 24818 15516 26454
rect 15568 26240 15620 26246
rect 15568 26182 15620 26188
rect 15580 25838 15608 26182
rect 15568 25832 15620 25838
rect 15568 25774 15620 25780
rect 15200 24676 15252 24682
rect 15200 24618 15252 24624
rect 15108 24268 15160 24274
rect 15108 24210 15160 24216
rect 15120 23798 15148 24210
rect 15212 23866 15240 24618
rect 15292 24268 15344 24274
rect 15396 24256 15424 24806
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15396 24228 15516 24256
rect 15292 24210 15344 24216
rect 15200 23860 15252 23866
rect 15200 23802 15252 23808
rect 15108 23792 15160 23798
rect 15108 23734 15160 23740
rect 15304 22710 15332 24210
rect 15488 22982 15516 24228
rect 15568 24064 15620 24070
rect 15568 24006 15620 24012
rect 15580 23866 15608 24006
rect 15568 23860 15620 23866
rect 15568 23802 15620 23808
rect 15476 22976 15528 22982
rect 15476 22918 15528 22924
rect 15292 22704 15344 22710
rect 15292 22646 15344 22652
rect 15568 22636 15620 22642
rect 15568 22578 15620 22584
rect 15016 22568 15068 22574
rect 15016 22510 15068 22516
rect 14924 21616 14976 21622
rect 14924 21558 14976 21564
rect 14740 21480 14792 21486
rect 14740 21422 14792 21428
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14752 20602 14780 21422
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14936 20534 14964 21558
rect 14924 20528 14976 20534
rect 14924 20470 14976 20476
rect 15028 19496 15056 22510
rect 15476 22432 15528 22438
rect 15476 22374 15528 22380
rect 15488 22234 15516 22374
rect 15476 22228 15528 22234
rect 15476 22170 15528 22176
rect 15580 22098 15608 22578
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 15200 21956 15252 21962
rect 15200 21898 15252 21904
rect 15212 21162 15240 21898
rect 15120 21146 15240 21162
rect 15108 21140 15240 21146
rect 15160 21134 15240 21140
rect 15108 21082 15160 21088
rect 15476 20528 15528 20534
rect 15476 20470 15528 20476
rect 14660 19468 15056 19496
rect 14660 19310 14688 19468
rect 15488 19446 15516 20470
rect 15476 19440 15528 19446
rect 15476 19382 15528 19388
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14648 19304 14700 19310
rect 14462 19272 14518 19281
rect 14648 19246 14700 19252
rect 14462 19207 14518 19216
rect 14660 18873 14688 19246
rect 14646 18864 14702 18873
rect 14646 18799 14702 18808
rect 14752 17746 14780 19314
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 15120 18970 15148 19246
rect 15108 18964 15160 18970
rect 15108 18906 15160 18912
rect 15384 18896 15436 18902
rect 15384 18838 15436 18844
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 15396 18766 15424 18838
rect 15016 18760 15068 18766
rect 15016 18702 15068 18708
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15028 18222 15056 18702
rect 15580 18698 15608 18838
rect 15292 18692 15344 18698
rect 15292 18634 15344 18640
rect 15568 18692 15620 18698
rect 15568 18634 15620 18640
rect 15304 18290 15332 18634
rect 15476 18352 15528 18358
rect 15476 18294 15528 18300
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15016 18216 15068 18222
rect 15016 18158 15068 18164
rect 15488 18154 15516 18294
rect 14832 18148 14884 18154
rect 14832 18090 14884 18096
rect 15476 18148 15528 18154
rect 15476 18090 15528 18096
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 14016 17338 14044 17614
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 14016 16046 14044 17138
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14752 16250 14780 16390
rect 14740 16244 14792 16250
rect 14740 16186 14792 16192
rect 14844 16046 14872 18090
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15016 17740 15068 17746
rect 15016 17682 15068 17688
rect 15028 16658 15056 17682
rect 15304 17338 15332 18022
rect 15488 17678 15516 18090
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15292 17128 15344 17134
rect 15120 17076 15292 17082
rect 15120 17070 15344 17076
rect 15120 17066 15332 17070
rect 15108 17060 15332 17066
rect 15160 17054 15332 17060
rect 15108 17002 15160 17008
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 14924 16584 14976 16590
rect 15212 16538 15240 16934
rect 14976 16532 15240 16538
rect 14924 16526 15240 16532
rect 14936 16510 15240 16526
rect 15488 16504 15516 17614
rect 15568 16516 15620 16522
rect 15488 16476 15568 16504
rect 15488 16182 15516 16476
rect 15568 16458 15620 16464
rect 15476 16176 15528 16182
rect 15476 16118 15528 16124
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14108 15094 14136 15982
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13554 13084 13862 13093
rect 13554 13082 13560 13084
rect 13616 13082 13640 13084
rect 13696 13082 13720 13084
rect 13776 13082 13800 13084
rect 13856 13082 13862 13084
rect 13616 13030 13618 13082
rect 13798 13030 13800 13082
rect 13554 13028 13560 13030
rect 13616 13028 13640 13030
rect 13696 13028 13720 13030
rect 13776 13028 13800 13030
rect 13856 13028 13862 13030
rect 13554 13019 13862 13028
rect 13924 12986 13952 13466
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13910 12880 13966 12889
rect 13910 12815 13966 12824
rect 13924 12782 13952 12815
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13832 12306 13860 12582
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13554 11996 13862 12005
rect 13554 11994 13560 11996
rect 13616 11994 13640 11996
rect 13696 11994 13720 11996
rect 13776 11994 13800 11996
rect 13856 11994 13862 11996
rect 13616 11942 13618 11994
rect 13798 11942 13800 11994
rect 13554 11940 13560 11942
rect 13616 11940 13640 11942
rect 13696 11940 13720 11942
rect 13776 11940 13800 11942
rect 13856 11940 13862 11942
rect 13554 11931 13862 11940
rect 13820 11824 13872 11830
rect 13634 11792 13690 11801
rect 13820 11766 13872 11772
rect 13634 11727 13636 11736
rect 13688 11727 13690 11736
rect 13636 11698 13688 11704
rect 13832 11558 13860 11766
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13554 10908 13862 10917
rect 13554 10906 13560 10908
rect 13616 10906 13640 10908
rect 13696 10906 13720 10908
rect 13776 10906 13800 10908
rect 13856 10906 13862 10908
rect 13616 10854 13618 10906
rect 13798 10854 13800 10906
rect 13554 10852 13560 10854
rect 13616 10852 13640 10854
rect 13696 10852 13720 10854
rect 13776 10852 13800 10854
rect 13856 10852 13862 10854
rect 13554 10843 13862 10852
rect 13554 9820 13862 9829
rect 13554 9818 13560 9820
rect 13616 9818 13640 9820
rect 13696 9818 13720 9820
rect 13776 9818 13800 9820
rect 13856 9818 13862 9820
rect 13616 9766 13618 9818
rect 13798 9766 13800 9818
rect 13554 9764 13560 9766
rect 13616 9764 13640 9766
rect 13696 9764 13720 9766
rect 13776 9764 13800 9766
rect 13856 9764 13862 9766
rect 13554 9755 13862 9764
rect 13728 9376 13780 9382
rect 13924 9364 13952 12174
rect 14016 11898 14044 14758
rect 14108 14414 14136 15030
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14200 14074 14228 15438
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14384 14482 14412 15302
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 15488 14414 15516 16118
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14476 14074 14504 14214
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14292 13326 14320 13874
rect 14476 13546 14504 14010
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 14384 13518 14504 13546
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 14108 12850 14136 13194
rect 14186 12880 14242 12889
rect 14096 12844 14148 12850
rect 14186 12815 14242 12824
rect 14096 12786 14148 12792
rect 14108 12374 14136 12786
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14004 11892 14056 11898
rect 14004 11834 14056 11840
rect 14108 11762 14136 12310
rect 14200 11898 14228 12815
rect 14292 12646 14320 13262
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 13780 9336 13952 9364
rect 13728 9318 13780 9324
rect 13554 8732 13862 8741
rect 13554 8730 13560 8732
rect 13616 8730 13640 8732
rect 13696 8730 13720 8732
rect 13776 8730 13800 8732
rect 13856 8730 13862 8732
rect 13616 8678 13618 8730
rect 13798 8678 13800 8730
rect 13554 8676 13560 8678
rect 13616 8676 13640 8678
rect 13696 8676 13720 8678
rect 13776 8676 13800 8678
rect 13856 8676 13862 8678
rect 13554 8667 13862 8676
rect 13924 8634 13952 9336
rect 14016 9110 14044 9862
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14004 9104 14056 9110
rect 14004 9046 14056 9052
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13832 8022 13860 8434
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 13554 7644 13862 7653
rect 13554 7642 13560 7644
rect 13616 7642 13640 7644
rect 13696 7642 13720 7644
rect 13776 7642 13800 7644
rect 13856 7642 13862 7644
rect 13616 7590 13618 7642
rect 13798 7590 13800 7642
rect 13554 7588 13560 7590
rect 13616 7588 13640 7590
rect 13696 7588 13720 7590
rect 13776 7588 13800 7590
rect 13856 7588 13862 7590
rect 13554 7579 13862 7588
rect 13924 7002 13952 7890
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14016 7410 14044 7686
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 13912 6996 13964 7002
rect 13912 6938 13964 6944
rect 14016 6798 14044 7142
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 13554 6556 13862 6565
rect 13554 6554 13560 6556
rect 13616 6554 13640 6556
rect 13696 6554 13720 6556
rect 13776 6554 13800 6556
rect 13856 6554 13862 6556
rect 13616 6502 13618 6554
rect 13798 6502 13800 6554
rect 13554 6500 13560 6502
rect 13616 6500 13640 6502
rect 13696 6500 13720 6502
rect 13776 6500 13800 6502
rect 13856 6500 13862 6502
rect 13554 6491 13862 6500
rect 14016 6458 14044 6734
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 13554 5468 13862 5477
rect 13554 5466 13560 5468
rect 13616 5466 13640 5468
rect 13696 5466 13720 5468
rect 13776 5466 13800 5468
rect 13856 5466 13862 5468
rect 13616 5414 13618 5466
rect 13798 5414 13800 5466
rect 13554 5412 13560 5414
rect 13616 5412 13640 5414
rect 13696 5412 13720 5414
rect 13776 5412 13800 5414
rect 13856 5412 13862 5414
rect 13554 5403 13862 5412
rect 13924 4826 13952 6122
rect 14016 5914 14044 6258
rect 14108 6118 14136 9522
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14016 4826 14044 5850
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 13556 4690 13584 4762
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13554 4380 13862 4389
rect 13554 4378 13560 4380
rect 13616 4378 13640 4380
rect 13696 4378 13720 4380
rect 13776 4378 13800 4380
rect 13856 4378 13862 4380
rect 13616 4326 13618 4378
rect 13798 4326 13800 4378
rect 13554 4324 13560 4326
rect 13616 4324 13640 4326
rect 13696 4324 13720 4326
rect 13776 4324 13800 4326
rect 13856 4324 13862 4326
rect 13554 4315 13862 4324
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12360 3194 12388 3402
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12452 3126 12480 3674
rect 13280 3194 13308 3878
rect 13464 3738 13492 4082
rect 13648 3738 13676 4218
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13554 3292 13862 3301
rect 13554 3290 13560 3292
rect 13616 3290 13640 3292
rect 13696 3290 13720 3292
rect 13776 3290 13800 3292
rect 13856 3290 13862 3292
rect 13616 3238 13618 3290
rect 13798 3238 13800 3290
rect 13554 3236 13560 3238
rect 13616 3236 13640 3238
rect 13696 3236 13720 3238
rect 13776 3236 13800 3238
rect 13856 3236 13862 3238
rect 13554 3227 13862 3236
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 10403 2748 10711 2757
rect 10403 2746 10409 2748
rect 10465 2746 10489 2748
rect 10545 2746 10569 2748
rect 10625 2746 10649 2748
rect 10705 2746 10711 2748
rect 10465 2694 10467 2746
rect 10647 2694 10649 2746
rect 10403 2692 10409 2694
rect 10465 2692 10489 2694
rect 10545 2692 10569 2694
rect 10625 2692 10649 2694
rect 10705 2692 10711 2694
rect 10403 2683 10711 2692
rect 14200 2446 14228 11018
rect 14384 10130 14412 13518
rect 14740 13456 14792 13462
rect 14740 13398 14792 13404
rect 14464 13388 14516 13394
rect 14464 13330 14516 13336
rect 14476 12714 14504 13330
rect 14752 13190 14780 13398
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14464 12708 14516 12714
rect 14464 12650 14516 12656
rect 14462 12336 14518 12345
rect 14462 12271 14464 12280
rect 14516 12271 14518 12280
rect 14464 12242 14516 12248
rect 14568 12170 14596 12786
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14568 11694 14596 12106
rect 14752 11801 14780 13126
rect 14936 12986 14964 13194
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 15028 12889 15056 13670
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15120 12986 15148 13126
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15014 12880 15070 12889
rect 14924 12844 14976 12850
rect 15014 12815 15070 12824
rect 14924 12786 14976 12792
rect 14936 12238 14964 12786
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 14844 11830 14872 12174
rect 14936 12102 14964 12174
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 15028 11898 15056 12106
rect 15016 11892 15068 11898
rect 15304 11880 15332 12242
rect 15396 12170 15424 13262
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15580 12986 15608 13126
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15672 12918 15700 26930
rect 17040 26784 17092 26790
rect 17040 26726 17092 26732
rect 16705 26684 17013 26693
rect 16705 26682 16711 26684
rect 16767 26682 16791 26684
rect 16847 26682 16871 26684
rect 16927 26682 16951 26684
rect 17007 26682 17013 26684
rect 16767 26630 16769 26682
rect 16949 26630 16951 26682
rect 16705 26628 16711 26630
rect 16767 26628 16791 26630
rect 16847 26628 16871 26630
rect 16927 26628 16951 26630
rect 17007 26628 17013 26630
rect 16705 26619 17013 26628
rect 17052 25974 17080 26726
rect 17040 25968 17092 25974
rect 17040 25910 17092 25916
rect 16580 25832 16632 25838
rect 16580 25774 16632 25780
rect 16304 25356 16356 25362
rect 16304 25298 16356 25304
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 15752 24608 15804 24614
rect 15752 24550 15804 24556
rect 15764 16674 15792 24550
rect 15842 24304 15898 24313
rect 15842 24239 15844 24248
rect 15896 24239 15898 24248
rect 15844 24210 15896 24216
rect 15936 23520 15988 23526
rect 15936 23462 15988 23468
rect 15948 23050 15976 23462
rect 16040 23322 16068 24754
rect 16028 23316 16080 23322
rect 16316 23304 16344 25298
rect 16488 24608 16540 24614
rect 16488 24550 16540 24556
rect 16500 24410 16528 24550
rect 16488 24404 16540 24410
rect 16488 24346 16540 24352
rect 16028 23258 16080 23264
rect 16132 23276 16344 23304
rect 15936 23044 15988 23050
rect 15936 22986 15988 22992
rect 15844 22976 15896 22982
rect 15844 22918 15896 22924
rect 15856 22438 15884 22918
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 15844 20868 15896 20874
rect 15844 20810 15896 20816
rect 15856 20058 15884 20810
rect 15948 20534 15976 22986
rect 16028 22568 16080 22574
rect 16028 22510 16080 22516
rect 16040 21486 16068 22510
rect 16132 22234 16160 23276
rect 16212 23180 16264 23186
rect 16212 23122 16264 23128
rect 16120 22228 16172 22234
rect 16120 22170 16172 22176
rect 16224 22030 16252 23122
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16304 23044 16356 23050
rect 16304 22986 16356 22992
rect 16316 22778 16344 22986
rect 16408 22778 16436 23054
rect 16304 22772 16356 22778
rect 16304 22714 16356 22720
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 16316 22522 16344 22714
rect 16316 22494 16436 22522
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 16028 21480 16080 21486
rect 16028 21422 16080 21428
rect 15936 20528 15988 20534
rect 15936 20470 15988 20476
rect 16040 20482 16068 21422
rect 16132 21146 16160 21966
rect 16224 21690 16252 21966
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 16132 20602 16160 21082
rect 16120 20596 16172 20602
rect 16120 20538 16172 20544
rect 16316 20482 16344 22374
rect 16408 21146 16436 22494
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 16500 21622 16528 21830
rect 16488 21616 16540 21622
rect 16488 21558 16540 21564
rect 16592 21554 16620 25774
rect 16705 25596 17013 25605
rect 16705 25594 16711 25596
rect 16767 25594 16791 25596
rect 16847 25594 16871 25596
rect 16927 25594 16951 25596
rect 17007 25594 17013 25596
rect 16767 25542 16769 25594
rect 16949 25542 16951 25594
rect 16705 25540 16711 25542
rect 16767 25540 16791 25542
rect 16847 25540 16871 25542
rect 16927 25540 16951 25542
rect 17007 25540 17013 25542
rect 16705 25531 17013 25540
rect 17144 25498 17172 26930
rect 20720 26920 20772 26926
rect 20720 26862 20772 26868
rect 19616 26784 19668 26790
rect 19616 26726 19668 26732
rect 17316 26376 17368 26382
rect 17316 26318 17368 26324
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 17684 26376 17736 26382
rect 17684 26318 17736 26324
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 17132 25492 17184 25498
rect 17132 25434 17184 25440
rect 17328 25294 17356 26318
rect 17408 26240 17460 26246
rect 17408 26182 17460 26188
rect 17420 25294 17448 26182
rect 17512 25498 17540 26318
rect 17696 25702 17724 26318
rect 18236 25968 18288 25974
rect 18236 25910 18288 25916
rect 17684 25696 17736 25702
rect 17684 25638 17736 25644
rect 17500 25492 17552 25498
rect 17500 25434 17552 25440
rect 17316 25288 17368 25294
rect 17316 25230 17368 25236
rect 17408 25288 17460 25294
rect 17408 25230 17460 25236
rect 16705 24508 17013 24517
rect 16705 24506 16711 24508
rect 16767 24506 16791 24508
rect 16847 24506 16871 24508
rect 16927 24506 16951 24508
rect 17007 24506 17013 24508
rect 16767 24454 16769 24506
rect 16949 24454 16951 24506
rect 16705 24452 16711 24454
rect 16767 24452 16791 24454
rect 16847 24452 16871 24454
rect 16927 24452 16951 24454
rect 17007 24452 17013 24454
rect 16705 24443 17013 24452
rect 17328 24070 17356 25230
rect 17696 25226 17724 25638
rect 17776 25356 17828 25362
rect 17776 25298 17828 25304
rect 17684 25220 17736 25226
rect 17684 25162 17736 25168
rect 17500 24880 17552 24886
rect 17500 24822 17552 24828
rect 17512 24410 17540 24822
rect 17500 24404 17552 24410
rect 17500 24346 17552 24352
rect 17316 24064 17368 24070
rect 17316 24006 17368 24012
rect 17328 23662 17356 24006
rect 17040 23656 17092 23662
rect 17040 23598 17092 23604
rect 17316 23656 17368 23662
rect 17316 23598 17368 23604
rect 16705 23420 17013 23429
rect 16705 23418 16711 23420
rect 16767 23418 16791 23420
rect 16847 23418 16871 23420
rect 16927 23418 16951 23420
rect 17007 23418 17013 23420
rect 16767 23366 16769 23418
rect 16949 23366 16951 23418
rect 16705 23364 16711 23366
rect 16767 23364 16791 23366
rect 16847 23364 16871 23366
rect 16927 23364 16951 23366
rect 17007 23364 17013 23366
rect 16705 23355 17013 23364
rect 17052 23322 17080 23598
rect 17040 23316 17092 23322
rect 17040 23258 17092 23264
rect 17328 23186 17356 23598
rect 17316 23180 17368 23186
rect 17316 23122 17368 23128
rect 17408 23180 17460 23186
rect 17408 23122 17460 23128
rect 16705 22332 17013 22341
rect 16705 22330 16711 22332
rect 16767 22330 16791 22332
rect 16847 22330 16871 22332
rect 16927 22330 16951 22332
rect 17007 22330 17013 22332
rect 16767 22278 16769 22330
rect 16949 22278 16951 22330
rect 16705 22276 16711 22278
rect 16767 22276 16791 22278
rect 16847 22276 16871 22278
rect 16927 22276 16951 22278
rect 17007 22276 17013 22278
rect 16705 22267 17013 22276
rect 17420 22094 17448 23122
rect 17788 23118 17816 25298
rect 18248 25242 18276 25910
rect 18432 25838 18460 26318
rect 18512 26308 18564 26314
rect 18512 26250 18564 26256
rect 18524 25974 18552 26250
rect 18512 25968 18564 25974
rect 18512 25910 18564 25916
rect 18420 25832 18472 25838
rect 18420 25774 18472 25780
rect 18432 25294 18460 25774
rect 19248 25696 19300 25702
rect 19248 25638 19300 25644
rect 19260 25294 19288 25638
rect 19628 25362 19656 26726
rect 19856 26140 20164 26149
rect 19856 26138 19862 26140
rect 19918 26138 19942 26140
rect 19998 26138 20022 26140
rect 20078 26138 20102 26140
rect 20158 26138 20164 26140
rect 19918 26086 19920 26138
rect 20100 26086 20102 26138
rect 19856 26084 19862 26086
rect 19918 26084 19942 26086
rect 19998 26084 20022 26086
rect 20078 26084 20102 26086
rect 20158 26084 20164 26086
rect 19856 26075 20164 26084
rect 20628 25832 20680 25838
rect 20628 25774 20680 25780
rect 20260 25696 20312 25702
rect 20260 25638 20312 25644
rect 19616 25356 19668 25362
rect 19616 25298 19668 25304
rect 18064 25214 18276 25242
rect 18328 25288 18380 25294
rect 18328 25230 18380 25236
rect 18420 25288 18472 25294
rect 18420 25230 18472 25236
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 18064 25158 18092 25214
rect 18052 25152 18104 25158
rect 18052 25094 18104 25100
rect 18144 25152 18196 25158
rect 18144 25094 18196 25100
rect 17868 24744 17920 24750
rect 17868 24686 17920 24692
rect 17880 24342 17908 24686
rect 17960 24608 18012 24614
rect 17960 24550 18012 24556
rect 17868 24336 17920 24342
rect 17868 24278 17920 24284
rect 17972 24206 18000 24550
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 17960 24200 18012 24206
rect 17960 24142 18012 24148
rect 17880 23712 17908 24142
rect 17972 23866 18000 24142
rect 17960 23860 18012 23866
rect 17960 23802 18012 23808
rect 17960 23724 18012 23730
rect 17880 23684 17960 23712
rect 17960 23666 18012 23672
rect 17776 23112 17828 23118
rect 17776 23054 17828 23060
rect 17868 22228 17920 22234
rect 17868 22170 17920 22176
rect 17328 22066 17448 22094
rect 17040 21888 17092 21894
rect 17040 21830 17092 21836
rect 16580 21548 16632 21554
rect 16580 21490 16632 21496
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 16396 21004 16448 21010
rect 16396 20946 16448 20952
rect 16488 21004 16540 21010
rect 16592 20992 16620 21490
rect 17052 21486 17080 21830
rect 17040 21480 17092 21486
rect 17040 21422 17092 21428
rect 16705 21244 17013 21253
rect 16705 21242 16711 21244
rect 16767 21242 16791 21244
rect 16847 21242 16871 21244
rect 16927 21242 16951 21244
rect 17007 21242 17013 21244
rect 16767 21190 16769 21242
rect 16949 21190 16951 21242
rect 16705 21188 16711 21190
rect 16767 21188 16791 21190
rect 16847 21188 16871 21190
rect 16927 21188 16951 21190
rect 17007 21188 17013 21190
rect 16705 21179 17013 21188
rect 16540 20964 16620 20992
rect 16488 20946 16540 20952
rect 16408 20534 16436 20946
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 15948 18630 15976 20470
rect 16040 20466 16160 20482
rect 16224 20466 16344 20482
rect 16396 20528 16448 20534
rect 16396 20470 16448 20476
rect 16040 20460 16172 20466
rect 16040 20454 16120 20460
rect 16120 20402 16172 20408
rect 16212 20460 16344 20466
rect 16264 20454 16344 20460
rect 16212 20402 16264 20408
rect 16224 18970 16252 20402
rect 16592 20262 16620 20964
rect 17052 20602 17080 21422
rect 17040 20596 17092 20602
rect 17040 20538 17092 20544
rect 17040 20392 17092 20398
rect 17328 20380 17356 22066
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17408 21888 17460 21894
rect 17408 21830 17460 21836
rect 17420 21010 17448 21830
rect 17408 21004 17460 21010
rect 17408 20946 17460 20952
rect 17512 20602 17540 21966
rect 17776 20936 17828 20942
rect 17776 20878 17828 20884
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17684 20460 17736 20466
rect 17684 20402 17736 20408
rect 17092 20352 17356 20380
rect 17040 20334 17092 20340
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 16210 18864 16266 18873
rect 16210 18799 16212 18808
rect 16264 18799 16266 18808
rect 16212 18770 16264 18776
rect 16118 18728 16174 18737
rect 16118 18663 16174 18672
rect 16132 18630 16160 18663
rect 15936 18624 15988 18630
rect 15936 18566 15988 18572
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 15948 18358 15976 18566
rect 16132 18426 16160 18566
rect 16120 18420 16172 18426
rect 16120 18362 16172 18368
rect 15936 18352 15988 18358
rect 15936 18294 15988 18300
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15856 17882 15884 18226
rect 15844 17876 15896 17882
rect 15844 17818 15896 17824
rect 16224 17746 16252 18770
rect 16316 18766 16344 19654
rect 16500 19514 16528 19790
rect 16592 19514 16620 20198
rect 16705 20156 17013 20165
rect 16705 20154 16711 20156
rect 16767 20154 16791 20156
rect 16847 20154 16871 20156
rect 16927 20154 16951 20156
rect 17007 20154 17013 20156
rect 16767 20102 16769 20154
rect 16949 20102 16951 20154
rect 16705 20100 16711 20102
rect 16767 20100 16791 20102
rect 16847 20100 16871 20102
rect 16927 20100 16951 20102
rect 17007 20100 17013 20102
rect 16705 20091 17013 20100
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16580 19508 16632 19514
rect 16580 19450 16632 19456
rect 16500 18766 16528 19450
rect 16948 19168 17000 19174
rect 17052 19156 17080 20334
rect 17316 19712 17368 19718
rect 17316 19654 17368 19660
rect 17328 19514 17356 19654
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 17000 19128 17080 19156
rect 16948 19110 17000 19116
rect 16705 19068 17013 19077
rect 16705 19066 16711 19068
rect 16767 19066 16791 19068
rect 16847 19066 16871 19068
rect 16927 19066 16951 19068
rect 17007 19066 17013 19068
rect 16767 19014 16769 19066
rect 16949 19014 16951 19066
rect 16705 19012 16711 19014
rect 16767 19012 16791 19014
rect 16847 19012 16871 19014
rect 16927 19012 16951 19014
rect 17007 19012 17013 19014
rect 16705 19003 17013 19012
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 17052 18714 17080 19128
rect 17144 18834 17172 19246
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 16580 18692 16632 18698
rect 16580 18634 16632 18640
rect 16672 18692 16724 18698
rect 17052 18686 17356 18714
rect 16672 18634 16724 18640
rect 16592 18170 16620 18634
rect 16684 18358 16712 18634
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 16672 18352 16724 18358
rect 16672 18294 16724 18300
rect 16500 18142 16620 18170
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 15764 16646 15884 16674
rect 15856 14074 15884 16646
rect 16224 15502 16252 17682
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16500 17490 16528 18142
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16592 17678 16620 18022
rect 16705 17980 17013 17989
rect 16705 17978 16711 17980
rect 16767 17978 16791 17980
rect 16847 17978 16871 17980
rect 16927 17978 16951 17980
rect 17007 17978 17013 17980
rect 16767 17926 16769 17978
rect 16949 17926 16951 17978
rect 16705 17924 16711 17926
rect 16767 17924 16791 17926
rect 16847 17924 16871 17926
rect 16927 17924 16951 17926
rect 17007 17924 17013 17926
rect 16705 17915 17013 17924
rect 17052 17678 17080 18566
rect 17328 17728 17356 18686
rect 17408 18692 17460 18698
rect 17408 18634 17460 18640
rect 17420 18426 17448 18634
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17498 17776 17554 17785
rect 17408 17740 17460 17746
rect 17328 17700 17408 17728
rect 17498 17711 17554 17720
rect 17408 17682 17460 17688
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 16408 17270 16436 17478
rect 16500 17462 16620 17490
rect 16396 17264 16448 17270
rect 16396 17206 16448 17212
rect 16408 16794 16436 17206
rect 16396 16788 16448 16794
rect 16396 16730 16448 16736
rect 16592 16114 16620 17462
rect 17040 17128 17092 17134
rect 17040 17070 17092 17076
rect 16705 16892 17013 16901
rect 16705 16890 16711 16892
rect 16767 16890 16791 16892
rect 16847 16890 16871 16892
rect 16927 16890 16951 16892
rect 17007 16890 17013 16892
rect 16767 16838 16769 16890
rect 16949 16838 16951 16890
rect 16705 16836 16711 16838
rect 16767 16836 16791 16838
rect 16847 16836 16871 16838
rect 16927 16836 16951 16838
rect 17007 16836 17013 16838
rect 16705 16827 17013 16836
rect 17052 16674 17080 17070
rect 17420 17066 17448 17682
rect 17512 17678 17540 17711
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17408 17060 17460 17066
rect 17408 17002 17460 17008
rect 16960 16646 17080 16674
rect 17420 16658 17448 17002
rect 17408 16652 17460 16658
rect 16960 16250 16988 16646
rect 17408 16594 17460 16600
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 17052 16250 17080 16526
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16705 15804 17013 15813
rect 16705 15802 16711 15804
rect 16767 15802 16791 15804
rect 16847 15802 16871 15804
rect 16927 15802 16951 15804
rect 17007 15802 17013 15804
rect 16767 15750 16769 15802
rect 16949 15750 16951 15802
rect 16705 15748 16711 15750
rect 16767 15748 16791 15750
rect 16847 15748 16871 15750
rect 16927 15748 16951 15750
rect 17007 15748 17013 15750
rect 16705 15739 17013 15748
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 17236 15366 17264 16186
rect 17512 16114 17540 17614
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 16764 15088 16816 15094
rect 16762 15056 16764 15065
rect 16816 15056 16818 15065
rect 16762 14991 16818 15000
rect 16705 14716 17013 14725
rect 16705 14714 16711 14716
rect 16767 14714 16791 14716
rect 16847 14714 16871 14716
rect 16927 14714 16951 14716
rect 17007 14714 17013 14716
rect 16767 14662 16769 14714
rect 16949 14662 16951 14714
rect 16705 14660 16711 14662
rect 16767 14660 16791 14662
rect 16847 14660 16871 14662
rect 16927 14660 16951 14662
rect 17007 14660 17013 14662
rect 16705 14651 17013 14660
rect 17328 14074 17356 15846
rect 17604 14822 17632 20402
rect 17696 20262 17724 20402
rect 17684 20256 17736 20262
rect 17684 20198 17736 20204
rect 17684 19712 17736 19718
rect 17684 19654 17736 19660
rect 17696 18816 17724 19654
rect 17788 19514 17816 20878
rect 17880 19922 17908 22170
rect 17972 21622 18000 23666
rect 18156 23526 18184 25094
rect 18248 24886 18276 25214
rect 18340 24970 18368 25230
rect 18972 25152 19024 25158
rect 18972 25094 19024 25100
rect 18340 24942 18460 24970
rect 18236 24880 18288 24886
rect 18236 24822 18288 24828
rect 18248 23798 18276 24822
rect 18432 24682 18460 24942
rect 18880 24812 18932 24818
rect 18880 24754 18932 24760
rect 18420 24676 18472 24682
rect 18420 24618 18472 24624
rect 18788 24608 18840 24614
rect 18788 24550 18840 24556
rect 18602 24304 18658 24313
rect 18602 24239 18604 24248
rect 18656 24239 18658 24248
rect 18604 24210 18656 24216
rect 18236 23792 18288 23798
rect 18236 23734 18288 23740
rect 18144 23520 18196 23526
rect 18144 23462 18196 23468
rect 18512 23520 18564 23526
rect 18512 23462 18564 23468
rect 18524 23118 18552 23462
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 18512 22092 18564 22098
rect 18616 22080 18644 24210
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18708 23322 18736 24142
rect 18696 23316 18748 23322
rect 18696 23258 18748 23264
rect 18800 23118 18828 24550
rect 18892 23526 18920 24754
rect 18984 23662 19012 25094
rect 19260 24750 19288 25230
rect 19856 25052 20164 25061
rect 19856 25050 19862 25052
rect 19918 25050 19942 25052
rect 19998 25050 20022 25052
rect 20078 25050 20102 25052
rect 20158 25050 20164 25052
rect 19918 24998 19920 25050
rect 20100 24998 20102 25050
rect 19856 24996 19862 24998
rect 19918 24996 19942 24998
rect 19998 24996 20022 24998
rect 20078 24996 20102 24998
rect 20158 24996 20164 24998
rect 19856 24987 20164 24996
rect 19248 24744 19300 24750
rect 19248 24686 19300 24692
rect 19708 24744 19760 24750
rect 19708 24686 19760 24692
rect 19156 24608 19208 24614
rect 19156 24550 19208 24556
rect 19168 23798 19196 24550
rect 19156 23792 19208 23798
rect 19156 23734 19208 23740
rect 18972 23656 19024 23662
rect 18972 23598 19024 23604
rect 18880 23520 18932 23526
rect 18880 23462 18932 23468
rect 19064 23520 19116 23526
rect 19064 23462 19116 23468
rect 18788 23112 18840 23118
rect 18788 23054 18840 23060
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18800 22778 18828 22918
rect 18788 22772 18840 22778
rect 18788 22714 18840 22720
rect 18564 22052 18644 22080
rect 18512 22034 18564 22040
rect 17960 21616 18012 21622
rect 17960 21558 18012 21564
rect 17972 21078 18000 21558
rect 17960 21072 18012 21078
rect 17960 21014 18012 21020
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 18052 20868 18104 20874
rect 18052 20810 18104 20816
rect 18064 20466 18092 20810
rect 18432 20534 18460 20878
rect 18420 20528 18472 20534
rect 18420 20470 18472 20476
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 18328 20392 18380 20398
rect 18328 20334 18380 20340
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17776 19508 17828 19514
rect 17776 19450 17828 19456
rect 17776 18828 17828 18834
rect 17696 18788 17776 18816
rect 17696 18737 17724 18788
rect 17776 18770 17828 18776
rect 17682 18728 17738 18737
rect 17682 18663 17738 18672
rect 17696 18222 17724 18663
rect 17776 18352 17828 18358
rect 17776 18294 17828 18300
rect 17684 18216 17736 18222
rect 17684 18158 17736 18164
rect 17788 16658 17816 18294
rect 17880 17134 17908 19858
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18156 18630 18184 19110
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 18064 17678 18092 18022
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 18156 17542 18184 18158
rect 18340 17882 18368 20334
rect 18420 19508 18472 19514
rect 18420 19450 18472 19456
rect 18432 18698 18460 19450
rect 18524 18902 18552 22034
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 18708 21350 18736 21966
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18708 20466 18736 21286
rect 18892 20466 18920 23462
rect 18972 21004 19024 21010
rect 18972 20946 19024 20952
rect 18984 20466 19012 20946
rect 19076 20466 19104 23462
rect 19260 23118 19288 24686
rect 19340 24064 19392 24070
rect 19340 24006 19392 24012
rect 19352 23730 19380 24006
rect 19720 23866 19748 24686
rect 19856 23964 20164 23973
rect 19856 23962 19862 23964
rect 19918 23962 19942 23964
rect 19998 23962 20022 23964
rect 20078 23962 20102 23964
rect 20158 23962 20164 23964
rect 19918 23910 19920 23962
rect 20100 23910 20102 23962
rect 19856 23908 19862 23910
rect 19918 23908 19942 23910
rect 19998 23908 20022 23910
rect 20078 23908 20102 23910
rect 20158 23908 20164 23910
rect 19856 23899 20164 23908
rect 19708 23860 19760 23866
rect 19708 23802 19760 23808
rect 19340 23724 19392 23730
rect 19340 23666 19392 23672
rect 19892 23520 19944 23526
rect 19720 23480 19892 23508
rect 19248 23112 19300 23118
rect 19248 23054 19300 23060
rect 19260 22710 19288 23054
rect 19248 22704 19300 22710
rect 19248 22646 19300 22652
rect 19260 22098 19288 22646
rect 19248 22092 19300 22098
rect 19248 22034 19300 22040
rect 19260 21554 19288 22034
rect 19340 21956 19392 21962
rect 19340 21898 19392 21904
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19352 20602 19380 21898
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 19064 20460 19116 20466
rect 19064 20402 19116 20408
rect 19076 20346 19104 20402
rect 18708 20318 19104 20346
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18512 18896 18564 18902
rect 18512 18838 18564 18844
rect 18420 18692 18472 18698
rect 18420 18634 18472 18640
rect 18432 18290 18460 18634
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17776 16652 17828 16658
rect 17776 16594 17828 16600
rect 17880 16182 17908 17070
rect 17868 16176 17920 16182
rect 17868 16118 17920 16124
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 17684 15428 17736 15434
rect 17684 15370 17736 15376
rect 17696 14890 17724 15370
rect 17788 15094 17816 15506
rect 17868 15428 17920 15434
rect 17868 15370 17920 15376
rect 17776 15088 17828 15094
rect 17776 15030 17828 15036
rect 17684 14884 17736 14890
rect 17684 14826 17736 14832
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 16316 13394 16344 13670
rect 16705 13628 17013 13637
rect 16705 13626 16711 13628
rect 16767 13626 16791 13628
rect 16847 13626 16871 13628
rect 16927 13626 16951 13628
rect 17007 13626 17013 13628
rect 16767 13574 16769 13626
rect 16949 13574 16951 13626
rect 16705 13572 16711 13574
rect 16767 13572 16791 13574
rect 16847 13572 16871 13574
rect 16927 13572 16951 13574
rect 17007 13572 17013 13574
rect 16705 13563 17013 13572
rect 17052 13530 17080 13874
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15384 12164 15436 12170
rect 15384 12106 15436 12112
rect 15384 11892 15436 11898
rect 15304 11852 15384 11880
rect 15016 11834 15068 11840
rect 15384 11834 15436 11840
rect 14832 11824 14884 11830
rect 14738 11792 14794 11801
rect 14648 11756 14700 11762
rect 14832 11766 14884 11772
rect 15488 11762 15516 12786
rect 15658 12336 15714 12345
rect 15658 12271 15660 12280
rect 15712 12271 15714 12280
rect 15660 12242 15712 12248
rect 15764 12102 15792 12854
rect 15934 12744 15990 12753
rect 15934 12679 15936 12688
rect 15988 12679 15990 12688
rect 15936 12650 15988 12656
rect 16040 12434 16068 13262
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16316 12434 16344 12582
rect 16040 12406 16344 12434
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15580 11801 15608 12038
rect 15566 11792 15622 11801
rect 14738 11727 14794 11736
rect 15016 11756 15068 11762
rect 14648 11698 14700 11704
rect 15384 11756 15436 11762
rect 15068 11716 15384 11744
rect 15016 11698 15068 11704
rect 15384 11698 15436 11704
rect 15476 11756 15528 11762
rect 15566 11727 15622 11736
rect 15476 11698 15528 11704
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14464 11144 14516 11150
rect 14568 11132 14596 11630
rect 14660 11218 14688 11698
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 15764 11150 15792 12038
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 14516 11104 14596 11132
rect 15752 11144 15804 11150
rect 14464 11086 14516 11092
rect 15752 11086 15804 11092
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15672 10130 15700 10406
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 14384 9722 14412 10066
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14660 9518 14688 9862
rect 14936 9722 14964 9998
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 14924 9716 14976 9722
rect 14924 9658 14976 9664
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14660 9110 14688 9454
rect 15120 9178 15148 9522
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 14648 9104 14700 9110
rect 14648 9046 14700 9052
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 7954 14596 8230
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14476 7546 14504 7822
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14660 7426 14688 9046
rect 15212 9042 15240 9522
rect 15304 9042 15332 9862
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14752 8362 14780 8570
rect 15028 8566 15056 8774
rect 15212 8634 15240 8978
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15016 8560 15068 8566
rect 15016 8502 15068 8508
rect 14740 8356 14792 8362
rect 14740 8298 14792 8304
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14476 7398 14688 7426
rect 14384 6934 14412 7346
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14476 6254 14504 7398
rect 15028 7206 15056 8502
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15120 6866 15148 7482
rect 15672 7410 15700 7822
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14660 6322 14688 6666
rect 15304 6322 15332 7142
rect 15672 6866 15700 7346
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 14292 5302 14320 6054
rect 15580 5914 15608 6054
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 14280 5296 14332 5302
rect 14280 5238 14332 5244
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14384 3058 14412 3470
rect 15028 3194 15056 3878
rect 15212 3738 15240 4422
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15200 3460 15252 3466
rect 15252 3420 15332 3448
rect 15200 3402 15252 3408
rect 15016 3188 15068 3194
rect 15016 3130 15068 3136
rect 15304 3126 15332 3420
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 15856 2774 15884 11494
rect 16040 10470 16068 12406
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16040 9586 16068 10406
rect 16132 10266 16160 10406
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 16040 9042 16068 9522
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 16040 7886 16068 8366
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15948 5914 15976 6598
rect 16120 6384 16172 6390
rect 16120 6326 16172 6332
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15948 4486 15976 5646
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 15948 3738 15976 4422
rect 16040 4078 16068 4626
rect 16132 4214 16160 6326
rect 16120 4208 16172 4214
rect 16120 4150 16172 4156
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 16132 3194 16160 4150
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 16316 2774 16344 11834
rect 16408 11694 16436 12786
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 16705 12540 17013 12549
rect 16705 12538 16711 12540
rect 16767 12538 16791 12540
rect 16847 12538 16871 12540
rect 16927 12538 16951 12540
rect 17007 12538 17013 12540
rect 16767 12486 16769 12538
rect 16949 12486 16951 12538
rect 16705 12484 16711 12486
rect 16767 12484 16791 12486
rect 16847 12484 16871 12486
rect 16927 12484 16951 12486
rect 17007 12484 17013 12486
rect 16705 12475 17013 12484
rect 17236 12442 17264 12718
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 16705 11452 17013 11461
rect 16705 11450 16711 11452
rect 16767 11450 16791 11452
rect 16847 11450 16871 11452
rect 16927 11450 16951 11452
rect 17007 11450 17013 11452
rect 16767 11398 16769 11450
rect 16949 11398 16951 11450
rect 16705 11396 16711 11398
rect 16767 11396 16791 11398
rect 16847 11396 16871 11398
rect 16927 11396 16951 11398
rect 17007 11396 17013 11398
rect 16705 11387 17013 11396
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 16705 10364 17013 10373
rect 16705 10362 16711 10364
rect 16767 10362 16791 10364
rect 16847 10362 16871 10364
rect 16927 10362 16951 10364
rect 17007 10362 17013 10364
rect 16767 10310 16769 10362
rect 16949 10310 16951 10362
rect 16705 10308 16711 10310
rect 16767 10308 16791 10310
rect 16847 10308 16871 10310
rect 16927 10308 16951 10310
rect 17007 10308 17013 10310
rect 16705 10299 17013 10308
rect 17052 9654 17080 10950
rect 17236 10062 17264 11698
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17328 10810 17356 10950
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17420 10690 17448 11154
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17512 10810 17540 11086
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17328 10662 17448 10690
rect 17224 10056 17276 10062
rect 17144 10004 17224 10010
rect 17144 9998 17276 10004
rect 17144 9982 17264 9998
rect 17144 9722 17172 9982
rect 17328 9926 17356 10662
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17236 9722 17264 9862
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16408 9110 16436 9318
rect 16705 9276 17013 9285
rect 16705 9274 16711 9276
rect 16767 9274 16791 9276
rect 16847 9274 16871 9276
rect 16927 9274 16951 9276
rect 17007 9274 17013 9276
rect 16767 9222 16769 9274
rect 16949 9222 16951 9274
rect 16705 9220 16711 9222
rect 16767 9220 16791 9222
rect 16847 9220 16871 9222
rect 16927 9220 16951 9222
rect 17007 9220 17013 9222
rect 16705 9211 17013 9220
rect 16396 9104 16448 9110
rect 16396 9046 16448 9052
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16500 7886 16528 8570
rect 16592 8498 16620 8774
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16488 7880 16540 7886
rect 16488 7822 16540 7828
rect 16500 7546 16528 7822
rect 16592 7818 16620 8434
rect 16705 8188 17013 8197
rect 16705 8186 16711 8188
rect 16767 8186 16791 8188
rect 16847 8186 16871 8188
rect 16927 8186 16951 8188
rect 17007 8186 17013 8188
rect 16767 8134 16769 8186
rect 16949 8134 16951 8186
rect 16705 8132 16711 8134
rect 16767 8132 16791 8134
rect 16847 8132 16871 8134
rect 16927 8132 16951 8134
rect 17007 8132 17013 8134
rect 16705 8123 17013 8132
rect 17052 7954 17080 8910
rect 17144 8906 17172 9658
rect 17132 8900 17184 8906
rect 17132 8842 17184 8848
rect 17144 8430 17172 8842
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17236 8634 17264 8774
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 16580 7812 16632 7818
rect 16580 7754 16632 7760
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 16592 7426 16620 7754
rect 16500 7398 16620 7426
rect 16500 7274 16528 7398
rect 17144 7392 17172 8366
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 17236 7818 17264 8230
rect 17224 7812 17276 7818
rect 17224 7754 17276 7760
rect 17328 7410 17356 9862
rect 17604 9518 17632 14758
rect 17880 13802 17908 15370
rect 17972 15042 18000 17478
rect 18524 17338 18552 18838
rect 18512 17332 18564 17338
rect 18512 17274 18564 17280
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18524 16794 18552 17138
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18432 16114 18460 16594
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18328 15904 18380 15910
rect 18328 15846 18380 15852
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 17972 15014 18092 15042
rect 17868 13796 17920 13802
rect 17696 13756 17868 13784
rect 17696 12306 17724 13756
rect 17868 13738 17920 13744
rect 17776 13524 17828 13530
rect 17828 13484 17908 13512
rect 17776 13466 17828 13472
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17696 10538 17724 12242
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 17684 10532 17736 10538
rect 17684 10474 17736 10480
rect 17788 10418 17816 10610
rect 17696 10390 17816 10418
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17604 8906 17632 9454
rect 17696 9382 17724 10390
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17696 9042 17724 9318
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17592 8900 17644 8906
rect 17592 8842 17644 8848
rect 17604 8566 17632 8842
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17592 7812 17644 7818
rect 17592 7754 17644 7760
rect 17604 7478 17632 7754
rect 17880 7562 17908 13484
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17972 12102 18000 13262
rect 18064 12306 18092 15014
rect 18156 14958 18184 15642
rect 18340 15366 18368 15846
rect 18432 15570 18460 16050
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 18524 15502 18552 16594
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 18236 15360 18288 15366
rect 18236 15302 18288 15308
rect 18328 15360 18380 15366
rect 18328 15302 18380 15308
rect 18248 15094 18276 15302
rect 18236 15088 18288 15094
rect 18236 15030 18288 15036
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18156 14618 18184 14894
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18248 14482 18276 15030
rect 18236 14476 18288 14482
rect 18236 14418 18288 14424
rect 18340 14006 18368 15302
rect 18328 14000 18380 14006
rect 18328 13942 18380 13948
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18524 12918 18552 13330
rect 18616 13326 18644 19994
rect 18708 17785 18736 20318
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18800 19174 18828 19790
rect 18880 19304 18932 19310
rect 18880 19246 18932 19252
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18892 18630 18920 19246
rect 18880 18624 18932 18630
rect 18880 18566 18932 18572
rect 18892 17814 18920 18566
rect 18880 17808 18932 17814
rect 18694 17776 18750 17785
rect 18880 17750 18932 17756
rect 18694 17711 18750 17720
rect 18708 15910 18736 17711
rect 18788 17264 18840 17270
rect 18788 17206 18840 17212
rect 18800 16590 18828 17206
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18800 16046 18828 16526
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18892 16114 18920 16390
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18708 15502 18736 15846
rect 18892 15502 18920 16050
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18892 14550 18920 15438
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18512 12912 18564 12918
rect 18248 12860 18512 12866
rect 18248 12854 18564 12860
rect 18248 12838 18552 12854
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17972 9178 18000 12038
rect 18248 11830 18276 12838
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18432 11762 18460 12582
rect 18800 12238 18828 12582
rect 18984 12434 19012 20198
rect 19616 19168 19668 19174
rect 19616 19110 19668 19116
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19248 18624 19300 18630
rect 19248 18566 19300 18572
rect 19260 18426 19288 18566
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19064 17196 19116 17202
rect 19064 17138 19116 17144
rect 19076 15706 19104 17138
rect 19352 16794 19380 18906
rect 19628 18766 19656 19110
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19524 18216 19576 18222
rect 19524 18158 19576 18164
rect 19536 17882 19564 18158
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19720 17218 19748 23480
rect 19892 23462 19944 23468
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 20088 23322 20116 23462
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 20272 23186 20300 25638
rect 20640 24614 20668 25774
rect 20732 25362 20760 26862
rect 20904 26444 20956 26450
rect 20904 26386 20956 26392
rect 20812 25900 20864 25906
rect 20812 25842 20864 25848
rect 20720 25356 20772 25362
rect 20720 25298 20772 25304
rect 20732 24886 20760 25298
rect 20720 24880 20772 24886
rect 20720 24822 20772 24828
rect 20628 24608 20680 24614
rect 20628 24550 20680 24556
rect 20640 24070 20668 24550
rect 20824 24410 20852 25842
rect 20916 25838 20944 26386
rect 20904 25832 20956 25838
rect 20904 25774 20956 25780
rect 20916 25362 20944 25774
rect 20904 25356 20956 25362
rect 20904 25298 20956 25304
rect 20916 24954 20944 25298
rect 20904 24948 20956 24954
rect 20904 24890 20956 24896
rect 20812 24404 20864 24410
rect 20812 24346 20864 24352
rect 20352 24064 20404 24070
rect 20352 24006 20404 24012
rect 20628 24064 20680 24070
rect 20628 24006 20680 24012
rect 20364 23730 20392 24006
rect 20352 23724 20404 23730
rect 20352 23666 20404 23672
rect 20640 23254 20668 24006
rect 20812 23724 20864 23730
rect 20812 23666 20864 23672
rect 20628 23248 20680 23254
rect 20628 23190 20680 23196
rect 20260 23180 20312 23186
rect 20260 23122 20312 23128
rect 19856 22876 20164 22885
rect 19856 22874 19862 22876
rect 19918 22874 19942 22876
rect 19998 22874 20022 22876
rect 20078 22874 20102 22876
rect 20158 22874 20164 22876
rect 19918 22822 19920 22874
rect 20100 22822 20102 22874
rect 19856 22820 19862 22822
rect 19918 22820 19942 22822
rect 19998 22820 20022 22822
rect 20078 22820 20102 22822
rect 20158 22820 20164 22822
rect 19856 22811 20164 22820
rect 19856 21788 20164 21797
rect 19856 21786 19862 21788
rect 19918 21786 19942 21788
rect 19998 21786 20022 21788
rect 20078 21786 20102 21788
rect 20158 21786 20164 21788
rect 19918 21734 19920 21786
rect 20100 21734 20102 21786
rect 19856 21732 19862 21734
rect 19918 21732 19942 21734
rect 19998 21732 20022 21734
rect 20078 21732 20102 21734
rect 20158 21732 20164 21734
rect 19856 21723 20164 21732
rect 19856 20700 20164 20709
rect 19856 20698 19862 20700
rect 19918 20698 19942 20700
rect 19998 20698 20022 20700
rect 20078 20698 20102 20700
rect 20158 20698 20164 20700
rect 19918 20646 19920 20698
rect 20100 20646 20102 20698
rect 19856 20644 19862 20646
rect 19918 20644 19942 20646
rect 19998 20644 20022 20646
rect 20078 20644 20102 20646
rect 20158 20644 20164 20646
rect 19856 20635 20164 20644
rect 20272 20466 20300 23122
rect 20824 22778 20852 23666
rect 21008 23050 21036 26930
rect 22468 26784 22520 26790
rect 22468 26726 22520 26732
rect 22100 26308 22152 26314
rect 22100 26250 22152 26256
rect 21180 25696 21232 25702
rect 21180 25638 21232 25644
rect 21456 25696 21508 25702
rect 21456 25638 21508 25644
rect 21192 24274 21220 25638
rect 21468 25362 21496 25638
rect 22112 25498 22140 26250
rect 22480 25974 22508 26726
rect 23007 26684 23315 26693
rect 23007 26682 23013 26684
rect 23069 26682 23093 26684
rect 23149 26682 23173 26684
rect 23229 26682 23253 26684
rect 23309 26682 23315 26684
rect 23069 26630 23071 26682
rect 23251 26630 23253 26682
rect 23007 26628 23013 26630
rect 23069 26628 23093 26630
rect 23149 26628 23173 26630
rect 23229 26628 23253 26630
rect 23309 26628 23315 26630
rect 23007 26619 23315 26628
rect 22836 26444 22888 26450
rect 22836 26386 22888 26392
rect 22744 26240 22796 26246
rect 22744 26182 22796 26188
rect 22756 25974 22784 26182
rect 22468 25968 22520 25974
rect 22468 25910 22520 25916
rect 22744 25968 22796 25974
rect 22744 25910 22796 25916
rect 22100 25492 22152 25498
rect 22100 25434 22152 25440
rect 21456 25356 21508 25362
rect 21456 25298 21508 25304
rect 22560 25356 22612 25362
rect 22560 25298 22612 25304
rect 21364 25152 21416 25158
rect 21364 25094 21416 25100
rect 21272 24744 21324 24750
rect 21272 24686 21324 24692
rect 21284 24410 21312 24686
rect 21272 24404 21324 24410
rect 21272 24346 21324 24352
rect 21180 24268 21232 24274
rect 21180 24210 21232 24216
rect 21270 23760 21326 23769
rect 21376 23746 21404 25094
rect 21916 24812 21968 24818
rect 21916 24754 21968 24760
rect 21928 24721 21956 24754
rect 21914 24712 21970 24721
rect 21914 24647 21970 24656
rect 22100 24608 22152 24614
rect 22376 24608 22428 24614
rect 22100 24550 22152 24556
rect 22296 24568 22376 24596
rect 22008 24268 22060 24274
rect 22112 24256 22140 24550
rect 22060 24228 22140 24256
rect 22008 24210 22060 24216
rect 21732 24064 21784 24070
rect 21732 24006 21784 24012
rect 21744 23866 21772 24006
rect 21732 23860 21784 23866
rect 21732 23802 21784 23808
rect 21326 23718 21404 23746
rect 21270 23695 21326 23704
rect 20996 23044 21048 23050
rect 20996 22986 21048 22992
rect 21088 22976 21140 22982
rect 21088 22918 21140 22924
rect 20812 22772 20864 22778
rect 20812 22714 20864 22720
rect 20904 22432 20956 22438
rect 20904 22374 20956 22380
rect 20916 22094 20944 22374
rect 20732 22066 20944 22094
rect 20732 22030 20760 22066
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20352 21888 20404 21894
rect 20352 21830 20404 21836
rect 20364 21690 20392 21830
rect 20352 21684 20404 21690
rect 20352 21626 20404 21632
rect 20996 21616 21048 21622
rect 20996 21558 21048 21564
rect 20904 21480 20956 21486
rect 20904 21422 20956 21428
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 19856 19612 20164 19621
rect 19856 19610 19862 19612
rect 19918 19610 19942 19612
rect 19998 19610 20022 19612
rect 20078 19610 20102 19612
rect 20158 19610 20164 19612
rect 19918 19558 19920 19610
rect 20100 19558 20102 19610
rect 19856 19556 19862 19558
rect 19918 19556 19942 19558
rect 19998 19556 20022 19558
rect 20078 19556 20102 19558
rect 20158 19556 20164 19558
rect 19856 19547 20164 19556
rect 20732 19310 20760 19654
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20732 18834 20760 19110
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 19856 18524 20164 18533
rect 19856 18522 19862 18524
rect 19918 18522 19942 18524
rect 19998 18522 20022 18524
rect 20078 18522 20102 18524
rect 20158 18522 20164 18524
rect 19918 18470 19920 18522
rect 20100 18470 20102 18522
rect 19856 18468 19862 18470
rect 19918 18468 19942 18470
rect 19998 18468 20022 18470
rect 20078 18468 20102 18470
rect 20158 18468 20164 18470
rect 19856 18459 20164 18468
rect 20732 18222 20760 18770
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 19892 18080 19944 18086
rect 19892 18022 19944 18028
rect 19904 17678 19932 18022
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19856 17436 20164 17445
rect 19856 17434 19862 17436
rect 19918 17434 19942 17436
rect 19998 17434 20022 17436
rect 20078 17434 20102 17436
rect 20158 17434 20164 17436
rect 19918 17382 19920 17434
rect 20100 17382 20102 17434
rect 19856 17380 19862 17382
rect 19918 17380 19942 17382
rect 19998 17380 20022 17382
rect 20078 17380 20102 17382
rect 20158 17380 20164 17382
rect 19856 17371 20164 17380
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19536 17190 19748 17218
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19064 15700 19116 15706
rect 19064 15642 19116 15648
rect 19168 15434 19196 16050
rect 19352 15706 19380 16526
rect 19444 16182 19472 17138
rect 19432 16176 19484 16182
rect 19432 16118 19484 16124
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19444 15586 19472 16118
rect 19352 15558 19472 15586
rect 19352 15502 19380 15558
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19156 15428 19208 15434
rect 19156 15370 19208 15376
rect 19444 15366 19472 15438
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19156 15088 19208 15094
rect 19156 15030 19208 15036
rect 19168 14346 19196 15030
rect 19444 14550 19472 15302
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19156 14340 19208 14346
rect 19156 14282 19208 14288
rect 19168 14006 19196 14282
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19156 14000 19208 14006
rect 19156 13942 19208 13948
rect 19168 13394 19196 13942
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 18892 12406 19012 12434
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18432 11218 18460 11698
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 18708 11354 18736 11630
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 18892 10810 18920 12406
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18984 11150 19012 12038
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 19260 11082 19288 14214
rect 19536 12434 19564 17190
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19984 16992 20036 16998
rect 19984 16934 20036 16940
rect 19720 16522 19748 16934
rect 19996 16522 20024 16934
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19984 16516 20036 16522
rect 19984 16458 20036 16464
rect 19856 16348 20164 16357
rect 19856 16346 19862 16348
rect 19918 16346 19942 16348
rect 19998 16346 20022 16348
rect 20078 16346 20102 16348
rect 20158 16346 20164 16348
rect 19918 16294 19920 16346
rect 20100 16294 20102 16346
rect 19856 16292 19862 16294
rect 19918 16292 19942 16294
rect 19998 16292 20022 16294
rect 20078 16292 20102 16294
rect 20158 16292 20164 16294
rect 19856 16283 20164 16292
rect 20732 16182 20760 18158
rect 20812 17740 20864 17746
rect 20812 17682 20864 17688
rect 20824 16590 20852 17682
rect 20916 17610 20944 21422
rect 21008 21146 21036 21558
rect 20996 21140 21048 21146
rect 20996 21082 21048 21088
rect 21008 20890 21036 21082
rect 21100 21010 21128 22918
rect 21284 22642 21312 23695
rect 22020 23662 22048 24210
rect 22192 24200 22244 24206
rect 22192 24142 22244 24148
rect 22100 24132 22152 24138
rect 22100 24074 22152 24080
rect 22112 23730 22140 24074
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 22008 23656 22060 23662
rect 22008 23598 22060 23604
rect 21916 23520 21968 23526
rect 21916 23462 21968 23468
rect 21456 23044 21508 23050
rect 21456 22986 21508 22992
rect 21468 22778 21496 22986
rect 21456 22772 21508 22778
rect 21456 22714 21508 22720
rect 21272 22636 21324 22642
rect 21272 22578 21324 22584
rect 21284 21554 21312 22578
rect 21928 22030 21956 23462
rect 22020 23322 22048 23598
rect 22008 23316 22060 23322
rect 22008 23258 22060 23264
rect 22204 23118 22232 24142
rect 22192 23112 22244 23118
rect 22192 23054 22244 23060
rect 22192 22704 22244 22710
rect 22192 22646 22244 22652
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 21916 22024 21968 22030
rect 21546 21992 21602 22001
rect 21916 21966 21968 21972
rect 21546 21927 21548 21936
rect 21600 21927 21602 21936
rect 21548 21898 21600 21904
rect 21272 21548 21324 21554
rect 21272 21490 21324 21496
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 21008 20862 21128 20890
rect 21284 20874 21312 21490
rect 22112 21010 22140 22578
rect 22204 22234 22232 22646
rect 22192 22228 22244 22234
rect 22192 22170 22244 22176
rect 22100 21004 22152 21010
rect 22100 20946 22152 20952
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 20996 20800 21048 20806
rect 20996 20742 21048 20748
rect 21008 20262 21036 20742
rect 20996 20256 21048 20262
rect 20996 20198 21048 20204
rect 20996 18692 21048 18698
rect 20996 18634 21048 18640
rect 21008 18426 21036 18634
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 21100 18306 21128 20862
rect 21272 20868 21324 20874
rect 21272 20810 21324 20816
rect 21284 19378 21312 20810
rect 21468 20262 21496 20878
rect 22112 20534 22140 20946
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 21008 18278 21128 18306
rect 21376 18290 21404 20198
rect 22100 19848 22152 19854
rect 22100 19790 22152 19796
rect 22112 19514 22140 19790
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 21916 19372 21968 19378
rect 21916 19314 21968 19320
rect 21928 18612 21956 19314
rect 22008 19304 22060 19310
rect 22008 19246 22060 19252
rect 22020 18834 22048 19246
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22008 18828 22060 18834
rect 22008 18770 22060 18776
rect 22008 18624 22060 18630
rect 21928 18584 22008 18612
rect 21928 18290 21956 18584
rect 22008 18566 22060 18572
rect 22112 18358 22140 19110
rect 22100 18352 22152 18358
rect 22100 18294 22152 18300
rect 21364 18284 21416 18290
rect 20904 17604 20956 17610
rect 20904 17546 20956 17552
rect 20916 16658 20944 17546
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20720 16176 20772 16182
rect 20720 16118 20772 16124
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 19984 15972 20036 15978
rect 19984 15914 20036 15920
rect 19996 15638 20024 15914
rect 19984 15632 20036 15638
rect 19984 15574 20036 15580
rect 20456 15502 20484 15982
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20444 15496 20496 15502
rect 20444 15438 20496 15444
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19628 14618 19656 15302
rect 19856 15260 20164 15269
rect 19856 15258 19862 15260
rect 19918 15258 19942 15260
rect 19998 15258 20022 15260
rect 20078 15258 20102 15260
rect 20158 15258 20164 15260
rect 19918 15206 19920 15258
rect 20100 15206 20102 15258
rect 19856 15204 19862 15206
rect 19918 15204 19942 15206
rect 19998 15204 20022 15206
rect 20078 15204 20102 15206
rect 20158 15204 20164 15206
rect 19856 15195 20164 15204
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19720 14074 19748 14894
rect 20364 14482 20392 15438
rect 20456 15026 20484 15438
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 20352 14476 20404 14482
rect 20352 14418 20404 14424
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 19856 14172 20164 14181
rect 19856 14170 19862 14172
rect 19918 14170 19942 14172
rect 19998 14170 20022 14172
rect 20078 14170 20102 14172
rect 20158 14170 20164 14172
rect 19918 14118 19920 14170
rect 20100 14118 20102 14170
rect 19856 14116 19862 14118
rect 19918 14116 19942 14118
rect 19998 14116 20022 14118
rect 20078 14116 20102 14118
rect 20158 14116 20164 14118
rect 19856 14107 20164 14116
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 19856 13084 20164 13093
rect 19856 13082 19862 13084
rect 19918 13082 19942 13084
rect 19998 13082 20022 13084
rect 20078 13082 20102 13084
rect 20158 13082 20164 13084
rect 19918 13030 19920 13082
rect 20100 13030 20102 13082
rect 19856 13028 19862 13030
rect 19918 13028 19942 13030
rect 19998 13028 20022 13030
rect 20078 13028 20102 13030
rect 20158 13028 20164 13030
rect 19856 13019 20164 13028
rect 20272 12918 20300 14214
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 20352 12776 20404 12782
rect 20352 12718 20404 12724
rect 19352 12406 19564 12434
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19260 10810 19288 11018
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19156 10736 19208 10742
rect 19352 10690 19380 12406
rect 19524 11076 19576 11082
rect 19524 11018 19576 11024
rect 19536 10810 19564 11018
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19208 10684 19380 10690
rect 19156 10678 19380 10684
rect 19168 10662 19380 10678
rect 19522 10704 19578 10713
rect 19432 10668 19484 10674
rect 19522 10639 19524 10648
rect 19432 10610 19484 10616
rect 19576 10639 19578 10648
rect 19524 10610 19576 10616
rect 19444 10266 19472 10610
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 18432 9042 18460 10066
rect 19628 9518 19656 12718
rect 20364 12434 20392 12718
rect 20180 12406 20392 12434
rect 20180 12238 20208 12406
rect 20456 12322 20484 13806
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20272 12294 20484 12322
rect 20272 12238 20300 12294
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 19856 11996 20164 12005
rect 19856 11994 19862 11996
rect 19918 11994 19942 11996
rect 19998 11994 20022 11996
rect 20078 11994 20102 11996
rect 20158 11994 20164 11996
rect 19918 11942 19920 11994
rect 20100 11942 20102 11994
rect 19856 11940 19862 11942
rect 19918 11940 19942 11942
rect 19998 11940 20022 11942
rect 20078 11940 20102 11942
rect 20158 11940 20164 11942
rect 19856 11931 20164 11940
rect 19708 11008 19760 11014
rect 19708 10950 19760 10956
rect 19720 9654 19748 10950
rect 19856 10908 20164 10917
rect 19856 10906 19862 10908
rect 19918 10906 19942 10908
rect 19998 10906 20022 10908
rect 20078 10906 20102 10908
rect 20158 10906 20164 10908
rect 19918 10854 19920 10906
rect 20100 10854 20102 10906
rect 19856 10852 19862 10854
rect 19918 10852 19942 10854
rect 19998 10852 20022 10854
rect 20078 10852 20102 10854
rect 20158 10852 20164 10854
rect 19856 10843 20164 10852
rect 20272 10130 20300 12174
rect 20352 12164 20404 12170
rect 20352 12106 20404 12112
rect 20364 11558 20392 12106
rect 20548 11762 20576 12786
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20352 11552 20404 11558
rect 20352 11494 20404 11500
rect 20364 10674 20392 11494
rect 20640 10810 20668 16050
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20732 14890 20760 15370
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20824 14006 20852 16526
rect 20812 14000 20864 14006
rect 20812 13942 20864 13948
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20732 12170 20760 13126
rect 20916 12442 20944 16594
rect 21008 16522 21036 18278
rect 21364 18226 21416 18232
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21364 17196 21416 17202
rect 21364 17138 21416 17144
rect 21548 17196 21600 17202
rect 21548 17138 21600 17144
rect 20996 16516 21048 16522
rect 20996 16458 21048 16464
rect 21008 15026 21036 16458
rect 21376 16250 21404 17138
rect 21364 16244 21416 16250
rect 21364 16186 21416 16192
rect 21364 15904 21416 15910
rect 21364 15846 21416 15852
rect 21376 15026 21404 15846
rect 21560 15026 21588 17138
rect 21744 16046 21772 17614
rect 21824 16584 21876 16590
rect 21824 16526 21876 16532
rect 21836 16250 21864 16526
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21928 16130 21956 18226
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 22112 17678 22140 18022
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 22204 17542 22232 17818
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22100 16992 22152 16998
rect 22100 16934 22152 16940
rect 22112 16182 22140 16934
rect 21836 16102 21956 16130
rect 22100 16176 22152 16182
rect 22100 16118 22152 16124
rect 21732 16040 21784 16046
rect 21732 15982 21784 15988
rect 21744 15706 21772 15982
rect 21836 15978 21864 16102
rect 21824 15972 21876 15978
rect 21824 15914 21876 15920
rect 21732 15700 21784 15706
rect 21732 15642 21784 15648
rect 21836 15502 21864 15914
rect 22296 15570 22324 24568
rect 22376 24550 22428 24556
rect 22376 23724 22428 23730
rect 22376 23666 22428 23672
rect 22388 23322 22416 23666
rect 22572 23526 22600 25298
rect 22652 25220 22704 25226
rect 22652 25162 22704 25168
rect 22664 23866 22692 25162
rect 22756 24818 22784 25910
rect 22744 24812 22796 24818
rect 22744 24754 22796 24760
rect 22652 23860 22704 23866
rect 22652 23802 22704 23808
rect 22756 23769 22784 24754
rect 22742 23760 22798 23769
rect 22664 23730 22742 23746
rect 22652 23724 22742 23730
rect 22704 23718 22742 23724
rect 22742 23695 22798 23704
rect 22652 23666 22704 23672
rect 22744 23656 22796 23662
rect 22744 23598 22796 23604
rect 22652 23588 22704 23594
rect 22652 23530 22704 23536
rect 22560 23520 22612 23526
rect 22560 23462 22612 23468
rect 22376 23316 22428 23322
rect 22376 23258 22428 23264
rect 22560 23248 22612 23254
rect 22560 23190 22612 23196
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22480 22710 22508 22918
rect 22468 22704 22520 22710
rect 22468 22646 22520 22652
rect 22572 22438 22600 23190
rect 22560 22432 22612 22438
rect 22560 22374 22612 22380
rect 22376 22160 22428 22166
rect 22376 22102 22428 22108
rect 22388 17882 22416 22102
rect 22572 22098 22600 22374
rect 22560 22092 22612 22098
rect 22560 22034 22612 22040
rect 22560 21956 22612 21962
rect 22560 21898 22612 21904
rect 22572 21434 22600 21898
rect 22664 21554 22692 23530
rect 22756 23186 22784 23598
rect 22744 23180 22796 23186
rect 22744 23122 22796 23128
rect 22744 22976 22796 22982
rect 22744 22918 22796 22924
rect 22756 21962 22784 22918
rect 22848 22094 22876 26386
rect 26158 26140 26466 26149
rect 26158 26138 26164 26140
rect 26220 26138 26244 26140
rect 26300 26138 26324 26140
rect 26380 26138 26404 26140
rect 26460 26138 26466 26140
rect 26220 26086 26222 26138
rect 26402 26086 26404 26138
rect 26158 26084 26164 26086
rect 26220 26084 26244 26086
rect 26300 26084 26324 26086
rect 26380 26084 26404 26086
rect 26460 26084 26466 26086
rect 26158 26075 26466 26084
rect 23664 25696 23716 25702
rect 23664 25638 23716 25644
rect 23007 25596 23315 25605
rect 23007 25594 23013 25596
rect 23069 25594 23093 25596
rect 23149 25594 23173 25596
rect 23229 25594 23253 25596
rect 23309 25594 23315 25596
rect 23069 25542 23071 25594
rect 23251 25542 23253 25594
rect 23007 25540 23013 25542
rect 23069 25540 23093 25542
rect 23149 25540 23173 25542
rect 23229 25540 23253 25542
rect 23309 25540 23315 25542
rect 23007 25531 23315 25540
rect 23676 25498 23704 25638
rect 23664 25492 23716 25498
rect 23664 25434 23716 25440
rect 26332 25424 26384 25430
rect 26332 25366 26384 25372
rect 25688 25288 25740 25294
rect 26344 25265 26372 25366
rect 25688 25230 25740 25236
rect 26330 25256 26386 25265
rect 24400 25152 24452 25158
rect 24400 25094 24452 25100
rect 24412 24886 24440 25094
rect 24400 24880 24452 24886
rect 24400 24822 24452 24828
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23007 24508 23315 24517
rect 23007 24506 23013 24508
rect 23069 24506 23093 24508
rect 23149 24506 23173 24508
rect 23229 24506 23253 24508
rect 23309 24506 23315 24508
rect 23069 24454 23071 24506
rect 23251 24454 23253 24506
rect 23007 24452 23013 24454
rect 23069 24452 23093 24454
rect 23149 24452 23173 24454
rect 23229 24452 23253 24454
rect 23309 24452 23315 24454
rect 23007 24443 23315 24452
rect 22928 24200 22980 24206
rect 22928 24142 22980 24148
rect 22940 23322 22968 24142
rect 23400 23526 23428 24550
rect 23664 24064 23716 24070
rect 23664 24006 23716 24012
rect 23676 23866 23704 24006
rect 23664 23860 23716 23866
rect 23664 23802 23716 23808
rect 23388 23520 23440 23526
rect 23388 23462 23440 23468
rect 23007 23420 23315 23429
rect 23007 23418 23013 23420
rect 23069 23418 23093 23420
rect 23149 23418 23173 23420
rect 23229 23418 23253 23420
rect 23309 23418 23315 23420
rect 23069 23366 23071 23418
rect 23251 23366 23253 23418
rect 23007 23364 23013 23366
rect 23069 23364 23093 23366
rect 23149 23364 23173 23366
rect 23229 23364 23253 23366
rect 23309 23364 23315 23366
rect 23007 23355 23315 23364
rect 22928 23316 22980 23322
rect 22928 23258 22980 23264
rect 23400 22778 23428 23462
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 23007 22332 23315 22341
rect 23007 22330 23013 22332
rect 23069 22330 23093 22332
rect 23149 22330 23173 22332
rect 23229 22330 23253 22332
rect 23309 22330 23315 22332
rect 23069 22278 23071 22330
rect 23251 22278 23253 22330
rect 23007 22276 23013 22278
rect 23069 22276 23093 22278
rect 23149 22276 23173 22278
rect 23229 22276 23253 22278
rect 23309 22276 23315 22278
rect 23007 22267 23315 22276
rect 25700 22094 25728 25230
rect 26330 25191 26386 25200
rect 26158 25052 26466 25061
rect 26158 25050 26164 25052
rect 26220 25050 26244 25052
rect 26300 25050 26324 25052
rect 26380 25050 26404 25052
rect 26460 25050 26466 25052
rect 26220 24998 26222 25050
rect 26402 24998 26404 25050
rect 26158 24996 26164 24998
rect 26220 24996 26244 24998
rect 26300 24996 26324 24998
rect 26380 24996 26404 24998
rect 26460 24996 26466 24998
rect 26158 24987 26466 24996
rect 26158 23964 26466 23973
rect 26158 23962 26164 23964
rect 26220 23962 26244 23964
rect 26300 23962 26324 23964
rect 26380 23962 26404 23964
rect 26460 23962 26466 23964
rect 26220 23910 26222 23962
rect 26402 23910 26404 23962
rect 26158 23908 26164 23910
rect 26220 23908 26244 23910
rect 26300 23908 26324 23910
rect 26380 23908 26404 23910
rect 26460 23908 26466 23910
rect 26158 23899 26466 23908
rect 26158 22876 26466 22885
rect 26158 22874 26164 22876
rect 26220 22874 26244 22876
rect 26300 22874 26324 22876
rect 26380 22874 26404 22876
rect 26460 22874 26466 22876
rect 26220 22822 26222 22874
rect 26402 22822 26404 22874
rect 26158 22820 26164 22822
rect 26220 22820 26244 22822
rect 26300 22820 26324 22822
rect 26380 22820 26404 22822
rect 26460 22820 26466 22822
rect 26158 22811 26466 22820
rect 22848 22066 22968 22094
rect 22744 21956 22796 21962
rect 22744 21898 22796 21904
rect 22836 21888 22888 21894
rect 22836 21830 22888 21836
rect 22848 21690 22876 21830
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 22572 21406 22692 21434
rect 22664 20398 22692 21406
rect 22836 20460 22888 20466
rect 22836 20402 22888 20408
rect 22652 20392 22704 20398
rect 22652 20334 22704 20340
rect 22664 19922 22692 20334
rect 22652 19916 22704 19922
rect 22652 19858 22704 19864
rect 22664 18222 22692 19858
rect 22848 19446 22876 20402
rect 22940 19938 22968 22066
rect 25516 22066 25728 22094
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 23007 21244 23315 21253
rect 23007 21242 23013 21244
rect 23069 21242 23093 21244
rect 23149 21242 23173 21244
rect 23229 21242 23253 21244
rect 23309 21242 23315 21244
rect 23069 21190 23071 21242
rect 23251 21190 23253 21242
rect 23007 21188 23013 21190
rect 23069 21188 23093 21190
rect 23149 21188 23173 21190
rect 23229 21188 23253 21190
rect 23309 21188 23315 21190
rect 23007 21179 23315 21188
rect 23400 21146 23428 21490
rect 23388 21140 23440 21146
rect 23308 21100 23388 21128
rect 23308 20602 23336 21100
rect 23388 21082 23440 21088
rect 23296 20596 23348 20602
rect 23296 20538 23348 20544
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 23007 20156 23315 20165
rect 23007 20154 23013 20156
rect 23069 20154 23093 20156
rect 23149 20154 23173 20156
rect 23229 20154 23253 20156
rect 23309 20154 23315 20156
rect 23069 20102 23071 20154
rect 23251 20102 23253 20154
rect 23007 20100 23013 20102
rect 23069 20100 23093 20102
rect 23149 20100 23173 20102
rect 23229 20100 23253 20102
rect 23309 20100 23315 20102
rect 23007 20091 23315 20100
rect 23400 20058 23428 20470
rect 23848 20460 23900 20466
rect 23848 20402 23900 20408
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 24032 20460 24084 20466
rect 24032 20402 24084 20408
rect 25136 20460 25188 20466
rect 25136 20402 25188 20408
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 22940 19910 23060 19938
rect 23032 19854 23060 19910
rect 23020 19848 23072 19854
rect 23480 19848 23532 19854
rect 23020 19790 23072 19796
rect 23400 19796 23480 19802
rect 23400 19790 23532 19796
rect 22836 19440 22888 19446
rect 22836 19382 22888 19388
rect 23032 19378 23060 19790
rect 23400 19774 23520 19790
rect 22744 19372 22796 19378
rect 22744 19314 22796 19320
rect 23020 19372 23072 19378
rect 23020 19314 23072 19320
rect 22652 18216 22704 18222
rect 22652 18158 22704 18164
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22652 17876 22704 17882
rect 22652 17818 22704 17824
rect 22664 17678 22692 17818
rect 22468 17672 22520 17678
rect 22468 17614 22520 17620
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 22480 17338 22508 17614
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 21364 15020 21416 15026
rect 21364 14962 21416 14968
rect 21548 15020 21600 15026
rect 21548 14962 21600 14968
rect 21272 14952 21324 14958
rect 21272 14894 21324 14900
rect 21284 14464 21312 14894
rect 21456 14476 21508 14482
rect 21284 14436 21404 14464
rect 20996 12640 21048 12646
rect 20996 12582 21048 12588
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20720 12164 20772 12170
rect 20720 12106 20772 12112
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 20824 11150 20852 11630
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20916 11014 20944 11494
rect 20904 11008 20956 11014
rect 20904 10950 20956 10956
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 19856 9820 20164 9829
rect 19856 9818 19862 9820
rect 19918 9818 19942 9820
rect 19998 9818 20022 9820
rect 20078 9818 20102 9820
rect 20158 9818 20164 9820
rect 19918 9766 19920 9818
rect 20100 9766 20102 9818
rect 19856 9764 19862 9766
rect 19918 9764 19942 9766
rect 19998 9764 20022 9766
rect 20078 9764 20102 9766
rect 20158 9764 20164 9766
rect 19856 9755 20164 9764
rect 19708 9648 19760 9654
rect 19708 9590 19760 9596
rect 19616 9512 19668 9518
rect 19616 9454 19668 9460
rect 18972 9444 19024 9450
rect 18972 9386 19024 9392
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 17788 7534 17908 7562
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 17224 7404 17276 7410
rect 17144 7364 17224 7392
rect 17224 7346 17276 7352
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16488 7268 16540 7274
rect 16488 7210 16540 7216
rect 16592 6866 16620 7278
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 16705 7100 17013 7109
rect 16705 7098 16711 7100
rect 16767 7098 16791 7100
rect 16847 7098 16871 7100
rect 16927 7098 16951 7100
rect 17007 7098 17013 7100
rect 16767 7046 16769 7098
rect 16949 7046 16951 7098
rect 16705 7044 16711 7046
rect 16767 7044 16791 7046
rect 16847 7044 16871 7046
rect 16927 7044 16951 7046
rect 17007 7044 17013 7046
rect 16705 7035 17013 7044
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 16960 6458 16988 6598
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 17052 6322 17080 6598
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16592 5370 16620 6054
rect 16705 6012 17013 6021
rect 16705 6010 16711 6012
rect 16767 6010 16791 6012
rect 16847 6010 16871 6012
rect 16927 6010 16951 6012
rect 17007 6010 17013 6012
rect 16767 5958 16769 6010
rect 16949 5958 16951 6010
rect 16705 5956 16711 5958
rect 16767 5956 16791 5958
rect 16847 5956 16871 5958
rect 16927 5956 16951 5958
rect 17007 5956 17013 5958
rect 16705 5947 17013 5956
rect 17052 5778 17080 6258
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 17052 5234 17080 5714
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 16705 4924 17013 4933
rect 16705 4922 16711 4924
rect 16767 4922 16791 4924
rect 16847 4922 16871 4924
rect 16927 4922 16951 4924
rect 17007 4922 17013 4924
rect 16767 4870 16769 4922
rect 16949 4870 16951 4922
rect 16705 4868 16711 4870
rect 16767 4868 16791 4870
rect 16847 4868 16871 4870
rect 16927 4868 16951 4870
rect 17007 4868 17013 4870
rect 16705 4859 17013 4868
rect 16764 4752 16816 4758
rect 16764 4694 16816 4700
rect 16776 4486 16804 4694
rect 17052 4690 17080 4966
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 17144 4146 17172 7142
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16408 3194 16436 3878
rect 16705 3836 17013 3845
rect 16705 3834 16711 3836
rect 16767 3834 16791 3836
rect 16847 3834 16871 3836
rect 16927 3834 16951 3836
rect 17007 3834 17013 3836
rect 16767 3782 16769 3834
rect 16949 3782 16951 3834
rect 16705 3780 16711 3782
rect 16767 3780 16791 3782
rect 16847 3780 16871 3782
rect 16927 3780 16951 3782
rect 17007 3780 17013 3782
rect 16705 3771 17013 3780
rect 16580 3460 16632 3466
rect 16580 3402 16632 3408
rect 17040 3460 17092 3466
rect 17236 3448 17264 7346
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17420 6458 17448 6598
rect 17512 6458 17540 6802
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17592 5568 17644 5574
rect 17592 5510 17644 5516
rect 17604 5370 17632 5510
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17788 4554 17816 7534
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17972 6186 18000 6598
rect 18064 6390 18092 7686
rect 18340 7206 18368 8366
rect 18524 7954 18552 8978
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18616 8362 18644 8774
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18512 7948 18564 7954
rect 18512 7890 18564 7896
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 18052 6384 18104 6390
rect 18052 6326 18104 6332
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17880 5234 17908 5646
rect 17972 5574 18000 6122
rect 18064 5778 18092 6326
rect 18340 6322 18368 7142
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 18064 5658 18092 5714
rect 18064 5630 18184 5658
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 18156 5234 18184 5630
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 17776 4548 17828 4554
rect 17776 4490 17828 4496
rect 17788 4146 17816 4490
rect 17880 4146 17908 5170
rect 18156 5098 18184 5170
rect 18248 5098 18276 5510
rect 18340 5166 18368 6258
rect 18524 5778 18552 7890
rect 18616 7426 18644 8298
rect 18708 7546 18736 8774
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18616 7398 18736 7426
rect 18604 6656 18656 6662
rect 18604 6598 18656 6604
rect 18616 6254 18644 6598
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18708 5794 18736 7398
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18800 5914 18828 6734
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 18512 5772 18564 5778
rect 18708 5766 18828 5794
rect 18984 5778 19012 9386
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19260 9178 19288 9318
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 19076 6390 19104 8570
rect 19260 8430 19288 8910
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19352 7886 19380 8774
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19260 7546 19288 7686
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19064 6384 19116 6390
rect 19064 6326 19116 6332
rect 19536 5778 19564 6394
rect 19628 5778 19656 9318
rect 19720 8566 19748 9590
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 19856 8732 20164 8741
rect 19856 8730 19862 8732
rect 19918 8730 19942 8732
rect 19998 8730 20022 8732
rect 20078 8730 20102 8732
rect 20158 8730 20164 8732
rect 19918 8678 19920 8730
rect 20100 8678 20102 8730
rect 19856 8676 19862 8678
rect 19918 8676 19942 8678
rect 19998 8676 20022 8678
rect 20078 8676 20102 8678
rect 20158 8676 20164 8678
rect 19856 8667 20164 8676
rect 19708 8560 19760 8566
rect 19708 8502 19760 8508
rect 19856 7644 20164 7653
rect 19856 7642 19862 7644
rect 19918 7642 19942 7644
rect 19998 7642 20022 7644
rect 20078 7642 20102 7644
rect 20158 7642 20164 7644
rect 19918 7590 19920 7642
rect 20100 7590 20102 7642
rect 19856 7588 19862 7590
rect 19918 7588 19942 7590
rect 19998 7588 20022 7590
rect 20078 7588 20102 7590
rect 20158 7588 20164 7590
rect 19856 7579 20164 7588
rect 20732 7546 20760 8842
rect 20824 8634 20852 10542
rect 20916 10538 20944 10950
rect 21008 10742 21036 12582
rect 21088 11212 21140 11218
rect 21088 11154 21140 11160
rect 20996 10736 21048 10742
rect 20996 10678 21048 10684
rect 20904 10532 20956 10538
rect 20904 10474 20956 10480
rect 21100 9518 21128 11154
rect 21272 11008 21324 11014
rect 21272 10950 21324 10956
rect 21284 10713 21312 10950
rect 21270 10704 21326 10713
rect 21270 10639 21326 10648
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 21100 8634 21128 9454
rect 21192 9450 21220 9862
rect 21180 9444 21232 9450
rect 21180 9386 21232 9392
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 21192 8294 21220 9386
rect 21284 8566 21312 10639
rect 21272 8560 21324 8566
rect 21272 8502 21324 8508
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 19856 6556 20164 6565
rect 19856 6554 19862 6556
rect 19918 6554 19942 6556
rect 19998 6554 20022 6556
rect 20078 6554 20102 6556
rect 20158 6554 20164 6556
rect 19918 6502 19920 6554
rect 20100 6502 20102 6554
rect 19856 6500 19862 6502
rect 19918 6500 19942 6502
rect 19998 6500 20022 6502
rect 20078 6500 20102 6502
rect 20158 6500 20164 6502
rect 19856 6491 20164 6500
rect 21284 6118 21312 7686
rect 21376 7478 21404 14436
rect 21456 14418 21508 14424
rect 21468 14006 21496 14418
rect 21456 14000 21508 14006
rect 21456 13942 21508 13948
rect 21560 13870 21588 14962
rect 21824 14340 21876 14346
rect 21824 14282 21876 14288
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 21652 13938 21680 14214
rect 21836 14074 21864 14282
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 21732 14000 21784 14006
rect 21732 13942 21784 13948
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21548 13864 21600 13870
rect 21548 13806 21600 13812
rect 21744 13530 21772 13942
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 22204 13530 22232 13738
rect 21732 13524 21784 13530
rect 21732 13466 21784 13472
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22112 12646 22140 13262
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22112 12442 22140 12582
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22296 11830 22324 15506
rect 22468 14408 22520 14414
rect 22468 14350 22520 14356
rect 22480 13870 22508 14350
rect 22468 13864 22520 13870
rect 22388 13812 22468 13814
rect 22388 13806 22520 13812
rect 22388 13786 22508 13806
rect 22388 13682 22416 13786
rect 22468 13728 22520 13734
rect 22388 13676 22468 13682
rect 22388 13670 22520 13676
rect 22388 13654 22508 13670
rect 22572 13512 22600 15642
rect 22756 14414 22784 19314
rect 23007 19068 23315 19077
rect 23007 19066 23013 19068
rect 23069 19066 23093 19068
rect 23149 19066 23173 19068
rect 23229 19066 23253 19068
rect 23309 19066 23315 19068
rect 23069 19014 23071 19066
rect 23251 19014 23253 19066
rect 23007 19012 23013 19014
rect 23069 19012 23093 19014
rect 23149 19012 23173 19014
rect 23229 19012 23253 19014
rect 23309 19012 23315 19014
rect 23007 19003 23315 19012
rect 22836 18216 22888 18222
rect 22836 18158 22888 18164
rect 22848 17678 22876 18158
rect 23007 17980 23315 17989
rect 23007 17978 23013 17980
rect 23069 17978 23093 17980
rect 23149 17978 23173 17980
rect 23229 17978 23253 17980
rect 23309 17978 23315 17980
rect 23069 17926 23071 17978
rect 23251 17926 23253 17978
rect 23007 17924 23013 17926
rect 23069 17924 23093 17926
rect 23149 17924 23173 17926
rect 23229 17924 23253 17926
rect 23309 17924 23315 17926
rect 23007 17915 23315 17924
rect 23400 17678 23428 19774
rect 23676 19378 23704 20198
rect 23860 19854 23888 20402
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 23848 19712 23900 19718
rect 23848 19654 23900 19660
rect 23664 19372 23716 19378
rect 23664 19314 23716 19320
rect 23480 19304 23532 19310
rect 23480 19246 23532 19252
rect 23492 18970 23520 19246
rect 23664 19168 23716 19174
rect 23664 19110 23716 19116
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23676 18834 23704 19110
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 23756 18352 23808 18358
rect 23756 18294 23808 18300
rect 23768 17882 23796 18294
rect 23756 17876 23808 17882
rect 23756 17818 23808 17824
rect 22836 17672 22888 17678
rect 22836 17614 22888 17620
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23664 17536 23716 17542
rect 23664 17478 23716 17484
rect 23007 16892 23315 16901
rect 23007 16890 23013 16892
rect 23069 16890 23093 16892
rect 23149 16890 23173 16892
rect 23229 16890 23253 16892
rect 23309 16890 23315 16892
rect 23069 16838 23071 16890
rect 23251 16838 23253 16890
rect 23007 16836 23013 16838
rect 23069 16836 23093 16838
rect 23149 16836 23173 16838
rect 23229 16836 23253 16838
rect 23309 16836 23315 16838
rect 23007 16827 23315 16836
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 23400 16182 23428 16390
rect 23388 16176 23440 16182
rect 23388 16118 23440 16124
rect 23007 15804 23315 15813
rect 23007 15802 23013 15804
rect 23069 15802 23093 15804
rect 23149 15802 23173 15804
rect 23229 15802 23253 15804
rect 23309 15802 23315 15804
rect 23069 15750 23071 15802
rect 23251 15750 23253 15802
rect 23007 15748 23013 15750
rect 23069 15748 23093 15750
rect 23149 15748 23173 15750
rect 23229 15748 23253 15750
rect 23309 15748 23315 15750
rect 23007 15739 23315 15748
rect 23492 15706 23520 16594
rect 23572 16516 23624 16522
rect 23572 16458 23624 16464
rect 23584 16114 23612 16458
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 23480 15700 23532 15706
rect 23480 15642 23532 15648
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 23112 15360 23164 15366
rect 23112 15302 23164 15308
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22756 13938 22784 14350
rect 22744 13932 22796 13938
rect 22744 13874 22796 13880
rect 22836 13932 22888 13938
rect 22836 13874 22888 13880
rect 22652 13728 22704 13734
rect 22652 13670 22704 13676
rect 22388 13484 22600 13512
rect 22284 11824 22336 11830
rect 22284 11766 22336 11772
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 22020 11218 22048 11494
rect 21548 11212 21600 11218
rect 21548 11154 21600 11160
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21468 9994 21496 11086
rect 21560 10674 21588 11154
rect 21548 10668 21600 10674
rect 21548 10610 21600 10616
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 21836 10266 21864 10406
rect 22112 10266 22140 11698
rect 22204 11218 22324 11234
rect 22192 11212 22324 11218
rect 22244 11206 22324 11212
rect 22192 11154 22244 11160
rect 22296 11082 22324 11206
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 22388 10062 22416 13484
rect 22664 13410 22692 13670
rect 22848 13530 22876 13874
rect 22836 13524 22888 13530
rect 22836 13466 22888 13472
rect 22468 13388 22520 13394
rect 22468 13330 22520 13336
rect 22572 13382 22692 13410
rect 22480 12306 22508 13330
rect 22572 13190 22600 13382
rect 22744 13252 22796 13258
rect 22744 13194 22796 13200
rect 22560 13184 22612 13190
rect 22560 13126 22612 13132
rect 22756 12986 22784 13194
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 22468 12300 22520 12306
rect 22468 12242 22520 12248
rect 22480 11762 22508 12242
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 22480 11218 22508 11698
rect 22560 11552 22612 11558
rect 22560 11494 22612 11500
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22480 10810 22508 11154
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 22572 10606 22600 11494
rect 22652 11076 22704 11082
rect 22652 11018 22704 11024
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 21824 10056 21876 10062
rect 21824 9998 21876 10004
rect 22376 10056 22428 10062
rect 22376 9998 22428 10004
rect 21456 9988 21508 9994
rect 21456 9930 21508 9936
rect 21468 8906 21496 9930
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 21456 8900 21508 8906
rect 21456 8842 21508 8848
rect 21468 7750 21496 8842
rect 21652 7954 21680 9318
rect 21836 8634 21864 9998
rect 22388 9674 22416 9998
rect 22664 9926 22692 11018
rect 22652 9920 22704 9926
rect 22652 9862 22704 9868
rect 22388 9646 22600 9674
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 21928 8634 21956 8774
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21916 8628 21968 8634
rect 21916 8570 21968 8576
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21456 7744 21508 7750
rect 21456 7686 21508 7692
rect 21364 7472 21416 7478
rect 21364 7414 21416 7420
rect 21652 7410 21680 7890
rect 21836 7546 21864 8570
rect 22572 8090 22600 9646
rect 22664 9586 22692 9862
rect 22652 9580 22704 9586
rect 22652 9522 22704 9528
rect 22560 8084 22612 8090
rect 22560 8026 22612 8032
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 21732 7472 21784 7478
rect 21732 7414 21784 7420
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21744 7002 21772 7414
rect 21732 6996 21784 7002
rect 21732 6938 21784 6944
rect 21928 6798 21956 7686
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 21928 6662 21956 6734
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 22020 6186 22048 7278
rect 22112 6798 22140 7686
rect 22204 6798 22232 7822
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22296 7206 22324 7686
rect 22284 7200 22336 7206
rect 22284 7142 22336 7148
rect 22296 6798 22324 7142
rect 22756 7002 22784 11766
rect 22836 11552 22888 11558
rect 22836 11494 22888 11500
rect 22848 9722 22876 11494
rect 22836 9716 22888 9722
rect 22836 9658 22888 9664
rect 22940 7460 22968 15302
rect 23124 15026 23152 15302
rect 23112 15020 23164 15026
rect 23112 14962 23164 14968
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 23007 14716 23315 14725
rect 23007 14714 23013 14716
rect 23069 14714 23093 14716
rect 23149 14714 23173 14716
rect 23229 14714 23253 14716
rect 23309 14714 23315 14716
rect 23069 14662 23071 14714
rect 23251 14662 23253 14714
rect 23007 14660 23013 14662
rect 23069 14660 23093 14662
rect 23149 14660 23173 14662
rect 23229 14660 23253 14662
rect 23309 14660 23315 14662
rect 23007 14651 23315 14660
rect 23400 14618 23428 14758
rect 23296 14612 23348 14618
rect 23296 14554 23348 14560
rect 23388 14612 23440 14618
rect 23388 14554 23440 14560
rect 23204 14408 23256 14414
rect 23204 14350 23256 14356
rect 23216 13870 23244 14350
rect 23308 14346 23336 14554
rect 23296 14340 23348 14346
rect 23296 14282 23348 14288
rect 23204 13864 23256 13870
rect 23204 13806 23256 13812
rect 23308 13814 23336 14282
rect 23400 14278 23428 14554
rect 23480 14476 23532 14482
rect 23480 14418 23532 14424
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23400 13938 23428 14214
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23308 13786 23428 13814
rect 23400 13734 23428 13786
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23007 13628 23315 13637
rect 23007 13626 23013 13628
rect 23069 13626 23093 13628
rect 23149 13626 23173 13628
rect 23229 13626 23253 13628
rect 23309 13626 23315 13628
rect 23069 13574 23071 13626
rect 23251 13574 23253 13626
rect 23007 13572 23013 13574
rect 23069 13572 23093 13574
rect 23149 13572 23173 13574
rect 23229 13572 23253 13574
rect 23309 13572 23315 13574
rect 23007 13563 23315 13572
rect 23400 13512 23428 13670
rect 23308 13484 23428 13512
rect 23308 12646 23336 13484
rect 23492 13394 23520 14418
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23388 13184 23440 13190
rect 23388 13126 23440 13132
rect 23296 12640 23348 12646
rect 23296 12582 23348 12588
rect 23007 12540 23315 12549
rect 23007 12538 23013 12540
rect 23069 12538 23093 12540
rect 23149 12538 23173 12540
rect 23229 12538 23253 12540
rect 23309 12538 23315 12540
rect 23069 12486 23071 12538
rect 23251 12486 23253 12538
rect 23007 12484 23013 12486
rect 23069 12484 23093 12486
rect 23149 12484 23173 12486
rect 23229 12484 23253 12486
rect 23309 12484 23315 12486
rect 23007 12475 23315 12484
rect 23007 11452 23315 11461
rect 23007 11450 23013 11452
rect 23069 11450 23093 11452
rect 23149 11450 23173 11452
rect 23229 11450 23253 11452
rect 23309 11450 23315 11452
rect 23069 11398 23071 11450
rect 23251 11398 23253 11450
rect 23007 11396 23013 11398
rect 23069 11396 23093 11398
rect 23149 11396 23173 11398
rect 23229 11396 23253 11398
rect 23309 11396 23315 11398
rect 23007 11387 23315 11396
rect 23400 11150 23428 13126
rect 23492 12850 23520 13330
rect 23480 12844 23532 12850
rect 23480 12786 23532 12792
rect 23480 11688 23532 11694
rect 23480 11630 23532 11636
rect 23492 11354 23520 11630
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 23007 10364 23315 10373
rect 23007 10362 23013 10364
rect 23069 10362 23093 10364
rect 23149 10362 23173 10364
rect 23229 10362 23253 10364
rect 23309 10362 23315 10364
rect 23069 10310 23071 10362
rect 23251 10310 23253 10362
rect 23007 10308 23013 10310
rect 23069 10308 23093 10310
rect 23149 10308 23173 10310
rect 23229 10308 23253 10310
rect 23309 10308 23315 10310
rect 23007 10299 23315 10308
rect 23400 10266 23428 11086
rect 23388 10260 23440 10266
rect 23388 10202 23440 10208
rect 23007 9276 23315 9285
rect 23007 9274 23013 9276
rect 23069 9274 23093 9276
rect 23149 9274 23173 9276
rect 23229 9274 23253 9276
rect 23309 9274 23315 9276
rect 23069 9222 23071 9274
rect 23251 9222 23253 9274
rect 23007 9220 23013 9222
rect 23069 9220 23093 9222
rect 23149 9220 23173 9222
rect 23229 9220 23253 9222
rect 23309 9220 23315 9222
rect 23007 9211 23315 9220
rect 23572 8832 23624 8838
rect 23676 8820 23704 17478
rect 23860 15194 23888 19654
rect 23952 17678 23980 20402
rect 24044 19514 24072 20402
rect 24492 20052 24544 20058
rect 24492 19994 24544 20000
rect 24504 19854 24532 19994
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24124 19712 24176 19718
rect 24124 19654 24176 19660
rect 24032 19508 24084 19514
rect 24032 19450 24084 19456
rect 24136 17882 24164 19654
rect 24504 19310 24532 19790
rect 24492 19304 24544 19310
rect 24492 19246 24544 19252
rect 24492 18624 24544 18630
rect 24492 18566 24544 18572
rect 24504 18426 24532 18566
rect 24492 18420 24544 18426
rect 24492 18362 24544 18368
rect 24124 17876 24176 17882
rect 24124 17818 24176 17824
rect 23940 17672 23992 17678
rect 23940 17614 23992 17620
rect 24780 17202 24808 19790
rect 24860 18216 24912 18222
rect 24860 18158 24912 18164
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 24768 17196 24820 17202
rect 24768 17138 24820 17144
rect 23952 16794 23980 17138
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 24872 16250 24900 18158
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 24492 16108 24544 16114
rect 24492 16050 24544 16056
rect 24032 15904 24084 15910
rect 24032 15846 24084 15852
rect 24044 15706 24072 15846
rect 24032 15700 24084 15706
rect 24032 15642 24084 15648
rect 23768 15166 23888 15194
rect 23768 12918 23796 15166
rect 24504 15094 24532 16050
rect 24492 15088 24544 15094
rect 24492 15030 24544 15036
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 24216 14408 24268 14414
rect 24216 14350 24268 14356
rect 24032 14000 24084 14006
rect 24032 13942 24084 13948
rect 24044 13326 24072 13942
rect 24228 13530 24256 14350
rect 24596 14074 24624 14554
rect 25056 14414 25084 14758
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 24584 14068 24636 14074
rect 24584 14010 24636 14016
rect 24400 13864 24452 13870
rect 24400 13806 24452 13812
rect 24412 13530 24440 13806
rect 24216 13524 24268 13530
rect 24216 13466 24268 13472
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 24044 12918 24072 13262
rect 24688 12986 24716 14350
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 24964 13530 24992 14214
rect 25056 13530 25084 14350
rect 25148 13546 25176 20402
rect 25228 19848 25280 19854
rect 25228 19790 25280 19796
rect 25240 19378 25268 19790
rect 25412 19712 25464 19718
rect 25412 19654 25464 19660
rect 25228 19372 25280 19378
rect 25228 19314 25280 19320
rect 25240 18766 25268 19314
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 25424 17746 25452 19654
rect 25412 17740 25464 17746
rect 25412 17682 25464 17688
rect 25516 16574 25544 22066
rect 26158 21788 26466 21797
rect 26158 21786 26164 21788
rect 26220 21786 26244 21788
rect 26300 21786 26324 21788
rect 26380 21786 26404 21788
rect 26460 21786 26466 21788
rect 26220 21734 26222 21786
rect 26402 21734 26404 21786
rect 26158 21732 26164 21734
rect 26220 21732 26244 21734
rect 26300 21732 26324 21734
rect 26380 21732 26404 21734
rect 26460 21732 26466 21734
rect 26158 21723 26466 21732
rect 25688 21548 25740 21554
rect 25688 21490 25740 21496
rect 25700 20602 25728 21490
rect 25872 21344 25924 21350
rect 25872 21286 25924 21292
rect 25884 21185 25912 21286
rect 25870 21176 25926 21185
rect 25870 21111 25926 21120
rect 26158 20700 26466 20709
rect 26158 20698 26164 20700
rect 26220 20698 26244 20700
rect 26300 20698 26324 20700
rect 26380 20698 26404 20700
rect 26460 20698 26466 20700
rect 26220 20646 26222 20698
rect 26402 20646 26404 20698
rect 26158 20644 26164 20646
rect 26220 20644 26244 20646
rect 26300 20644 26324 20646
rect 26380 20644 26404 20646
rect 26460 20644 26466 20646
rect 26158 20635 26466 20644
rect 25688 20596 25740 20602
rect 25688 20538 25740 20544
rect 26158 19612 26466 19621
rect 26158 19610 26164 19612
rect 26220 19610 26244 19612
rect 26300 19610 26324 19612
rect 26380 19610 26404 19612
rect 26460 19610 26466 19612
rect 26220 19558 26222 19610
rect 26402 19558 26404 19610
rect 26158 19556 26164 19558
rect 26220 19556 26244 19558
rect 26300 19556 26324 19558
rect 26380 19556 26404 19558
rect 26460 19556 26466 19558
rect 26158 19547 26466 19556
rect 26158 18524 26466 18533
rect 26158 18522 26164 18524
rect 26220 18522 26244 18524
rect 26300 18522 26324 18524
rect 26380 18522 26404 18524
rect 26460 18522 26466 18524
rect 26220 18470 26222 18522
rect 26402 18470 26404 18522
rect 26158 18468 26164 18470
rect 26220 18468 26244 18470
rect 26300 18468 26324 18470
rect 26380 18468 26404 18470
rect 26460 18468 26466 18470
rect 26158 18459 26466 18468
rect 26158 17436 26466 17445
rect 26158 17434 26164 17436
rect 26220 17434 26244 17436
rect 26300 17434 26324 17436
rect 26380 17434 26404 17436
rect 26460 17434 26466 17436
rect 26220 17382 26222 17434
rect 26402 17382 26404 17434
rect 26158 17380 26164 17382
rect 26220 17380 26244 17382
rect 26300 17380 26324 17382
rect 26380 17380 26404 17382
rect 26460 17380 26466 17382
rect 26158 17371 26466 17380
rect 26332 17128 26384 17134
rect 26330 17096 26332 17105
rect 26384 17096 26386 17105
rect 26330 17031 26386 17040
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25424 16546 25544 16574
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25240 15094 25268 15302
rect 25228 15088 25280 15094
rect 25228 15030 25280 15036
rect 25320 13728 25372 13734
rect 25320 13670 25372 13676
rect 24952 13524 25004 13530
rect 24952 13466 25004 13472
rect 25044 13524 25096 13530
rect 25148 13518 25268 13546
rect 25044 13466 25096 13472
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 24032 12912 24084 12918
rect 24032 12854 24084 12860
rect 24044 11830 24072 12854
rect 24780 11898 24808 13262
rect 25148 12646 25176 13330
rect 25240 12782 25268 13518
rect 25332 13326 25360 13670
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25228 12776 25280 12782
rect 25424 12753 25452 16546
rect 25608 16266 25636 16934
rect 26158 16348 26466 16357
rect 26158 16346 26164 16348
rect 26220 16346 26244 16348
rect 26300 16346 26324 16348
rect 26380 16346 26404 16348
rect 26460 16346 26466 16348
rect 26220 16294 26222 16346
rect 26402 16294 26404 16346
rect 26158 16292 26164 16294
rect 26220 16292 26244 16294
rect 26300 16292 26324 16294
rect 26380 16292 26404 16294
rect 26460 16292 26466 16294
rect 26158 16283 26466 16292
rect 25516 16238 25636 16266
rect 25516 16182 25544 16238
rect 25504 16176 25556 16182
rect 25504 16118 25556 16124
rect 25780 16040 25832 16046
rect 25780 15982 25832 15988
rect 25792 15026 25820 15982
rect 26158 15260 26466 15269
rect 26158 15258 26164 15260
rect 26220 15258 26244 15260
rect 26300 15258 26324 15260
rect 26380 15258 26404 15260
rect 26460 15258 26466 15260
rect 26220 15206 26222 15258
rect 26402 15206 26404 15258
rect 26158 15204 26164 15206
rect 26220 15204 26244 15206
rect 26300 15204 26324 15206
rect 26380 15204 26404 15206
rect 26460 15204 26466 15206
rect 26158 15195 26466 15204
rect 27080 15162 27108 28809
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 25780 15020 25832 15026
rect 25780 14962 25832 14968
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25700 14006 25728 14214
rect 26158 14172 26466 14181
rect 26158 14170 26164 14172
rect 26220 14170 26244 14172
rect 26300 14170 26324 14172
rect 26380 14170 26404 14172
rect 26460 14170 26466 14172
rect 26220 14118 26222 14170
rect 26402 14118 26404 14170
rect 26158 14116 26164 14118
rect 26220 14116 26244 14118
rect 26300 14116 26324 14118
rect 26380 14116 26404 14118
rect 26460 14116 26466 14118
rect 26158 14107 26466 14116
rect 25688 14000 25740 14006
rect 25688 13942 25740 13948
rect 25688 13864 25740 13870
rect 25688 13806 25740 13812
rect 25700 13530 25728 13806
rect 25688 13524 25740 13530
rect 25688 13466 25740 13472
rect 25872 13456 25924 13462
rect 25872 13398 25924 13404
rect 25688 13320 25740 13326
rect 25884 13297 25912 13398
rect 25688 13262 25740 13268
rect 25870 13288 25926 13297
rect 25228 12718 25280 12724
rect 25410 12744 25466 12753
rect 25410 12679 25466 12688
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 25700 11898 25728 13262
rect 25870 13223 25926 13232
rect 26158 13084 26466 13093
rect 26158 13082 26164 13084
rect 26220 13082 26244 13084
rect 26300 13082 26324 13084
rect 26380 13082 26404 13084
rect 26460 13082 26466 13084
rect 26220 13030 26222 13082
rect 26402 13030 26404 13082
rect 26158 13028 26164 13030
rect 26220 13028 26244 13030
rect 26300 13028 26324 13030
rect 26380 13028 26404 13030
rect 26460 13028 26466 13030
rect 26158 13019 26466 13028
rect 26158 11996 26466 12005
rect 26158 11994 26164 11996
rect 26220 11994 26244 11996
rect 26300 11994 26324 11996
rect 26380 11994 26404 11996
rect 26460 11994 26466 11996
rect 26220 11942 26222 11994
rect 26402 11942 26404 11994
rect 26158 11940 26164 11942
rect 26220 11940 26244 11942
rect 26300 11940 26324 11942
rect 26380 11940 26404 11942
rect 26460 11940 26466 11942
rect 26158 11931 26466 11940
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 25688 11892 25740 11898
rect 25688 11834 25740 11840
rect 24032 11824 24084 11830
rect 24032 11766 24084 11772
rect 24044 11054 24072 11766
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 24044 11026 24164 11054
rect 24136 10742 24164 11026
rect 24400 11008 24452 11014
rect 24400 10950 24452 10956
rect 23848 10736 23900 10742
rect 23848 10678 23900 10684
rect 24124 10736 24176 10742
rect 24124 10678 24176 10684
rect 23860 10130 23888 10678
rect 24412 10606 24440 10950
rect 24216 10600 24268 10606
rect 24216 10542 24268 10548
rect 24400 10600 24452 10606
rect 24400 10542 24452 10548
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 24228 10266 24256 10542
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 23848 10124 23900 10130
rect 23848 10066 23900 10072
rect 23860 9994 23888 10066
rect 24216 10056 24268 10062
rect 24216 9998 24268 10004
rect 23848 9988 23900 9994
rect 23848 9930 23900 9936
rect 23940 9988 23992 9994
rect 23940 9930 23992 9936
rect 23860 9654 23888 9930
rect 23848 9648 23900 9654
rect 23848 9590 23900 9596
rect 23860 8974 23888 9590
rect 23848 8968 23900 8974
rect 23848 8910 23900 8916
rect 23624 8792 23704 8820
rect 23572 8774 23624 8780
rect 23952 8634 23980 9930
rect 24228 8974 24256 9998
rect 24412 9722 24440 10542
rect 24400 9716 24452 9722
rect 24400 9658 24452 9664
rect 24964 9586 24992 10542
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 25148 9586 25176 9998
rect 25332 9654 25360 11290
rect 25688 11144 25740 11150
rect 25688 11086 25740 11092
rect 25504 10464 25556 10470
rect 25504 10406 25556 10412
rect 25516 9994 25544 10406
rect 25504 9988 25556 9994
rect 25504 9930 25556 9936
rect 25320 9648 25372 9654
rect 25320 9590 25372 9596
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 25136 9580 25188 9586
rect 25136 9522 25188 9528
rect 25332 9058 25360 9590
rect 25700 9382 25728 11086
rect 26158 10908 26466 10917
rect 26158 10906 26164 10908
rect 26220 10906 26244 10908
rect 26300 10906 26324 10908
rect 26380 10906 26404 10908
rect 26460 10906 26466 10908
rect 26220 10854 26222 10906
rect 26402 10854 26404 10906
rect 26158 10852 26164 10854
rect 26220 10852 26244 10854
rect 26300 10852 26324 10854
rect 26380 10852 26404 10854
rect 26460 10852 26466 10854
rect 26158 10843 26466 10852
rect 25780 10600 25832 10606
rect 25780 10542 25832 10548
rect 25792 10266 25820 10542
rect 25780 10260 25832 10266
rect 25780 10202 25832 10208
rect 25872 10056 25924 10062
rect 25872 9998 25924 10004
rect 25884 9722 25912 9998
rect 26158 9820 26466 9829
rect 26158 9818 26164 9820
rect 26220 9818 26244 9820
rect 26300 9818 26324 9820
rect 26380 9818 26404 9820
rect 26460 9818 26466 9820
rect 26220 9766 26222 9818
rect 26402 9766 26404 9818
rect 26158 9764 26164 9766
rect 26220 9764 26244 9766
rect 26300 9764 26324 9766
rect 26380 9764 26404 9766
rect 26460 9764 26466 9766
rect 26158 9755 26466 9764
rect 25872 9716 25924 9722
rect 25872 9658 25924 9664
rect 25688 9376 25740 9382
rect 25688 9318 25740 9324
rect 25332 9030 25452 9058
rect 24216 8968 24268 8974
rect 24216 8910 24268 8916
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 24228 8566 24256 8910
rect 25320 8900 25372 8906
rect 25320 8842 25372 8848
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 24216 8560 24268 8566
rect 24216 8502 24268 8508
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 23007 8188 23315 8197
rect 23007 8186 23013 8188
rect 23069 8186 23093 8188
rect 23149 8186 23173 8188
rect 23229 8186 23253 8188
rect 23309 8186 23315 8188
rect 23069 8134 23071 8186
rect 23251 8134 23253 8186
rect 23007 8132 23013 8134
rect 23069 8132 23093 8134
rect 23149 8132 23173 8134
rect 23229 8132 23253 8134
rect 23309 8132 23315 8134
rect 23007 8123 23315 8132
rect 23020 7472 23072 7478
rect 22940 7432 23020 7460
rect 23020 7414 23072 7420
rect 23007 7100 23315 7109
rect 23007 7098 23013 7100
rect 23069 7098 23093 7100
rect 23149 7098 23173 7100
rect 23229 7098 23253 7100
rect 23309 7098 23315 7100
rect 23069 7046 23071 7098
rect 23251 7046 23253 7098
rect 23007 7044 23013 7046
rect 23069 7044 23093 7046
rect 23149 7044 23173 7046
rect 23229 7044 23253 7046
rect 23309 7044 23315 7046
rect 23007 7035 23315 7044
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 22376 6928 22428 6934
rect 22376 6870 22428 6876
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22284 6792 22336 6798
rect 22284 6734 22336 6740
rect 22008 6180 22060 6186
rect 22008 6122 22060 6128
rect 21272 6112 21324 6118
rect 21272 6054 21324 6060
rect 21548 6112 21600 6118
rect 21548 6054 21600 6060
rect 18512 5714 18564 5720
rect 18420 5636 18472 5642
rect 18420 5578 18472 5584
rect 18432 5302 18460 5578
rect 18420 5296 18472 5302
rect 18420 5238 18472 5244
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 18236 5092 18288 5098
rect 18236 5034 18288 5040
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 18064 4146 18092 4558
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 17092 3420 17264 3448
rect 17040 3402 17092 3408
rect 16592 3194 16620 3402
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 17052 3126 17080 3402
rect 17880 3194 17908 4082
rect 18064 3738 18092 4082
rect 18524 4078 18552 5714
rect 18800 5710 18828 5766
rect 18972 5772 19024 5778
rect 18972 5714 19024 5720
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19616 5772 19668 5778
rect 19616 5714 19668 5720
rect 18696 5704 18748 5710
rect 18696 5646 18748 5652
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18708 5574 18736 5646
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18708 5370 18736 5510
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 18800 4826 18828 5646
rect 21284 5574 21312 6054
rect 21560 5778 21588 6054
rect 21548 5772 21600 5778
rect 21548 5714 21600 5720
rect 22112 5574 22140 6734
rect 22204 6118 22232 6734
rect 22388 6458 22416 6870
rect 22560 6724 22612 6730
rect 22560 6666 22612 6672
rect 22376 6452 22428 6458
rect 22376 6394 22428 6400
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22572 5914 22600 6666
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 21272 5568 21324 5574
rect 21272 5510 21324 5516
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 18972 5160 19024 5166
rect 18972 5102 19024 5108
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 18248 3534 18276 3878
rect 18892 3602 18920 4966
rect 18984 4826 19012 5102
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 19076 4622 19104 5510
rect 19856 5468 20164 5477
rect 19856 5466 19862 5468
rect 19918 5466 19942 5468
rect 19998 5466 20022 5468
rect 20078 5466 20102 5468
rect 20158 5466 20164 5468
rect 19918 5414 19920 5466
rect 20100 5414 20102 5466
rect 19856 5412 19862 5414
rect 19918 5412 19942 5414
rect 19998 5412 20022 5414
rect 20078 5412 20102 5414
rect 20158 5412 20164 5414
rect 19856 5403 20164 5412
rect 21284 5302 21312 5510
rect 21272 5296 21324 5302
rect 21272 5238 21324 5244
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 19856 4380 20164 4389
rect 19856 4378 19862 4380
rect 19918 4378 19942 4380
rect 19998 4378 20022 4380
rect 20078 4378 20102 4380
rect 20158 4378 20164 4380
rect 19918 4326 19920 4378
rect 20100 4326 20102 4378
rect 19856 4324 19862 4326
rect 19918 4324 19942 4326
rect 19998 4324 20022 4326
rect 20078 4324 20102 4326
rect 20158 4324 20164 4326
rect 19856 4315 20164 4324
rect 21284 4214 21312 5238
rect 22572 5166 22600 5850
rect 22756 5710 22784 6938
rect 22928 6928 22980 6934
rect 23112 6928 23164 6934
rect 22980 6888 23112 6916
rect 22928 6870 22980 6876
rect 23112 6870 23164 6876
rect 22928 6792 22980 6798
rect 23112 6792 23164 6798
rect 22980 6752 23112 6780
rect 22928 6734 22980 6740
rect 23112 6734 23164 6740
rect 22836 6384 22888 6390
rect 22836 6326 22888 6332
rect 22848 6118 22876 6326
rect 23400 6202 23428 8366
rect 23676 7954 23704 8434
rect 24964 7954 24992 8774
rect 25136 8424 25188 8430
rect 25136 8366 25188 8372
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 24952 7948 25004 7954
rect 24952 7890 25004 7896
rect 23676 7342 23704 7890
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24136 7546 24164 7686
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 23664 7336 23716 7342
rect 23664 7278 23716 7284
rect 23676 6458 23704 7278
rect 25148 7002 25176 8366
rect 25228 8288 25280 8294
rect 25228 8230 25280 8236
rect 25240 7478 25268 8230
rect 25332 7954 25360 8842
rect 25320 7948 25372 7954
rect 25320 7890 25372 7896
rect 25424 7546 25452 9030
rect 25700 8634 25728 9318
rect 26158 8732 26466 8741
rect 26158 8730 26164 8732
rect 26220 8730 26244 8732
rect 26300 8730 26324 8732
rect 26380 8730 26404 8732
rect 26460 8730 26466 8732
rect 26220 8678 26222 8730
rect 26402 8678 26404 8730
rect 26158 8676 26164 8678
rect 26220 8676 26244 8678
rect 26300 8676 26324 8678
rect 26380 8676 26404 8678
rect 26460 8676 26466 8678
rect 26158 8667 26466 8676
rect 25688 8628 25740 8634
rect 25688 8570 25740 8576
rect 25962 8256 26018 8265
rect 25962 8191 26018 8200
rect 25976 7954 26004 8191
rect 25964 7948 26016 7954
rect 25964 7890 26016 7896
rect 26158 7644 26466 7653
rect 26158 7642 26164 7644
rect 26220 7642 26244 7644
rect 26300 7642 26324 7644
rect 26380 7642 26404 7644
rect 26460 7642 26466 7644
rect 26220 7590 26222 7642
rect 26402 7590 26404 7642
rect 26158 7588 26164 7590
rect 26220 7588 26244 7590
rect 26300 7588 26324 7590
rect 26380 7588 26404 7590
rect 26460 7588 26466 7590
rect 26158 7579 26466 7588
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25228 7472 25280 7478
rect 25228 7414 25280 7420
rect 23848 6996 23900 7002
rect 23848 6938 23900 6944
rect 25136 6996 25188 7002
rect 25136 6938 25188 6944
rect 23860 6662 23888 6938
rect 25424 6866 25452 7482
rect 25412 6860 25464 6866
rect 25412 6802 25464 6808
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 26158 6556 26466 6565
rect 26158 6554 26164 6556
rect 26220 6554 26244 6556
rect 26300 6554 26324 6556
rect 26380 6554 26404 6556
rect 26460 6554 26466 6556
rect 26220 6502 26222 6554
rect 26402 6502 26404 6554
rect 26158 6500 26164 6502
rect 26220 6500 26244 6502
rect 26300 6500 26324 6502
rect 26380 6500 26404 6502
rect 26460 6500 26466 6502
rect 26158 6491 26466 6500
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23676 6322 23704 6394
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23400 6186 23612 6202
rect 23400 6180 23624 6186
rect 23400 6174 23572 6180
rect 23572 6122 23624 6128
rect 22836 6112 22888 6118
rect 22836 6054 22888 6060
rect 23480 6112 23532 6118
rect 23480 6054 23532 6060
rect 23007 6012 23315 6021
rect 23007 6010 23013 6012
rect 23069 6010 23093 6012
rect 23149 6010 23173 6012
rect 23229 6010 23253 6012
rect 23309 6010 23315 6012
rect 23069 5958 23071 6010
rect 23251 5958 23253 6010
rect 23007 5956 23013 5958
rect 23069 5956 23093 5958
rect 23149 5956 23173 5958
rect 23229 5956 23253 5958
rect 23309 5956 23315 5958
rect 23007 5947 23315 5956
rect 22744 5704 22796 5710
rect 22744 5646 22796 5652
rect 23492 5370 23520 6054
rect 23676 5778 23704 6258
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 23664 5772 23716 5778
rect 23664 5714 23716 5720
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 22560 5160 22612 5166
rect 22560 5102 22612 5108
rect 21272 4208 21324 4214
rect 21272 4150 21324 4156
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18340 3194 18368 3334
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 17040 3120 17092 3126
rect 17040 3062 17092 3068
rect 18892 2990 18920 3538
rect 21284 3466 21312 4150
rect 22572 4078 22600 5102
rect 23007 4924 23315 4933
rect 23007 4922 23013 4924
rect 23069 4922 23093 4924
rect 23149 4922 23173 4924
rect 23229 4922 23253 4924
rect 23309 4922 23315 4924
rect 23069 4870 23071 4922
rect 23251 4870 23253 4922
rect 23007 4868 23013 4870
rect 23069 4868 23093 4870
rect 23149 4868 23173 4870
rect 23229 4868 23253 4870
rect 23309 4868 23315 4870
rect 23007 4859 23315 4868
rect 23676 4146 23704 5714
rect 23664 4140 23716 4146
rect 23664 4082 23716 4088
rect 22560 4072 22612 4078
rect 22560 4014 22612 4020
rect 22836 4072 22888 4078
rect 22836 4014 22888 4020
rect 22848 3738 22876 4014
rect 23007 3836 23315 3845
rect 23007 3834 23013 3836
rect 23069 3834 23093 3836
rect 23149 3834 23173 3836
rect 23229 3834 23253 3836
rect 23309 3834 23315 3836
rect 23069 3782 23071 3834
rect 23251 3782 23253 3834
rect 23007 3780 23013 3782
rect 23069 3780 23093 3782
rect 23149 3780 23173 3782
rect 23229 3780 23253 3782
rect 23309 3780 23315 3782
rect 23007 3771 23315 3780
rect 22836 3732 22888 3738
rect 22836 3674 22888 3680
rect 20260 3460 20312 3466
rect 20260 3402 20312 3408
rect 21272 3460 21324 3466
rect 21272 3402 21324 3408
rect 19856 3292 20164 3301
rect 19856 3290 19862 3292
rect 19918 3290 19942 3292
rect 19998 3290 20022 3292
rect 20078 3290 20102 3292
rect 20158 3290 20164 3292
rect 19918 3238 19920 3290
rect 20100 3238 20102 3290
rect 19856 3236 19862 3238
rect 19918 3236 19942 3238
rect 19998 3236 20022 3238
rect 20078 3236 20102 3238
rect 20158 3236 20164 3238
rect 19856 3227 20164 3236
rect 18880 2984 18932 2990
rect 18880 2926 18932 2932
rect 15856 2746 15976 2774
rect 16316 2746 16436 2774
rect 15948 2446 15976 2746
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 16408 2378 16436 2746
rect 16705 2748 17013 2757
rect 16705 2746 16711 2748
rect 16767 2746 16791 2748
rect 16847 2746 16871 2748
rect 16927 2746 16951 2748
rect 17007 2746 17013 2748
rect 16767 2694 16769 2746
rect 16949 2694 16951 2746
rect 16705 2692 16711 2694
rect 16767 2692 16791 2694
rect 16847 2692 16871 2694
rect 16927 2692 16951 2694
rect 17007 2692 17013 2694
rect 16705 2683 17013 2692
rect 20272 2650 20300 3402
rect 23007 2748 23315 2757
rect 23007 2746 23013 2748
rect 23069 2746 23093 2748
rect 23149 2746 23173 2748
rect 23229 2746 23253 2748
rect 23309 2746 23315 2748
rect 23069 2694 23071 2746
rect 23251 2694 23253 2746
rect 23007 2692 23013 2694
rect 23069 2692 23093 2694
rect 23149 2692 23173 2694
rect 23229 2692 23253 2694
rect 23309 2692 23315 2694
rect 23007 2683 23315 2692
rect 25148 2650 25176 6190
rect 26158 5468 26466 5477
rect 26158 5466 26164 5468
rect 26220 5466 26244 5468
rect 26300 5466 26324 5468
rect 26380 5466 26404 5468
rect 26460 5466 26466 5468
rect 26220 5414 26222 5466
rect 26402 5414 26404 5466
rect 26158 5412 26164 5414
rect 26220 5412 26244 5414
rect 26300 5412 26324 5414
rect 26380 5412 26404 5414
rect 26460 5412 26466 5414
rect 26158 5403 26466 5412
rect 25964 4480 26016 4486
rect 25964 4422 26016 4428
rect 25976 4185 26004 4422
rect 26158 4380 26466 4389
rect 26158 4378 26164 4380
rect 26220 4378 26244 4380
rect 26300 4378 26324 4380
rect 26380 4378 26404 4380
rect 26460 4378 26466 4380
rect 26220 4326 26222 4378
rect 26402 4326 26404 4378
rect 26158 4324 26164 4326
rect 26220 4324 26244 4326
rect 26300 4324 26324 4326
rect 26380 4324 26404 4326
rect 26460 4324 26466 4326
rect 26158 4315 26466 4324
rect 25962 4176 26018 4185
rect 25962 4111 26018 4120
rect 26158 3292 26466 3301
rect 26158 3290 26164 3292
rect 26220 3290 26244 3292
rect 26300 3290 26324 3292
rect 26380 3290 26404 3292
rect 26460 3290 26466 3292
rect 26220 3238 26222 3290
rect 26402 3238 26404 3290
rect 26158 3236 26164 3238
rect 26220 3236 26244 3238
rect 26300 3236 26324 3238
rect 26380 3236 26404 3238
rect 26460 3236 26466 3238
rect 26158 3227 26466 3236
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 25136 2644 25188 2650
rect 25136 2586 25188 2592
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 11704 2372 11756 2378
rect 11704 2314 11756 2320
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 16396 2372 16448 2378
rect 16396 2314 16448 2320
rect 32 800 60 2314
rect 3988 1170 4016 2314
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7252 2204 7560 2213
rect 7252 2202 7258 2204
rect 7314 2202 7338 2204
rect 7394 2202 7418 2204
rect 7474 2202 7498 2204
rect 7554 2202 7560 2204
rect 7314 2150 7316 2202
rect 7496 2150 7498 2202
rect 7252 2148 7258 2150
rect 7314 2148 7338 2150
rect 7394 2148 7418 2150
rect 7474 2148 7498 2150
rect 7554 2148 7560 2150
rect 7252 2139 7560 2148
rect 3896 1142 4016 1170
rect 3896 800 3924 1142
rect 7760 800 7788 2246
rect 11716 1170 11744 2314
rect 13554 2204 13862 2213
rect 13554 2202 13560 2204
rect 13616 2202 13640 2204
rect 13696 2202 13720 2204
rect 13776 2202 13800 2204
rect 13856 2202 13862 2204
rect 13616 2150 13618 2202
rect 13798 2150 13800 2202
rect 13554 2148 13560 2150
rect 13616 2148 13640 2150
rect 13696 2148 13720 2150
rect 13776 2148 13800 2150
rect 13856 2148 13862 2150
rect 13554 2139 13862 2148
rect 15580 1170 15608 2314
rect 19856 2204 20164 2213
rect 19856 2202 19862 2204
rect 19918 2202 19942 2204
rect 19998 2202 20022 2204
rect 20078 2202 20102 2204
rect 20158 2202 20164 2204
rect 19918 2150 19920 2202
rect 20100 2150 20102 2202
rect 19856 2148 19862 2150
rect 19918 2148 19942 2150
rect 19998 2148 20022 2150
rect 20078 2148 20102 2150
rect 20158 2148 20164 2150
rect 19856 2139 20164 2148
rect 11624 1142 11744 1170
rect 15488 1142 15608 1170
rect 11624 800 11652 1142
rect 15488 800 15516 1142
rect 19996 870 20116 898
rect 19996 800 20024 870
rect 18 0 74 800
rect 3882 0 3938 800
rect 7746 0 7802 800
rect 11610 0 11666 800
rect 15474 0 15530 800
rect 19982 0 20038 800
rect 20088 762 20116 870
rect 20272 762 20300 2382
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 23860 800 23888 2246
rect 20088 734 20300 762
rect 23846 0 23902 800
rect 24780 105 24808 2246
rect 26158 2204 26466 2213
rect 26158 2202 26164 2204
rect 26220 2202 26244 2204
rect 26300 2202 26324 2204
rect 26380 2202 26404 2204
rect 26460 2202 26466 2204
rect 26220 2150 26222 2202
rect 26402 2150 26404 2202
rect 26158 2148 26164 2150
rect 26220 2148 26244 2150
rect 26300 2148 26324 2150
rect 26380 2148 26404 2150
rect 26460 2148 26466 2150
rect 26158 2139 26466 2148
rect 24766 96 24822 105
rect 24766 31 24822 40
<< via2 >>
rect 2778 29280 2834 29336
rect 7258 27226 7314 27228
rect 7338 27226 7394 27228
rect 7418 27226 7474 27228
rect 7498 27226 7554 27228
rect 7258 27174 7304 27226
rect 7304 27174 7314 27226
rect 7338 27174 7368 27226
rect 7368 27174 7380 27226
rect 7380 27174 7394 27226
rect 7418 27174 7432 27226
rect 7432 27174 7444 27226
rect 7444 27174 7474 27226
rect 7498 27174 7508 27226
rect 7508 27174 7554 27226
rect 7258 27172 7314 27174
rect 7338 27172 7394 27174
rect 7418 27172 7474 27174
rect 7498 27172 7554 27174
rect 13560 27226 13616 27228
rect 13640 27226 13696 27228
rect 13720 27226 13776 27228
rect 13800 27226 13856 27228
rect 13560 27174 13606 27226
rect 13606 27174 13616 27226
rect 13640 27174 13670 27226
rect 13670 27174 13682 27226
rect 13682 27174 13696 27226
rect 13720 27174 13734 27226
rect 13734 27174 13746 27226
rect 13746 27174 13776 27226
rect 13800 27174 13810 27226
rect 13810 27174 13856 27226
rect 13560 27172 13616 27174
rect 13640 27172 13696 27174
rect 13720 27172 13776 27174
rect 13800 27172 13856 27174
rect 19862 27226 19918 27228
rect 19942 27226 19998 27228
rect 20022 27226 20078 27228
rect 20102 27226 20158 27228
rect 19862 27174 19908 27226
rect 19908 27174 19918 27226
rect 19942 27174 19972 27226
rect 19972 27174 19984 27226
rect 19984 27174 19998 27226
rect 20022 27174 20036 27226
rect 20036 27174 20048 27226
rect 20048 27174 20078 27226
rect 20102 27174 20112 27226
rect 20112 27174 20158 27226
rect 19862 27172 19918 27174
rect 19942 27172 19998 27174
rect 20022 27172 20078 27174
rect 20102 27172 20158 27174
rect 26164 27226 26220 27228
rect 26244 27226 26300 27228
rect 26324 27226 26380 27228
rect 26404 27226 26460 27228
rect 26164 27174 26210 27226
rect 26210 27174 26220 27226
rect 26244 27174 26274 27226
rect 26274 27174 26286 27226
rect 26286 27174 26300 27226
rect 26324 27174 26338 27226
rect 26338 27174 26350 27226
rect 26350 27174 26380 27226
rect 26404 27174 26414 27226
rect 26414 27174 26460 27226
rect 26164 27172 26220 27174
rect 26244 27172 26300 27174
rect 26324 27172 26380 27174
rect 26404 27172 26460 27174
rect 938 25236 940 25256
rect 940 25236 992 25256
rect 992 25236 994 25256
rect 938 25200 994 25236
rect 938 21120 994 21176
rect 1490 16496 1546 16552
rect 938 12280 994 12336
rect 1306 8200 1362 8256
rect 4107 26682 4163 26684
rect 4187 26682 4243 26684
rect 4267 26682 4323 26684
rect 4347 26682 4403 26684
rect 4107 26630 4153 26682
rect 4153 26630 4163 26682
rect 4187 26630 4217 26682
rect 4217 26630 4229 26682
rect 4229 26630 4243 26682
rect 4267 26630 4281 26682
rect 4281 26630 4293 26682
rect 4293 26630 4323 26682
rect 4347 26630 4357 26682
rect 4357 26630 4403 26682
rect 4107 26628 4163 26630
rect 4187 26628 4243 26630
rect 4267 26628 4323 26630
rect 4347 26628 4403 26630
rect 4107 25594 4163 25596
rect 4187 25594 4243 25596
rect 4267 25594 4323 25596
rect 4347 25594 4403 25596
rect 4107 25542 4153 25594
rect 4153 25542 4163 25594
rect 4187 25542 4217 25594
rect 4217 25542 4229 25594
rect 4229 25542 4243 25594
rect 4267 25542 4281 25594
rect 4281 25542 4293 25594
rect 4293 25542 4323 25594
rect 4347 25542 4357 25594
rect 4357 25542 4403 25594
rect 4107 25540 4163 25542
rect 4187 25540 4243 25542
rect 4267 25540 4323 25542
rect 4347 25540 4403 25542
rect 4107 24506 4163 24508
rect 4187 24506 4243 24508
rect 4267 24506 4323 24508
rect 4347 24506 4403 24508
rect 4107 24454 4153 24506
rect 4153 24454 4163 24506
rect 4187 24454 4217 24506
rect 4217 24454 4229 24506
rect 4229 24454 4243 24506
rect 4267 24454 4281 24506
rect 4281 24454 4293 24506
rect 4293 24454 4323 24506
rect 4347 24454 4357 24506
rect 4357 24454 4403 24506
rect 4107 24452 4163 24454
rect 4187 24452 4243 24454
rect 4267 24452 4323 24454
rect 4347 24452 4403 24454
rect 4107 23418 4163 23420
rect 4187 23418 4243 23420
rect 4267 23418 4323 23420
rect 4347 23418 4403 23420
rect 4107 23366 4153 23418
rect 4153 23366 4163 23418
rect 4187 23366 4217 23418
rect 4217 23366 4229 23418
rect 4229 23366 4243 23418
rect 4267 23366 4281 23418
rect 4281 23366 4293 23418
rect 4293 23366 4323 23418
rect 4347 23366 4357 23418
rect 4357 23366 4403 23418
rect 4107 23364 4163 23366
rect 4187 23364 4243 23366
rect 4267 23364 4323 23366
rect 4347 23364 4403 23366
rect 4107 22330 4163 22332
rect 4187 22330 4243 22332
rect 4267 22330 4323 22332
rect 4347 22330 4403 22332
rect 4107 22278 4153 22330
rect 4153 22278 4163 22330
rect 4187 22278 4217 22330
rect 4217 22278 4229 22330
rect 4229 22278 4243 22330
rect 4267 22278 4281 22330
rect 4281 22278 4293 22330
rect 4293 22278 4323 22330
rect 4347 22278 4357 22330
rect 4357 22278 4403 22330
rect 4107 22276 4163 22278
rect 4187 22276 4243 22278
rect 4267 22276 4323 22278
rect 4347 22276 4403 22278
rect 4986 21936 5042 21992
rect 4107 21242 4163 21244
rect 4187 21242 4243 21244
rect 4267 21242 4323 21244
rect 4347 21242 4403 21244
rect 4107 21190 4153 21242
rect 4153 21190 4163 21242
rect 4187 21190 4217 21242
rect 4217 21190 4229 21242
rect 4229 21190 4243 21242
rect 4267 21190 4281 21242
rect 4281 21190 4293 21242
rect 4293 21190 4323 21242
rect 4347 21190 4357 21242
rect 4357 21190 4403 21242
rect 4107 21188 4163 21190
rect 4187 21188 4243 21190
rect 4267 21188 4323 21190
rect 4347 21188 4403 21190
rect 4107 20154 4163 20156
rect 4187 20154 4243 20156
rect 4267 20154 4323 20156
rect 4347 20154 4403 20156
rect 4107 20102 4153 20154
rect 4153 20102 4163 20154
rect 4187 20102 4217 20154
rect 4217 20102 4229 20154
rect 4229 20102 4243 20154
rect 4267 20102 4281 20154
rect 4281 20102 4293 20154
rect 4293 20102 4323 20154
rect 4347 20102 4357 20154
rect 4357 20102 4403 20154
rect 4107 20100 4163 20102
rect 4187 20100 4243 20102
rect 4267 20100 4323 20102
rect 4347 20100 4403 20102
rect 4107 19066 4163 19068
rect 4187 19066 4243 19068
rect 4267 19066 4323 19068
rect 4347 19066 4403 19068
rect 4107 19014 4153 19066
rect 4153 19014 4163 19066
rect 4187 19014 4217 19066
rect 4217 19014 4229 19066
rect 4229 19014 4243 19066
rect 4267 19014 4281 19066
rect 4281 19014 4293 19066
rect 4293 19014 4323 19066
rect 4347 19014 4357 19066
rect 4357 19014 4403 19066
rect 4107 19012 4163 19014
rect 4187 19012 4243 19014
rect 4267 19012 4323 19014
rect 4347 19012 4403 19014
rect 4107 17978 4163 17980
rect 4187 17978 4243 17980
rect 4267 17978 4323 17980
rect 4347 17978 4403 17980
rect 4107 17926 4153 17978
rect 4153 17926 4163 17978
rect 4187 17926 4217 17978
rect 4217 17926 4229 17978
rect 4229 17926 4243 17978
rect 4267 17926 4281 17978
rect 4281 17926 4293 17978
rect 4293 17926 4323 17978
rect 4347 17926 4357 17978
rect 4357 17926 4403 17978
rect 4107 17924 4163 17926
rect 4187 17924 4243 17926
rect 4267 17924 4323 17926
rect 4347 17924 4403 17926
rect 4107 16890 4163 16892
rect 4187 16890 4243 16892
rect 4267 16890 4323 16892
rect 4347 16890 4403 16892
rect 4107 16838 4153 16890
rect 4153 16838 4163 16890
rect 4187 16838 4217 16890
rect 4217 16838 4229 16890
rect 4229 16838 4243 16890
rect 4267 16838 4281 16890
rect 4281 16838 4293 16890
rect 4293 16838 4323 16890
rect 4347 16838 4357 16890
rect 4357 16838 4403 16890
rect 4107 16836 4163 16838
rect 4187 16836 4243 16838
rect 4267 16836 4323 16838
rect 4347 16836 4403 16838
rect 3238 15444 3240 15464
rect 3240 15444 3292 15464
rect 3292 15444 3294 15464
rect 3238 15408 3294 15444
rect 4107 15802 4163 15804
rect 4187 15802 4243 15804
rect 4267 15802 4323 15804
rect 4347 15802 4403 15804
rect 4107 15750 4153 15802
rect 4153 15750 4163 15802
rect 4187 15750 4217 15802
rect 4217 15750 4229 15802
rect 4229 15750 4243 15802
rect 4267 15750 4281 15802
rect 4281 15750 4293 15802
rect 4293 15750 4323 15802
rect 4347 15750 4357 15802
rect 4357 15750 4403 15802
rect 4107 15748 4163 15750
rect 4187 15748 4243 15750
rect 4267 15748 4323 15750
rect 4347 15748 4403 15750
rect 3146 14864 3202 14920
rect 4107 14714 4163 14716
rect 4187 14714 4243 14716
rect 4267 14714 4323 14716
rect 4347 14714 4403 14716
rect 4107 14662 4153 14714
rect 4153 14662 4163 14714
rect 4187 14662 4217 14714
rect 4217 14662 4229 14714
rect 4229 14662 4243 14714
rect 4267 14662 4281 14714
rect 4281 14662 4293 14714
rect 4293 14662 4323 14714
rect 4347 14662 4357 14714
rect 4357 14662 4403 14714
rect 4107 14660 4163 14662
rect 4187 14660 4243 14662
rect 4267 14660 4323 14662
rect 4347 14660 4403 14662
rect 4107 13626 4163 13628
rect 4187 13626 4243 13628
rect 4267 13626 4323 13628
rect 4347 13626 4403 13628
rect 4107 13574 4153 13626
rect 4153 13574 4163 13626
rect 4187 13574 4217 13626
rect 4217 13574 4229 13626
rect 4229 13574 4243 13626
rect 4267 13574 4281 13626
rect 4281 13574 4293 13626
rect 4293 13574 4323 13626
rect 4347 13574 4357 13626
rect 4357 13574 4403 13626
rect 4107 13572 4163 13574
rect 4187 13572 4243 13574
rect 4267 13572 4323 13574
rect 4347 13572 4403 13574
rect 4107 12538 4163 12540
rect 4187 12538 4243 12540
rect 4267 12538 4323 12540
rect 4347 12538 4403 12540
rect 4107 12486 4153 12538
rect 4153 12486 4163 12538
rect 4187 12486 4217 12538
rect 4217 12486 4229 12538
rect 4229 12486 4243 12538
rect 4267 12486 4281 12538
rect 4281 12486 4293 12538
rect 4293 12486 4323 12538
rect 4347 12486 4357 12538
rect 4357 12486 4403 12538
rect 4107 12484 4163 12486
rect 4187 12484 4243 12486
rect 4267 12484 4323 12486
rect 4347 12484 4403 12486
rect 7258 26138 7314 26140
rect 7338 26138 7394 26140
rect 7418 26138 7474 26140
rect 7498 26138 7554 26140
rect 7258 26086 7304 26138
rect 7304 26086 7314 26138
rect 7338 26086 7368 26138
rect 7368 26086 7380 26138
rect 7380 26086 7394 26138
rect 7418 26086 7432 26138
rect 7432 26086 7444 26138
rect 7444 26086 7474 26138
rect 7498 26086 7508 26138
rect 7508 26086 7554 26138
rect 7258 26084 7314 26086
rect 7338 26084 7394 26086
rect 7418 26084 7474 26086
rect 7498 26084 7554 26086
rect 6458 24656 6514 24712
rect 7258 25050 7314 25052
rect 7338 25050 7394 25052
rect 7418 25050 7474 25052
rect 7498 25050 7554 25052
rect 7258 24998 7304 25050
rect 7304 24998 7314 25050
rect 7338 24998 7368 25050
rect 7368 24998 7380 25050
rect 7380 24998 7394 25050
rect 7418 24998 7432 25050
rect 7432 24998 7444 25050
rect 7444 24998 7474 25050
rect 7498 24998 7508 25050
rect 7508 24998 7554 25050
rect 7258 24996 7314 24998
rect 7338 24996 7394 24998
rect 7418 24996 7474 24998
rect 7498 24996 7554 24998
rect 7562 24676 7618 24712
rect 7562 24656 7564 24676
rect 7564 24656 7616 24676
rect 7616 24656 7618 24676
rect 7258 23962 7314 23964
rect 7338 23962 7394 23964
rect 7418 23962 7474 23964
rect 7498 23962 7554 23964
rect 7258 23910 7304 23962
rect 7304 23910 7314 23962
rect 7338 23910 7368 23962
rect 7368 23910 7380 23962
rect 7380 23910 7394 23962
rect 7418 23910 7432 23962
rect 7432 23910 7444 23962
rect 7444 23910 7474 23962
rect 7498 23910 7508 23962
rect 7508 23910 7554 23962
rect 7258 23908 7314 23910
rect 7338 23908 7394 23910
rect 7418 23908 7474 23910
rect 7498 23908 7554 23910
rect 5262 19796 5264 19816
rect 5264 19796 5316 19816
rect 5316 19796 5318 19816
rect 5262 19760 5318 19796
rect 6182 19760 6238 19816
rect 938 4120 994 4176
rect 7258 22874 7314 22876
rect 7338 22874 7394 22876
rect 7418 22874 7474 22876
rect 7498 22874 7554 22876
rect 7258 22822 7304 22874
rect 7304 22822 7314 22874
rect 7338 22822 7368 22874
rect 7368 22822 7380 22874
rect 7380 22822 7394 22874
rect 7418 22822 7432 22874
rect 7432 22822 7444 22874
rect 7444 22822 7474 22874
rect 7498 22822 7508 22874
rect 7508 22822 7554 22874
rect 7258 22820 7314 22822
rect 7338 22820 7394 22822
rect 7418 22820 7474 22822
rect 7498 22820 7554 22822
rect 6918 20848 6974 20904
rect 7258 21786 7314 21788
rect 7338 21786 7394 21788
rect 7418 21786 7474 21788
rect 7498 21786 7554 21788
rect 7258 21734 7304 21786
rect 7304 21734 7314 21786
rect 7338 21734 7368 21786
rect 7368 21734 7380 21786
rect 7380 21734 7394 21786
rect 7418 21734 7432 21786
rect 7432 21734 7444 21786
rect 7444 21734 7474 21786
rect 7498 21734 7508 21786
rect 7508 21734 7554 21786
rect 7258 21732 7314 21734
rect 7338 21732 7394 21734
rect 7418 21732 7474 21734
rect 7498 21732 7554 21734
rect 7194 20868 7250 20904
rect 7194 20848 7196 20868
rect 7196 20848 7248 20868
rect 7248 20848 7250 20868
rect 7258 20698 7314 20700
rect 7338 20698 7394 20700
rect 7418 20698 7474 20700
rect 7498 20698 7554 20700
rect 7258 20646 7304 20698
rect 7304 20646 7314 20698
rect 7338 20646 7368 20698
rect 7368 20646 7380 20698
rect 7380 20646 7394 20698
rect 7418 20646 7432 20698
rect 7432 20646 7444 20698
rect 7444 20646 7474 20698
rect 7498 20646 7508 20698
rect 7508 20646 7554 20698
rect 7258 20644 7314 20646
rect 7338 20644 7394 20646
rect 7418 20644 7474 20646
rect 7498 20644 7554 20646
rect 7258 19610 7314 19612
rect 7338 19610 7394 19612
rect 7418 19610 7474 19612
rect 7498 19610 7554 19612
rect 7258 19558 7304 19610
rect 7304 19558 7314 19610
rect 7338 19558 7368 19610
rect 7368 19558 7380 19610
rect 7380 19558 7394 19610
rect 7418 19558 7432 19610
rect 7432 19558 7444 19610
rect 7444 19558 7474 19610
rect 7498 19558 7508 19610
rect 7508 19558 7554 19610
rect 7258 19556 7314 19558
rect 7338 19556 7394 19558
rect 7418 19556 7474 19558
rect 7498 19556 7554 19558
rect 10409 26682 10465 26684
rect 10489 26682 10545 26684
rect 10569 26682 10625 26684
rect 10649 26682 10705 26684
rect 10409 26630 10455 26682
rect 10455 26630 10465 26682
rect 10489 26630 10519 26682
rect 10519 26630 10531 26682
rect 10531 26630 10545 26682
rect 10569 26630 10583 26682
rect 10583 26630 10595 26682
rect 10595 26630 10625 26682
rect 10649 26630 10659 26682
rect 10659 26630 10705 26682
rect 10409 26628 10465 26630
rect 10489 26628 10545 26630
rect 10569 26628 10625 26630
rect 10649 26628 10705 26630
rect 10966 26424 11022 26480
rect 10409 25594 10465 25596
rect 10489 25594 10545 25596
rect 10569 25594 10625 25596
rect 10649 25594 10705 25596
rect 10409 25542 10455 25594
rect 10455 25542 10465 25594
rect 10489 25542 10519 25594
rect 10519 25542 10531 25594
rect 10531 25542 10545 25594
rect 10569 25542 10583 25594
rect 10583 25542 10595 25594
rect 10595 25542 10625 25594
rect 10649 25542 10659 25594
rect 10659 25542 10705 25594
rect 10409 25540 10465 25542
rect 10489 25540 10545 25542
rect 10569 25540 10625 25542
rect 10649 25540 10705 25542
rect 10409 24506 10465 24508
rect 10489 24506 10545 24508
rect 10569 24506 10625 24508
rect 10649 24506 10705 24508
rect 10409 24454 10455 24506
rect 10455 24454 10465 24506
rect 10489 24454 10519 24506
rect 10519 24454 10531 24506
rect 10531 24454 10545 24506
rect 10569 24454 10583 24506
rect 10583 24454 10595 24506
rect 10595 24454 10625 24506
rect 10649 24454 10659 24506
rect 10659 24454 10705 24506
rect 10409 24452 10465 24454
rect 10489 24452 10545 24454
rect 10569 24452 10625 24454
rect 10649 24452 10705 24454
rect 10409 23418 10465 23420
rect 10489 23418 10545 23420
rect 10569 23418 10625 23420
rect 10649 23418 10705 23420
rect 10409 23366 10455 23418
rect 10455 23366 10465 23418
rect 10489 23366 10519 23418
rect 10519 23366 10531 23418
rect 10531 23366 10545 23418
rect 10569 23366 10583 23418
rect 10583 23366 10595 23418
rect 10595 23366 10625 23418
rect 10649 23366 10659 23418
rect 10659 23366 10705 23418
rect 10409 23364 10465 23366
rect 10489 23364 10545 23366
rect 10569 23364 10625 23366
rect 10649 23364 10705 23366
rect 6918 19216 6974 19272
rect 7258 18522 7314 18524
rect 7338 18522 7394 18524
rect 7418 18522 7474 18524
rect 7498 18522 7554 18524
rect 7258 18470 7304 18522
rect 7304 18470 7314 18522
rect 7338 18470 7368 18522
rect 7368 18470 7380 18522
rect 7380 18470 7394 18522
rect 7418 18470 7432 18522
rect 7432 18470 7444 18522
rect 7444 18470 7474 18522
rect 7498 18470 7508 18522
rect 7508 18470 7554 18522
rect 7258 18468 7314 18470
rect 7338 18468 7394 18470
rect 7418 18468 7474 18470
rect 7498 18468 7554 18470
rect 5906 15428 5962 15464
rect 5906 15408 5908 15428
rect 5908 15408 5960 15428
rect 5960 15408 5962 15428
rect 4107 11450 4163 11452
rect 4187 11450 4243 11452
rect 4267 11450 4323 11452
rect 4347 11450 4403 11452
rect 4107 11398 4153 11450
rect 4153 11398 4163 11450
rect 4187 11398 4217 11450
rect 4217 11398 4229 11450
rect 4229 11398 4243 11450
rect 4267 11398 4281 11450
rect 4281 11398 4293 11450
rect 4293 11398 4323 11450
rect 4347 11398 4357 11450
rect 4357 11398 4403 11450
rect 4107 11396 4163 11398
rect 4187 11396 4243 11398
rect 4267 11396 4323 11398
rect 4347 11396 4403 11398
rect 4107 10362 4163 10364
rect 4187 10362 4243 10364
rect 4267 10362 4323 10364
rect 4347 10362 4403 10364
rect 4107 10310 4153 10362
rect 4153 10310 4163 10362
rect 4187 10310 4217 10362
rect 4217 10310 4229 10362
rect 4229 10310 4243 10362
rect 4267 10310 4281 10362
rect 4281 10310 4293 10362
rect 4293 10310 4323 10362
rect 4347 10310 4357 10362
rect 4357 10310 4403 10362
rect 4107 10308 4163 10310
rect 4187 10308 4243 10310
rect 4267 10308 4323 10310
rect 4347 10308 4403 10310
rect 5630 10648 5686 10704
rect 3882 9596 3884 9616
rect 3884 9596 3936 9616
rect 3936 9596 3938 9616
rect 3882 9560 3938 9596
rect 4107 9274 4163 9276
rect 4187 9274 4243 9276
rect 4267 9274 4323 9276
rect 4347 9274 4403 9276
rect 4107 9222 4153 9274
rect 4153 9222 4163 9274
rect 4187 9222 4217 9274
rect 4217 9222 4229 9274
rect 4229 9222 4243 9274
rect 4267 9222 4281 9274
rect 4281 9222 4293 9274
rect 4293 9222 4323 9274
rect 4347 9222 4357 9274
rect 4357 9222 4403 9274
rect 4107 9220 4163 9222
rect 4187 9220 4243 9222
rect 4267 9220 4323 9222
rect 4347 9220 4403 9222
rect 4802 9580 4858 9616
rect 4802 9560 4804 9580
rect 4804 9560 4856 9580
rect 4856 9560 4858 9580
rect 4107 8186 4163 8188
rect 4187 8186 4243 8188
rect 4267 8186 4323 8188
rect 4347 8186 4403 8188
rect 4107 8134 4153 8186
rect 4153 8134 4163 8186
rect 4187 8134 4217 8186
rect 4217 8134 4229 8186
rect 4229 8134 4243 8186
rect 4267 8134 4281 8186
rect 4281 8134 4293 8186
rect 4293 8134 4323 8186
rect 4347 8134 4357 8186
rect 4357 8134 4403 8186
rect 4107 8132 4163 8134
rect 4187 8132 4243 8134
rect 4267 8132 4323 8134
rect 4347 8132 4403 8134
rect 4107 7098 4163 7100
rect 4187 7098 4243 7100
rect 4267 7098 4323 7100
rect 4347 7098 4403 7100
rect 4107 7046 4153 7098
rect 4153 7046 4163 7098
rect 4187 7046 4217 7098
rect 4217 7046 4229 7098
rect 4229 7046 4243 7098
rect 4267 7046 4281 7098
rect 4281 7046 4293 7098
rect 4293 7046 4323 7098
rect 4347 7046 4357 7098
rect 4357 7046 4403 7098
rect 4107 7044 4163 7046
rect 4187 7044 4243 7046
rect 4267 7044 4323 7046
rect 4347 7044 4403 7046
rect 4107 6010 4163 6012
rect 4187 6010 4243 6012
rect 4267 6010 4323 6012
rect 4347 6010 4403 6012
rect 4107 5958 4153 6010
rect 4153 5958 4163 6010
rect 4187 5958 4217 6010
rect 4217 5958 4229 6010
rect 4229 5958 4243 6010
rect 4267 5958 4281 6010
rect 4281 5958 4293 6010
rect 4293 5958 4323 6010
rect 4347 5958 4357 6010
rect 4357 5958 4403 6010
rect 4107 5956 4163 5958
rect 4187 5956 4243 5958
rect 4267 5956 4323 5958
rect 4347 5956 4403 5958
rect 4107 4922 4163 4924
rect 4187 4922 4243 4924
rect 4267 4922 4323 4924
rect 4347 4922 4403 4924
rect 4107 4870 4153 4922
rect 4153 4870 4163 4922
rect 4187 4870 4217 4922
rect 4217 4870 4229 4922
rect 4229 4870 4243 4922
rect 4267 4870 4281 4922
rect 4281 4870 4293 4922
rect 4293 4870 4323 4922
rect 4347 4870 4357 4922
rect 4357 4870 4403 4922
rect 4107 4868 4163 4870
rect 4187 4868 4243 4870
rect 4267 4868 4323 4870
rect 4347 4868 4403 4870
rect 4107 3834 4163 3836
rect 4187 3834 4243 3836
rect 4267 3834 4323 3836
rect 4347 3834 4403 3836
rect 4107 3782 4153 3834
rect 4153 3782 4163 3834
rect 4187 3782 4217 3834
rect 4217 3782 4229 3834
rect 4229 3782 4243 3834
rect 4267 3782 4281 3834
rect 4281 3782 4293 3834
rect 4293 3782 4323 3834
rect 4347 3782 4357 3834
rect 4357 3782 4403 3834
rect 4107 3780 4163 3782
rect 4187 3780 4243 3782
rect 4267 3780 4323 3782
rect 4347 3780 4403 3782
rect 4107 2746 4163 2748
rect 4187 2746 4243 2748
rect 4267 2746 4323 2748
rect 4347 2746 4403 2748
rect 4107 2694 4153 2746
rect 4153 2694 4163 2746
rect 4187 2694 4217 2746
rect 4217 2694 4229 2746
rect 4229 2694 4243 2746
rect 4267 2694 4281 2746
rect 4281 2694 4293 2746
rect 4293 2694 4323 2746
rect 4347 2694 4357 2746
rect 4357 2694 4403 2746
rect 4107 2692 4163 2694
rect 4187 2692 4243 2694
rect 4267 2692 4323 2694
rect 4347 2692 4403 2694
rect 7258 17434 7314 17436
rect 7338 17434 7394 17436
rect 7418 17434 7474 17436
rect 7498 17434 7554 17436
rect 7258 17382 7304 17434
rect 7304 17382 7314 17434
rect 7338 17382 7368 17434
rect 7368 17382 7380 17434
rect 7380 17382 7394 17434
rect 7418 17382 7432 17434
rect 7432 17382 7444 17434
rect 7444 17382 7474 17434
rect 7498 17382 7508 17434
rect 7508 17382 7554 17434
rect 7258 17380 7314 17382
rect 7338 17380 7394 17382
rect 7418 17380 7474 17382
rect 7498 17380 7554 17382
rect 7258 16346 7314 16348
rect 7338 16346 7394 16348
rect 7418 16346 7474 16348
rect 7498 16346 7554 16348
rect 7258 16294 7304 16346
rect 7304 16294 7314 16346
rect 7338 16294 7368 16346
rect 7368 16294 7380 16346
rect 7380 16294 7394 16346
rect 7418 16294 7432 16346
rect 7432 16294 7444 16346
rect 7444 16294 7474 16346
rect 7498 16294 7508 16346
rect 7508 16294 7554 16346
rect 7258 16292 7314 16294
rect 7338 16292 7394 16294
rect 7418 16292 7474 16294
rect 7498 16292 7554 16294
rect 7258 15258 7314 15260
rect 7338 15258 7394 15260
rect 7418 15258 7474 15260
rect 7498 15258 7554 15260
rect 7258 15206 7304 15258
rect 7304 15206 7314 15258
rect 7338 15206 7368 15258
rect 7368 15206 7380 15258
rect 7380 15206 7394 15258
rect 7418 15206 7432 15258
rect 7432 15206 7444 15258
rect 7444 15206 7474 15258
rect 7498 15206 7508 15258
rect 7508 15206 7554 15258
rect 7258 15204 7314 15206
rect 7338 15204 7394 15206
rect 7418 15204 7474 15206
rect 7498 15204 7554 15206
rect 7258 14170 7314 14172
rect 7338 14170 7394 14172
rect 7418 14170 7474 14172
rect 7498 14170 7554 14172
rect 7258 14118 7304 14170
rect 7304 14118 7314 14170
rect 7338 14118 7368 14170
rect 7368 14118 7380 14170
rect 7380 14118 7394 14170
rect 7418 14118 7432 14170
rect 7432 14118 7444 14170
rect 7444 14118 7474 14170
rect 7498 14118 7508 14170
rect 7508 14118 7554 14170
rect 7258 14116 7314 14118
rect 7338 14116 7394 14118
rect 7418 14116 7474 14118
rect 7498 14116 7554 14118
rect 7258 13082 7314 13084
rect 7338 13082 7394 13084
rect 7418 13082 7474 13084
rect 7498 13082 7554 13084
rect 7258 13030 7304 13082
rect 7304 13030 7314 13082
rect 7338 13030 7368 13082
rect 7368 13030 7380 13082
rect 7380 13030 7394 13082
rect 7418 13030 7432 13082
rect 7432 13030 7444 13082
rect 7444 13030 7474 13082
rect 7498 13030 7508 13082
rect 7508 13030 7554 13082
rect 7258 13028 7314 13030
rect 7338 13028 7394 13030
rect 7418 13028 7474 13030
rect 7498 13028 7554 13030
rect 6734 10648 6790 10704
rect 7258 11994 7314 11996
rect 7338 11994 7394 11996
rect 7418 11994 7474 11996
rect 7498 11994 7554 11996
rect 7258 11942 7304 11994
rect 7304 11942 7314 11994
rect 7338 11942 7368 11994
rect 7368 11942 7380 11994
rect 7380 11942 7394 11994
rect 7418 11942 7432 11994
rect 7432 11942 7444 11994
rect 7444 11942 7474 11994
rect 7498 11942 7508 11994
rect 7508 11942 7554 11994
rect 7258 11940 7314 11942
rect 7338 11940 7394 11942
rect 7418 11940 7474 11942
rect 7498 11940 7554 11942
rect 7258 10906 7314 10908
rect 7338 10906 7394 10908
rect 7418 10906 7474 10908
rect 7498 10906 7554 10908
rect 7258 10854 7304 10906
rect 7304 10854 7314 10906
rect 7338 10854 7368 10906
rect 7368 10854 7380 10906
rect 7380 10854 7394 10906
rect 7418 10854 7432 10906
rect 7432 10854 7444 10906
rect 7444 10854 7474 10906
rect 7498 10854 7508 10906
rect 7508 10854 7554 10906
rect 7258 10852 7314 10854
rect 7338 10852 7394 10854
rect 7418 10852 7474 10854
rect 7498 10852 7554 10854
rect 6458 8472 6514 8528
rect 7258 9818 7314 9820
rect 7338 9818 7394 9820
rect 7418 9818 7474 9820
rect 7498 9818 7554 9820
rect 7258 9766 7304 9818
rect 7304 9766 7314 9818
rect 7338 9766 7368 9818
rect 7368 9766 7380 9818
rect 7380 9766 7394 9818
rect 7418 9766 7432 9818
rect 7432 9766 7444 9818
rect 7444 9766 7474 9818
rect 7498 9766 7508 9818
rect 7508 9766 7554 9818
rect 7258 9764 7314 9766
rect 7338 9764 7394 9766
rect 7418 9764 7474 9766
rect 7498 9764 7554 9766
rect 7258 8730 7314 8732
rect 7338 8730 7394 8732
rect 7418 8730 7474 8732
rect 7498 8730 7554 8732
rect 7258 8678 7304 8730
rect 7304 8678 7314 8730
rect 7338 8678 7368 8730
rect 7368 8678 7380 8730
rect 7380 8678 7394 8730
rect 7418 8678 7432 8730
rect 7432 8678 7444 8730
rect 7444 8678 7474 8730
rect 7498 8678 7508 8730
rect 7508 8678 7554 8730
rect 7258 8676 7314 8678
rect 7338 8676 7394 8678
rect 7418 8676 7474 8678
rect 7498 8676 7554 8678
rect 7258 7642 7314 7644
rect 7338 7642 7394 7644
rect 7418 7642 7474 7644
rect 7498 7642 7554 7644
rect 7258 7590 7304 7642
rect 7304 7590 7314 7642
rect 7338 7590 7368 7642
rect 7368 7590 7380 7642
rect 7380 7590 7394 7642
rect 7418 7590 7432 7642
rect 7432 7590 7444 7642
rect 7444 7590 7474 7642
rect 7498 7590 7508 7642
rect 7508 7590 7554 7642
rect 7258 7588 7314 7590
rect 7338 7588 7394 7590
rect 7418 7588 7474 7590
rect 7498 7588 7554 7590
rect 7258 6554 7314 6556
rect 7338 6554 7394 6556
rect 7418 6554 7474 6556
rect 7498 6554 7554 6556
rect 7258 6502 7304 6554
rect 7304 6502 7314 6554
rect 7338 6502 7368 6554
rect 7368 6502 7380 6554
rect 7380 6502 7394 6554
rect 7418 6502 7432 6554
rect 7432 6502 7444 6554
rect 7444 6502 7474 6554
rect 7498 6502 7508 6554
rect 7508 6502 7554 6554
rect 7258 6500 7314 6502
rect 7338 6500 7394 6502
rect 7418 6500 7474 6502
rect 7498 6500 7554 6502
rect 10409 22330 10465 22332
rect 10489 22330 10545 22332
rect 10569 22330 10625 22332
rect 10649 22330 10705 22332
rect 10409 22278 10455 22330
rect 10455 22278 10465 22330
rect 10489 22278 10519 22330
rect 10519 22278 10531 22330
rect 10531 22278 10545 22330
rect 10569 22278 10583 22330
rect 10583 22278 10595 22330
rect 10595 22278 10625 22330
rect 10649 22278 10659 22330
rect 10659 22278 10705 22330
rect 10409 22276 10465 22278
rect 10489 22276 10545 22278
rect 10569 22276 10625 22278
rect 10649 22276 10705 22278
rect 10409 21242 10465 21244
rect 10489 21242 10545 21244
rect 10569 21242 10625 21244
rect 10649 21242 10705 21244
rect 10409 21190 10455 21242
rect 10455 21190 10465 21242
rect 10489 21190 10519 21242
rect 10519 21190 10531 21242
rect 10531 21190 10545 21242
rect 10569 21190 10583 21242
rect 10583 21190 10595 21242
rect 10595 21190 10625 21242
rect 10649 21190 10659 21242
rect 10659 21190 10705 21242
rect 10409 21188 10465 21190
rect 10489 21188 10545 21190
rect 10569 21188 10625 21190
rect 10649 21188 10705 21190
rect 10409 20154 10465 20156
rect 10489 20154 10545 20156
rect 10569 20154 10625 20156
rect 10649 20154 10705 20156
rect 10409 20102 10455 20154
rect 10455 20102 10465 20154
rect 10489 20102 10519 20154
rect 10519 20102 10531 20154
rect 10531 20102 10545 20154
rect 10569 20102 10583 20154
rect 10583 20102 10595 20154
rect 10595 20102 10625 20154
rect 10649 20102 10659 20154
rect 10659 20102 10705 20154
rect 10409 20100 10465 20102
rect 10489 20100 10545 20102
rect 10569 20100 10625 20102
rect 10649 20100 10705 20102
rect 10409 19066 10465 19068
rect 10489 19066 10545 19068
rect 10569 19066 10625 19068
rect 10649 19066 10705 19068
rect 10409 19014 10455 19066
rect 10455 19014 10465 19066
rect 10489 19014 10519 19066
rect 10519 19014 10531 19066
rect 10531 19014 10545 19066
rect 10569 19014 10583 19066
rect 10583 19014 10595 19066
rect 10595 19014 10625 19066
rect 10649 19014 10659 19066
rect 10659 19014 10705 19066
rect 10409 19012 10465 19014
rect 10489 19012 10545 19014
rect 10569 19012 10625 19014
rect 10649 19012 10705 19014
rect 10409 17978 10465 17980
rect 10489 17978 10545 17980
rect 10569 17978 10625 17980
rect 10649 17978 10705 17980
rect 10409 17926 10455 17978
rect 10455 17926 10465 17978
rect 10489 17926 10519 17978
rect 10519 17926 10531 17978
rect 10531 17926 10545 17978
rect 10569 17926 10583 17978
rect 10583 17926 10595 17978
rect 10595 17926 10625 17978
rect 10649 17926 10659 17978
rect 10659 17926 10705 17978
rect 10409 17924 10465 17926
rect 10489 17924 10545 17926
rect 10569 17924 10625 17926
rect 10649 17924 10705 17926
rect 10409 16890 10465 16892
rect 10489 16890 10545 16892
rect 10569 16890 10625 16892
rect 10649 16890 10705 16892
rect 10409 16838 10455 16890
rect 10455 16838 10465 16890
rect 10489 16838 10519 16890
rect 10519 16838 10531 16890
rect 10531 16838 10545 16890
rect 10569 16838 10583 16890
rect 10583 16838 10595 16890
rect 10595 16838 10625 16890
rect 10649 16838 10659 16890
rect 10659 16838 10705 16890
rect 10409 16836 10465 16838
rect 10489 16836 10545 16838
rect 10569 16836 10625 16838
rect 10649 16836 10705 16838
rect 10409 15802 10465 15804
rect 10489 15802 10545 15804
rect 10569 15802 10625 15804
rect 10649 15802 10705 15804
rect 10409 15750 10455 15802
rect 10455 15750 10465 15802
rect 10489 15750 10519 15802
rect 10519 15750 10531 15802
rect 10531 15750 10545 15802
rect 10569 15750 10583 15802
rect 10583 15750 10595 15802
rect 10595 15750 10625 15802
rect 10649 15750 10659 15802
rect 10659 15750 10705 15802
rect 10409 15748 10465 15750
rect 10489 15748 10545 15750
rect 10569 15748 10625 15750
rect 10649 15748 10705 15750
rect 12898 26424 12954 26480
rect 13560 26138 13616 26140
rect 13640 26138 13696 26140
rect 13720 26138 13776 26140
rect 13800 26138 13856 26140
rect 13560 26086 13606 26138
rect 13606 26086 13616 26138
rect 13640 26086 13670 26138
rect 13670 26086 13682 26138
rect 13682 26086 13696 26138
rect 13720 26086 13734 26138
rect 13734 26086 13746 26138
rect 13746 26086 13776 26138
rect 13800 26086 13810 26138
rect 13810 26086 13856 26138
rect 13560 26084 13616 26086
rect 13640 26084 13696 26086
rect 13720 26084 13776 26086
rect 13800 26084 13856 26086
rect 14830 26424 14886 26480
rect 13560 25050 13616 25052
rect 13640 25050 13696 25052
rect 13720 25050 13776 25052
rect 13800 25050 13856 25052
rect 13560 24998 13606 25050
rect 13606 24998 13616 25050
rect 13640 24998 13670 25050
rect 13670 24998 13682 25050
rect 13682 24998 13696 25050
rect 13720 24998 13734 25050
rect 13734 24998 13746 25050
rect 13746 24998 13776 25050
rect 13800 24998 13810 25050
rect 13810 24998 13856 25050
rect 13560 24996 13616 24998
rect 13640 24996 13696 24998
rect 13720 24996 13776 24998
rect 13800 24996 13856 24998
rect 13560 23962 13616 23964
rect 13640 23962 13696 23964
rect 13720 23962 13776 23964
rect 13800 23962 13856 23964
rect 13560 23910 13606 23962
rect 13606 23910 13616 23962
rect 13640 23910 13670 23962
rect 13670 23910 13682 23962
rect 13682 23910 13696 23962
rect 13720 23910 13734 23962
rect 13734 23910 13746 23962
rect 13746 23910 13776 23962
rect 13800 23910 13810 23962
rect 13810 23910 13856 23962
rect 13560 23908 13616 23910
rect 13640 23908 13696 23910
rect 13720 23908 13776 23910
rect 13800 23908 13856 23910
rect 9954 15000 10010 15056
rect 10409 14714 10465 14716
rect 10489 14714 10545 14716
rect 10569 14714 10625 14716
rect 10649 14714 10705 14716
rect 10409 14662 10455 14714
rect 10455 14662 10465 14714
rect 10489 14662 10519 14714
rect 10519 14662 10531 14714
rect 10531 14662 10545 14714
rect 10569 14662 10583 14714
rect 10583 14662 10595 14714
rect 10595 14662 10625 14714
rect 10649 14662 10659 14714
rect 10659 14662 10705 14714
rect 10409 14660 10465 14662
rect 10489 14660 10545 14662
rect 10569 14660 10625 14662
rect 10649 14660 10705 14662
rect 10409 13626 10465 13628
rect 10489 13626 10545 13628
rect 10569 13626 10625 13628
rect 10649 13626 10705 13628
rect 10409 13574 10455 13626
rect 10455 13574 10465 13626
rect 10489 13574 10519 13626
rect 10519 13574 10531 13626
rect 10531 13574 10545 13626
rect 10569 13574 10583 13626
rect 10583 13574 10595 13626
rect 10595 13574 10625 13626
rect 10649 13574 10659 13626
rect 10659 13574 10705 13626
rect 10409 13572 10465 13574
rect 10489 13572 10545 13574
rect 10569 13572 10625 13574
rect 10649 13572 10705 13574
rect 10409 12538 10465 12540
rect 10489 12538 10545 12540
rect 10569 12538 10625 12540
rect 10649 12538 10705 12540
rect 10409 12486 10455 12538
rect 10455 12486 10465 12538
rect 10489 12486 10519 12538
rect 10519 12486 10531 12538
rect 10531 12486 10545 12538
rect 10569 12486 10583 12538
rect 10583 12486 10595 12538
rect 10595 12486 10625 12538
rect 10649 12486 10659 12538
rect 10659 12486 10705 12538
rect 10409 12484 10465 12486
rect 10489 12484 10545 12486
rect 10569 12484 10625 12486
rect 10649 12484 10705 12486
rect 8390 8472 8446 8528
rect 7258 5466 7314 5468
rect 7338 5466 7394 5468
rect 7418 5466 7474 5468
rect 7498 5466 7554 5468
rect 7258 5414 7304 5466
rect 7304 5414 7314 5466
rect 7338 5414 7368 5466
rect 7368 5414 7380 5466
rect 7380 5414 7394 5466
rect 7418 5414 7432 5466
rect 7432 5414 7444 5466
rect 7444 5414 7474 5466
rect 7498 5414 7508 5466
rect 7508 5414 7554 5466
rect 7258 5412 7314 5414
rect 7338 5412 7394 5414
rect 7418 5412 7474 5414
rect 7498 5412 7554 5414
rect 7258 4378 7314 4380
rect 7338 4378 7394 4380
rect 7418 4378 7474 4380
rect 7498 4378 7554 4380
rect 7258 4326 7304 4378
rect 7304 4326 7314 4378
rect 7338 4326 7368 4378
rect 7368 4326 7380 4378
rect 7380 4326 7394 4378
rect 7418 4326 7432 4378
rect 7432 4326 7444 4378
rect 7444 4326 7474 4378
rect 7498 4326 7508 4378
rect 7508 4326 7554 4378
rect 7258 4324 7314 4326
rect 7338 4324 7394 4326
rect 7418 4324 7474 4326
rect 7498 4324 7554 4326
rect 10409 11450 10465 11452
rect 10489 11450 10545 11452
rect 10569 11450 10625 11452
rect 10649 11450 10705 11452
rect 10409 11398 10455 11450
rect 10455 11398 10465 11450
rect 10489 11398 10519 11450
rect 10519 11398 10531 11450
rect 10531 11398 10545 11450
rect 10569 11398 10583 11450
rect 10583 11398 10595 11450
rect 10595 11398 10625 11450
rect 10649 11398 10659 11450
rect 10659 11398 10705 11450
rect 10409 11396 10465 11398
rect 10489 11396 10545 11398
rect 10569 11396 10625 11398
rect 10649 11396 10705 11398
rect 9862 10512 9918 10568
rect 10690 10512 10746 10568
rect 10409 10362 10465 10364
rect 10489 10362 10545 10364
rect 10569 10362 10625 10364
rect 10649 10362 10705 10364
rect 10409 10310 10455 10362
rect 10455 10310 10465 10362
rect 10489 10310 10519 10362
rect 10519 10310 10531 10362
rect 10531 10310 10545 10362
rect 10569 10310 10583 10362
rect 10583 10310 10595 10362
rect 10595 10310 10625 10362
rect 10649 10310 10659 10362
rect 10659 10310 10705 10362
rect 10409 10308 10465 10310
rect 10489 10308 10545 10310
rect 10569 10308 10625 10310
rect 10649 10308 10705 10310
rect 10409 9274 10465 9276
rect 10489 9274 10545 9276
rect 10569 9274 10625 9276
rect 10649 9274 10705 9276
rect 10409 9222 10455 9274
rect 10455 9222 10465 9274
rect 10489 9222 10519 9274
rect 10519 9222 10531 9274
rect 10531 9222 10545 9274
rect 10569 9222 10583 9274
rect 10583 9222 10595 9274
rect 10595 9222 10625 9274
rect 10649 9222 10659 9274
rect 10659 9222 10705 9274
rect 10409 9220 10465 9222
rect 10489 9220 10545 9222
rect 10569 9220 10625 9222
rect 10649 9220 10705 9222
rect 10409 8186 10465 8188
rect 10489 8186 10545 8188
rect 10569 8186 10625 8188
rect 10649 8186 10705 8188
rect 10409 8134 10455 8186
rect 10455 8134 10465 8186
rect 10489 8134 10519 8186
rect 10519 8134 10531 8186
rect 10531 8134 10545 8186
rect 10569 8134 10583 8186
rect 10583 8134 10595 8186
rect 10595 8134 10625 8186
rect 10649 8134 10659 8186
rect 10659 8134 10705 8186
rect 10409 8132 10465 8134
rect 10489 8132 10545 8134
rect 10569 8132 10625 8134
rect 10649 8132 10705 8134
rect 10409 7098 10465 7100
rect 10489 7098 10545 7100
rect 10569 7098 10625 7100
rect 10649 7098 10705 7100
rect 10409 7046 10455 7098
rect 10455 7046 10465 7098
rect 10489 7046 10519 7098
rect 10519 7046 10531 7098
rect 10531 7046 10545 7098
rect 10569 7046 10583 7098
rect 10583 7046 10595 7098
rect 10595 7046 10625 7098
rect 10649 7046 10659 7098
rect 10659 7046 10705 7098
rect 10409 7044 10465 7046
rect 10489 7044 10545 7046
rect 10569 7044 10625 7046
rect 10649 7044 10705 7046
rect 12714 17720 12770 17776
rect 13560 22874 13616 22876
rect 13640 22874 13696 22876
rect 13720 22874 13776 22876
rect 13800 22874 13856 22876
rect 13560 22822 13606 22874
rect 13606 22822 13616 22874
rect 13640 22822 13670 22874
rect 13670 22822 13682 22874
rect 13682 22822 13696 22874
rect 13720 22822 13734 22874
rect 13734 22822 13746 22874
rect 13746 22822 13776 22874
rect 13800 22822 13810 22874
rect 13810 22822 13856 22874
rect 13560 22820 13616 22822
rect 13640 22820 13696 22822
rect 13720 22820 13776 22822
rect 13800 22820 13856 22822
rect 13560 21786 13616 21788
rect 13640 21786 13696 21788
rect 13720 21786 13776 21788
rect 13800 21786 13856 21788
rect 13560 21734 13606 21786
rect 13606 21734 13616 21786
rect 13640 21734 13670 21786
rect 13670 21734 13682 21786
rect 13682 21734 13696 21786
rect 13720 21734 13734 21786
rect 13734 21734 13746 21786
rect 13746 21734 13776 21786
rect 13800 21734 13810 21786
rect 13810 21734 13856 21786
rect 13560 21732 13616 21734
rect 13640 21732 13696 21734
rect 13720 21732 13776 21734
rect 13800 21732 13856 21734
rect 13560 20698 13616 20700
rect 13640 20698 13696 20700
rect 13720 20698 13776 20700
rect 13800 20698 13856 20700
rect 13560 20646 13606 20698
rect 13606 20646 13616 20698
rect 13640 20646 13670 20698
rect 13670 20646 13682 20698
rect 13682 20646 13696 20698
rect 13720 20646 13734 20698
rect 13734 20646 13746 20698
rect 13746 20646 13776 20698
rect 13800 20646 13810 20698
rect 13810 20646 13856 20698
rect 13560 20644 13616 20646
rect 13640 20644 13696 20646
rect 13720 20644 13776 20646
rect 13800 20644 13856 20646
rect 13560 19610 13616 19612
rect 13640 19610 13696 19612
rect 13720 19610 13776 19612
rect 13800 19610 13856 19612
rect 13560 19558 13606 19610
rect 13606 19558 13616 19610
rect 13640 19558 13670 19610
rect 13670 19558 13682 19610
rect 13682 19558 13696 19610
rect 13720 19558 13734 19610
rect 13734 19558 13746 19610
rect 13746 19558 13776 19610
rect 13800 19558 13810 19610
rect 13810 19558 13856 19610
rect 13560 19556 13616 19558
rect 13640 19556 13696 19558
rect 13720 19556 13776 19558
rect 13800 19556 13856 19558
rect 13560 18522 13616 18524
rect 13640 18522 13696 18524
rect 13720 18522 13776 18524
rect 13800 18522 13856 18524
rect 13560 18470 13606 18522
rect 13606 18470 13616 18522
rect 13640 18470 13670 18522
rect 13670 18470 13682 18522
rect 13682 18470 13696 18522
rect 13720 18470 13734 18522
rect 13734 18470 13746 18522
rect 13746 18470 13776 18522
rect 13800 18470 13810 18522
rect 13810 18470 13856 18522
rect 13560 18468 13616 18470
rect 13640 18468 13696 18470
rect 13720 18468 13776 18470
rect 13800 18468 13856 18470
rect 13560 17434 13616 17436
rect 13640 17434 13696 17436
rect 13720 17434 13776 17436
rect 13800 17434 13856 17436
rect 13560 17382 13606 17434
rect 13606 17382 13616 17434
rect 13640 17382 13670 17434
rect 13670 17382 13682 17434
rect 13682 17382 13696 17434
rect 13720 17382 13734 17434
rect 13734 17382 13746 17434
rect 13746 17382 13776 17434
rect 13800 17382 13810 17434
rect 13810 17382 13856 17434
rect 13560 17380 13616 17382
rect 13640 17380 13696 17382
rect 13720 17380 13776 17382
rect 13800 17380 13856 17382
rect 13560 16346 13616 16348
rect 13640 16346 13696 16348
rect 13720 16346 13776 16348
rect 13800 16346 13856 16348
rect 13560 16294 13606 16346
rect 13606 16294 13616 16346
rect 13640 16294 13670 16346
rect 13670 16294 13682 16346
rect 13682 16294 13696 16346
rect 13720 16294 13734 16346
rect 13734 16294 13746 16346
rect 13746 16294 13776 16346
rect 13800 16294 13810 16346
rect 13810 16294 13856 16346
rect 13560 16292 13616 16294
rect 13640 16292 13696 16294
rect 13720 16292 13776 16294
rect 13800 16292 13856 16294
rect 13560 15258 13616 15260
rect 13640 15258 13696 15260
rect 13720 15258 13776 15260
rect 13800 15258 13856 15260
rect 13560 15206 13606 15258
rect 13606 15206 13616 15258
rect 13640 15206 13670 15258
rect 13670 15206 13682 15258
rect 13682 15206 13696 15258
rect 13720 15206 13734 15258
rect 13734 15206 13746 15258
rect 13746 15206 13776 15258
rect 13800 15206 13810 15258
rect 13810 15206 13856 15258
rect 13560 15204 13616 15206
rect 13640 15204 13696 15206
rect 13720 15204 13776 15206
rect 13800 15204 13856 15206
rect 7258 3290 7314 3292
rect 7338 3290 7394 3292
rect 7418 3290 7474 3292
rect 7498 3290 7554 3292
rect 7258 3238 7304 3290
rect 7304 3238 7314 3290
rect 7338 3238 7368 3290
rect 7368 3238 7380 3290
rect 7380 3238 7394 3290
rect 7418 3238 7432 3290
rect 7432 3238 7444 3290
rect 7444 3238 7474 3290
rect 7498 3238 7508 3290
rect 7508 3238 7554 3290
rect 7258 3236 7314 3238
rect 7338 3236 7394 3238
rect 7418 3236 7474 3238
rect 7498 3236 7554 3238
rect 10409 6010 10465 6012
rect 10489 6010 10545 6012
rect 10569 6010 10625 6012
rect 10649 6010 10705 6012
rect 10409 5958 10455 6010
rect 10455 5958 10465 6010
rect 10489 5958 10519 6010
rect 10519 5958 10531 6010
rect 10531 5958 10545 6010
rect 10569 5958 10583 6010
rect 10583 5958 10595 6010
rect 10595 5958 10625 6010
rect 10649 5958 10659 6010
rect 10659 5958 10705 6010
rect 10409 5956 10465 5958
rect 10489 5956 10545 5958
rect 10569 5956 10625 5958
rect 10649 5956 10705 5958
rect 10409 4922 10465 4924
rect 10489 4922 10545 4924
rect 10569 4922 10625 4924
rect 10649 4922 10705 4924
rect 10409 4870 10455 4922
rect 10455 4870 10465 4922
rect 10489 4870 10519 4922
rect 10519 4870 10531 4922
rect 10531 4870 10545 4922
rect 10569 4870 10583 4922
rect 10583 4870 10595 4922
rect 10595 4870 10625 4922
rect 10649 4870 10659 4922
rect 10659 4870 10705 4922
rect 10409 4868 10465 4870
rect 10489 4868 10545 4870
rect 10569 4868 10625 4870
rect 10649 4868 10705 4870
rect 10409 3834 10465 3836
rect 10489 3834 10545 3836
rect 10569 3834 10625 3836
rect 10649 3834 10705 3836
rect 10409 3782 10455 3834
rect 10455 3782 10465 3834
rect 10489 3782 10519 3834
rect 10519 3782 10531 3834
rect 10531 3782 10545 3834
rect 10569 3782 10583 3834
rect 10583 3782 10595 3834
rect 10595 3782 10625 3834
rect 10649 3782 10659 3834
rect 10659 3782 10705 3834
rect 10409 3780 10465 3782
rect 10489 3780 10545 3782
rect 10569 3780 10625 3782
rect 10649 3780 10705 3782
rect 13560 14170 13616 14172
rect 13640 14170 13696 14172
rect 13720 14170 13776 14172
rect 13800 14170 13856 14172
rect 13560 14118 13606 14170
rect 13606 14118 13616 14170
rect 13640 14118 13670 14170
rect 13670 14118 13682 14170
rect 13682 14118 13696 14170
rect 13720 14118 13734 14170
rect 13734 14118 13746 14170
rect 13746 14118 13776 14170
rect 13800 14118 13810 14170
rect 13810 14118 13856 14170
rect 13560 14116 13616 14118
rect 13640 14116 13696 14118
rect 13720 14116 13776 14118
rect 13800 14116 13856 14118
rect 14462 19216 14518 19272
rect 14646 18808 14702 18864
rect 13560 13082 13616 13084
rect 13640 13082 13696 13084
rect 13720 13082 13776 13084
rect 13800 13082 13856 13084
rect 13560 13030 13606 13082
rect 13606 13030 13616 13082
rect 13640 13030 13670 13082
rect 13670 13030 13682 13082
rect 13682 13030 13696 13082
rect 13720 13030 13734 13082
rect 13734 13030 13746 13082
rect 13746 13030 13776 13082
rect 13800 13030 13810 13082
rect 13810 13030 13856 13082
rect 13560 13028 13616 13030
rect 13640 13028 13696 13030
rect 13720 13028 13776 13030
rect 13800 13028 13856 13030
rect 13910 12824 13966 12880
rect 13560 11994 13616 11996
rect 13640 11994 13696 11996
rect 13720 11994 13776 11996
rect 13800 11994 13856 11996
rect 13560 11942 13606 11994
rect 13606 11942 13616 11994
rect 13640 11942 13670 11994
rect 13670 11942 13682 11994
rect 13682 11942 13696 11994
rect 13720 11942 13734 11994
rect 13734 11942 13746 11994
rect 13746 11942 13776 11994
rect 13800 11942 13810 11994
rect 13810 11942 13856 11994
rect 13560 11940 13616 11942
rect 13640 11940 13696 11942
rect 13720 11940 13776 11942
rect 13800 11940 13856 11942
rect 13634 11756 13690 11792
rect 13634 11736 13636 11756
rect 13636 11736 13688 11756
rect 13688 11736 13690 11756
rect 13560 10906 13616 10908
rect 13640 10906 13696 10908
rect 13720 10906 13776 10908
rect 13800 10906 13856 10908
rect 13560 10854 13606 10906
rect 13606 10854 13616 10906
rect 13640 10854 13670 10906
rect 13670 10854 13682 10906
rect 13682 10854 13696 10906
rect 13720 10854 13734 10906
rect 13734 10854 13746 10906
rect 13746 10854 13776 10906
rect 13800 10854 13810 10906
rect 13810 10854 13856 10906
rect 13560 10852 13616 10854
rect 13640 10852 13696 10854
rect 13720 10852 13776 10854
rect 13800 10852 13856 10854
rect 13560 9818 13616 9820
rect 13640 9818 13696 9820
rect 13720 9818 13776 9820
rect 13800 9818 13856 9820
rect 13560 9766 13606 9818
rect 13606 9766 13616 9818
rect 13640 9766 13670 9818
rect 13670 9766 13682 9818
rect 13682 9766 13696 9818
rect 13720 9766 13734 9818
rect 13734 9766 13746 9818
rect 13746 9766 13776 9818
rect 13800 9766 13810 9818
rect 13810 9766 13856 9818
rect 13560 9764 13616 9766
rect 13640 9764 13696 9766
rect 13720 9764 13776 9766
rect 13800 9764 13856 9766
rect 14186 12824 14242 12880
rect 13560 8730 13616 8732
rect 13640 8730 13696 8732
rect 13720 8730 13776 8732
rect 13800 8730 13856 8732
rect 13560 8678 13606 8730
rect 13606 8678 13616 8730
rect 13640 8678 13670 8730
rect 13670 8678 13682 8730
rect 13682 8678 13696 8730
rect 13720 8678 13734 8730
rect 13734 8678 13746 8730
rect 13746 8678 13776 8730
rect 13800 8678 13810 8730
rect 13810 8678 13856 8730
rect 13560 8676 13616 8678
rect 13640 8676 13696 8678
rect 13720 8676 13776 8678
rect 13800 8676 13856 8678
rect 13560 7642 13616 7644
rect 13640 7642 13696 7644
rect 13720 7642 13776 7644
rect 13800 7642 13856 7644
rect 13560 7590 13606 7642
rect 13606 7590 13616 7642
rect 13640 7590 13670 7642
rect 13670 7590 13682 7642
rect 13682 7590 13696 7642
rect 13720 7590 13734 7642
rect 13734 7590 13746 7642
rect 13746 7590 13776 7642
rect 13800 7590 13810 7642
rect 13810 7590 13856 7642
rect 13560 7588 13616 7590
rect 13640 7588 13696 7590
rect 13720 7588 13776 7590
rect 13800 7588 13856 7590
rect 13560 6554 13616 6556
rect 13640 6554 13696 6556
rect 13720 6554 13776 6556
rect 13800 6554 13856 6556
rect 13560 6502 13606 6554
rect 13606 6502 13616 6554
rect 13640 6502 13670 6554
rect 13670 6502 13682 6554
rect 13682 6502 13696 6554
rect 13720 6502 13734 6554
rect 13734 6502 13746 6554
rect 13746 6502 13776 6554
rect 13800 6502 13810 6554
rect 13810 6502 13856 6554
rect 13560 6500 13616 6502
rect 13640 6500 13696 6502
rect 13720 6500 13776 6502
rect 13800 6500 13856 6502
rect 13560 5466 13616 5468
rect 13640 5466 13696 5468
rect 13720 5466 13776 5468
rect 13800 5466 13856 5468
rect 13560 5414 13606 5466
rect 13606 5414 13616 5466
rect 13640 5414 13670 5466
rect 13670 5414 13682 5466
rect 13682 5414 13696 5466
rect 13720 5414 13734 5466
rect 13734 5414 13746 5466
rect 13746 5414 13776 5466
rect 13800 5414 13810 5466
rect 13810 5414 13856 5466
rect 13560 5412 13616 5414
rect 13640 5412 13696 5414
rect 13720 5412 13776 5414
rect 13800 5412 13856 5414
rect 13560 4378 13616 4380
rect 13640 4378 13696 4380
rect 13720 4378 13776 4380
rect 13800 4378 13856 4380
rect 13560 4326 13606 4378
rect 13606 4326 13616 4378
rect 13640 4326 13670 4378
rect 13670 4326 13682 4378
rect 13682 4326 13696 4378
rect 13720 4326 13734 4378
rect 13734 4326 13746 4378
rect 13746 4326 13776 4378
rect 13800 4326 13810 4378
rect 13810 4326 13856 4378
rect 13560 4324 13616 4326
rect 13640 4324 13696 4326
rect 13720 4324 13776 4326
rect 13800 4324 13856 4326
rect 13560 3290 13616 3292
rect 13640 3290 13696 3292
rect 13720 3290 13776 3292
rect 13800 3290 13856 3292
rect 13560 3238 13606 3290
rect 13606 3238 13616 3290
rect 13640 3238 13670 3290
rect 13670 3238 13682 3290
rect 13682 3238 13696 3290
rect 13720 3238 13734 3290
rect 13734 3238 13746 3290
rect 13746 3238 13776 3290
rect 13800 3238 13810 3290
rect 13810 3238 13856 3290
rect 13560 3236 13616 3238
rect 13640 3236 13696 3238
rect 13720 3236 13776 3238
rect 13800 3236 13856 3238
rect 10409 2746 10465 2748
rect 10489 2746 10545 2748
rect 10569 2746 10625 2748
rect 10649 2746 10705 2748
rect 10409 2694 10455 2746
rect 10455 2694 10465 2746
rect 10489 2694 10519 2746
rect 10519 2694 10531 2746
rect 10531 2694 10545 2746
rect 10569 2694 10583 2746
rect 10583 2694 10595 2746
rect 10595 2694 10625 2746
rect 10649 2694 10659 2746
rect 10659 2694 10705 2746
rect 10409 2692 10465 2694
rect 10489 2692 10545 2694
rect 10569 2692 10625 2694
rect 10649 2692 10705 2694
rect 14462 12300 14518 12336
rect 14462 12280 14464 12300
rect 14464 12280 14516 12300
rect 14516 12280 14518 12300
rect 15014 12824 15070 12880
rect 16711 26682 16767 26684
rect 16791 26682 16847 26684
rect 16871 26682 16927 26684
rect 16951 26682 17007 26684
rect 16711 26630 16757 26682
rect 16757 26630 16767 26682
rect 16791 26630 16821 26682
rect 16821 26630 16833 26682
rect 16833 26630 16847 26682
rect 16871 26630 16885 26682
rect 16885 26630 16897 26682
rect 16897 26630 16927 26682
rect 16951 26630 16961 26682
rect 16961 26630 17007 26682
rect 16711 26628 16767 26630
rect 16791 26628 16847 26630
rect 16871 26628 16927 26630
rect 16951 26628 17007 26630
rect 15842 24268 15898 24304
rect 15842 24248 15844 24268
rect 15844 24248 15896 24268
rect 15896 24248 15898 24268
rect 16711 25594 16767 25596
rect 16791 25594 16847 25596
rect 16871 25594 16927 25596
rect 16951 25594 17007 25596
rect 16711 25542 16757 25594
rect 16757 25542 16767 25594
rect 16791 25542 16821 25594
rect 16821 25542 16833 25594
rect 16833 25542 16847 25594
rect 16871 25542 16885 25594
rect 16885 25542 16897 25594
rect 16897 25542 16927 25594
rect 16951 25542 16961 25594
rect 16961 25542 17007 25594
rect 16711 25540 16767 25542
rect 16791 25540 16847 25542
rect 16871 25540 16927 25542
rect 16951 25540 17007 25542
rect 16711 24506 16767 24508
rect 16791 24506 16847 24508
rect 16871 24506 16927 24508
rect 16951 24506 17007 24508
rect 16711 24454 16757 24506
rect 16757 24454 16767 24506
rect 16791 24454 16821 24506
rect 16821 24454 16833 24506
rect 16833 24454 16847 24506
rect 16871 24454 16885 24506
rect 16885 24454 16897 24506
rect 16897 24454 16927 24506
rect 16951 24454 16961 24506
rect 16961 24454 17007 24506
rect 16711 24452 16767 24454
rect 16791 24452 16847 24454
rect 16871 24452 16927 24454
rect 16951 24452 17007 24454
rect 16711 23418 16767 23420
rect 16791 23418 16847 23420
rect 16871 23418 16927 23420
rect 16951 23418 17007 23420
rect 16711 23366 16757 23418
rect 16757 23366 16767 23418
rect 16791 23366 16821 23418
rect 16821 23366 16833 23418
rect 16833 23366 16847 23418
rect 16871 23366 16885 23418
rect 16885 23366 16897 23418
rect 16897 23366 16927 23418
rect 16951 23366 16961 23418
rect 16961 23366 17007 23418
rect 16711 23364 16767 23366
rect 16791 23364 16847 23366
rect 16871 23364 16927 23366
rect 16951 23364 17007 23366
rect 16711 22330 16767 22332
rect 16791 22330 16847 22332
rect 16871 22330 16927 22332
rect 16951 22330 17007 22332
rect 16711 22278 16757 22330
rect 16757 22278 16767 22330
rect 16791 22278 16821 22330
rect 16821 22278 16833 22330
rect 16833 22278 16847 22330
rect 16871 22278 16885 22330
rect 16885 22278 16897 22330
rect 16897 22278 16927 22330
rect 16951 22278 16961 22330
rect 16961 22278 17007 22330
rect 16711 22276 16767 22278
rect 16791 22276 16847 22278
rect 16871 22276 16927 22278
rect 16951 22276 17007 22278
rect 19862 26138 19918 26140
rect 19942 26138 19998 26140
rect 20022 26138 20078 26140
rect 20102 26138 20158 26140
rect 19862 26086 19908 26138
rect 19908 26086 19918 26138
rect 19942 26086 19972 26138
rect 19972 26086 19984 26138
rect 19984 26086 19998 26138
rect 20022 26086 20036 26138
rect 20036 26086 20048 26138
rect 20048 26086 20078 26138
rect 20102 26086 20112 26138
rect 20112 26086 20158 26138
rect 19862 26084 19918 26086
rect 19942 26084 19998 26086
rect 20022 26084 20078 26086
rect 20102 26084 20158 26086
rect 16711 21242 16767 21244
rect 16791 21242 16847 21244
rect 16871 21242 16927 21244
rect 16951 21242 17007 21244
rect 16711 21190 16757 21242
rect 16757 21190 16767 21242
rect 16791 21190 16821 21242
rect 16821 21190 16833 21242
rect 16833 21190 16847 21242
rect 16871 21190 16885 21242
rect 16885 21190 16897 21242
rect 16897 21190 16927 21242
rect 16951 21190 16961 21242
rect 16961 21190 17007 21242
rect 16711 21188 16767 21190
rect 16791 21188 16847 21190
rect 16871 21188 16927 21190
rect 16951 21188 17007 21190
rect 16210 18828 16266 18864
rect 16210 18808 16212 18828
rect 16212 18808 16264 18828
rect 16264 18808 16266 18828
rect 16118 18672 16174 18728
rect 16711 20154 16767 20156
rect 16791 20154 16847 20156
rect 16871 20154 16927 20156
rect 16951 20154 17007 20156
rect 16711 20102 16757 20154
rect 16757 20102 16767 20154
rect 16791 20102 16821 20154
rect 16821 20102 16833 20154
rect 16833 20102 16847 20154
rect 16871 20102 16885 20154
rect 16885 20102 16897 20154
rect 16897 20102 16927 20154
rect 16951 20102 16961 20154
rect 16961 20102 17007 20154
rect 16711 20100 16767 20102
rect 16791 20100 16847 20102
rect 16871 20100 16927 20102
rect 16951 20100 17007 20102
rect 16711 19066 16767 19068
rect 16791 19066 16847 19068
rect 16871 19066 16927 19068
rect 16951 19066 17007 19068
rect 16711 19014 16757 19066
rect 16757 19014 16767 19066
rect 16791 19014 16821 19066
rect 16821 19014 16833 19066
rect 16833 19014 16847 19066
rect 16871 19014 16885 19066
rect 16885 19014 16897 19066
rect 16897 19014 16927 19066
rect 16951 19014 16961 19066
rect 16961 19014 17007 19066
rect 16711 19012 16767 19014
rect 16791 19012 16847 19014
rect 16871 19012 16927 19014
rect 16951 19012 17007 19014
rect 16711 17978 16767 17980
rect 16791 17978 16847 17980
rect 16871 17978 16927 17980
rect 16951 17978 17007 17980
rect 16711 17926 16757 17978
rect 16757 17926 16767 17978
rect 16791 17926 16821 17978
rect 16821 17926 16833 17978
rect 16833 17926 16847 17978
rect 16871 17926 16885 17978
rect 16885 17926 16897 17978
rect 16897 17926 16927 17978
rect 16951 17926 16961 17978
rect 16961 17926 17007 17978
rect 16711 17924 16767 17926
rect 16791 17924 16847 17926
rect 16871 17924 16927 17926
rect 16951 17924 17007 17926
rect 17498 17720 17554 17776
rect 16711 16890 16767 16892
rect 16791 16890 16847 16892
rect 16871 16890 16927 16892
rect 16951 16890 17007 16892
rect 16711 16838 16757 16890
rect 16757 16838 16767 16890
rect 16791 16838 16821 16890
rect 16821 16838 16833 16890
rect 16833 16838 16847 16890
rect 16871 16838 16885 16890
rect 16885 16838 16897 16890
rect 16897 16838 16927 16890
rect 16951 16838 16961 16890
rect 16961 16838 17007 16890
rect 16711 16836 16767 16838
rect 16791 16836 16847 16838
rect 16871 16836 16927 16838
rect 16951 16836 17007 16838
rect 16711 15802 16767 15804
rect 16791 15802 16847 15804
rect 16871 15802 16927 15804
rect 16951 15802 17007 15804
rect 16711 15750 16757 15802
rect 16757 15750 16767 15802
rect 16791 15750 16821 15802
rect 16821 15750 16833 15802
rect 16833 15750 16847 15802
rect 16871 15750 16885 15802
rect 16885 15750 16897 15802
rect 16897 15750 16927 15802
rect 16951 15750 16961 15802
rect 16961 15750 17007 15802
rect 16711 15748 16767 15750
rect 16791 15748 16847 15750
rect 16871 15748 16927 15750
rect 16951 15748 17007 15750
rect 16762 15036 16764 15056
rect 16764 15036 16816 15056
rect 16816 15036 16818 15056
rect 16762 15000 16818 15036
rect 16711 14714 16767 14716
rect 16791 14714 16847 14716
rect 16871 14714 16927 14716
rect 16951 14714 17007 14716
rect 16711 14662 16757 14714
rect 16757 14662 16767 14714
rect 16791 14662 16821 14714
rect 16821 14662 16833 14714
rect 16833 14662 16847 14714
rect 16871 14662 16885 14714
rect 16885 14662 16897 14714
rect 16897 14662 16927 14714
rect 16951 14662 16961 14714
rect 16961 14662 17007 14714
rect 16711 14660 16767 14662
rect 16791 14660 16847 14662
rect 16871 14660 16927 14662
rect 16951 14660 17007 14662
rect 18602 24268 18658 24304
rect 18602 24248 18604 24268
rect 18604 24248 18656 24268
rect 18656 24248 18658 24268
rect 19862 25050 19918 25052
rect 19942 25050 19998 25052
rect 20022 25050 20078 25052
rect 20102 25050 20158 25052
rect 19862 24998 19908 25050
rect 19908 24998 19918 25050
rect 19942 24998 19972 25050
rect 19972 24998 19984 25050
rect 19984 24998 19998 25050
rect 20022 24998 20036 25050
rect 20036 24998 20048 25050
rect 20048 24998 20078 25050
rect 20102 24998 20112 25050
rect 20112 24998 20158 25050
rect 19862 24996 19918 24998
rect 19942 24996 19998 24998
rect 20022 24996 20078 24998
rect 20102 24996 20158 24998
rect 17682 18672 17738 18728
rect 19862 23962 19918 23964
rect 19942 23962 19998 23964
rect 20022 23962 20078 23964
rect 20102 23962 20158 23964
rect 19862 23910 19908 23962
rect 19908 23910 19918 23962
rect 19942 23910 19972 23962
rect 19972 23910 19984 23962
rect 19984 23910 19998 23962
rect 20022 23910 20036 23962
rect 20036 23910 20048 23962
rect 20048 23910 20078 23962
rect 20102 23910 20112 23962
rect 20112 23910 20158 23962
rect 19862 23908 19918 23910
rect 19942 23908 19998 23910
rect 20022 23908 20078 23910
rect 20102 23908 20158 23910
rect 16711 13626 16767 13628
rect 16791 13626 16847 13628
rect 16871 13626 16927 13628
rect 16951 13626 17007 13628
rect 16711 13574 16757 13626
rect 16757 13574 16767 13626
rect 16791 13574 16821 13626
rect 16821 13574 16833 13626
rect 16833 13574 16847 13626
rect 16871 13574 16885 13626
rect 16885 13574 16897 13626
rect 16897 13574 16927 13626
rect 16951 13574 16961 13626
rect 16961 13574 17007 13626
rect 16711 13572 16767 13574
rect 16791 13572 16847 13574
rect 16871 13572 16927 13574
rect 16951 13572 17007 13574
rect 14738 11736 14794 11792
rect 15658 12300 15714 12336
rect 15658 12280 15660 12300
rect 15660 12280 15712 12300
rect 15712 12280 15714 12300
rect 15934 12708 15990 12744
rect 15934 12688 15936 12708
rect 15936 12688 15988 12708
rect 15988 12688 15990 12708
rect 15566 11736 15622 11792
rect 16711 12538 16767 12540
rect 16791 12538 16847 12540
rect 16871 12538 16927 12540
rect 16951 12538 17007 12540
rect 16711 12486 16757 12538
rect 16757 12486 16767 12538
rect 16791 12486 16821 12538
rect 16821 12486 16833 12538
rect 16833 12486 16847 12538
rect 16871 12486 16885 12538
rect 16885 12486 16897 12538
rect 16897 12486 16927 12538
rect 16951 12486 16961 12538
rect 16961 12486 17007 12538
rect 16711 12484 16767 12486
rect 16791 12484 16847 12486
rect 16871 12484 16927 12486
rect 16951 12484 17007 12486
rect 16711 11450 16767 11452
rect 16791 11450 16847 11452
rect 16871 11450 16927 11452
rect 16951 11450 17007 11452
rect 16711 11398 16757 11450
rect 16757 11398 16767 11450
rect 16791 11398 16821 11450
rect 16821 11398 16833 11450
rect 16833 11398 16847 11450
rect 16871 11398 16885 11450
rect 16885 11398 16897 11450
rect 16897 11398 16927 11450
rect 16951 11398 16961 11450
rect 16961 11398 17007 11450
rect 16711 11396 16767 11398
rect 16791 11396 16847 11398
rect 16871 11396 16927 11398
rect 16951 11396 17007 11398
rect 16711 10362 16767 10364
rect 16791 10362 16847 10364
rect 16871 10362 16927 10364
rect 16951 10362 17007 10364
rect 16711 10310 16757 10362
rect 16757 10310 16767 10362
rect 16791 10310 16821 10362
rect 16821 10310 16833 10362
rect 16833 10310 16847 10362
rect 16871 10310 16885 10362
rect 16885 10310 16897 10362
rect 16897 10310 16927 10362
rect 16951 10310 16961 10362
rect 16961 10310 17007 10362
rect 16711 10308 16767 10310
rect 16791 10308 16847 10310
rect 16871 10308 16927 10310
rect 16951 10308 17007 10310
rect 16711 9274 16767 9276
rect 16791 9274 16847 9276
rect 16871 9274 16927 9276
rect 16951 9274 17007 9276
rect 16711 9222 16757 9274
rect 16757 9222 16767 9274
rect 16791 9222 16821 9274
rect 16821 9222 16833 9274
rect 16833 9222 16847 9274
rect 16871 9222 16885 9274
rect 16885 9222 16897 9274
rect 16897 9222 16927 9274
rect 16951 9222 16961 9274
rect 16961 9222 17007 9274
rect 16711 9220 16767 9222
rect 16791 9220 16847 9222
rect 16871 9220 16927 9222
rect 16951 9220 17007 9222
rect 16711 8186 16767 8188
rect 16791 8186 16847 8188
rect 16871 8186 16927 8188
rect 16951 8186 17007 8188
rect 16711 8134 16757 8186
rect 16757 8134 16767 8186
rect 16791 8134 16821 8186
rect 16821 8134 16833 8186
rect 16833 8134 16847 8186
rect 16871 8134 16885 8186
rect 16885 8134 16897 8186
rect 16897 8134 16927 8186
rect 16951 8134 16961 8186
rect 16961 8134 17007 8186
rect 16711 8132 16767 8134
rect 16791 8132 16847 8134
rect 16871 8132 16927 8134
rect 16951 8132 17007 8134
rect 18694 17720 18750 17776
rect 19862 22874 19918 22876
rect 19942 22874 19998 22876
rect 20022 22874 20078 22876
rect 20102 22874 20158 22876
rect 19862 22822 19908 22874
rect 19908 22822 19918 22874
rect 19942 22822 19972 22874
rect 19972 22822 19984 22874
rect 19984 22822 19998 22874
rect 20022 22822 20036 22874
rect 20036 22822 20048 22874
rect 20048 22822 20078 22874
rect 20102 22822 20112 22874
rect 20112 22822 20158 22874
rect 19862 22820 19918 22822
rect 19942 22820 19998 22822
rect 20022 22820 20078 22822
rect 20102 22820 20158 22822
rect 19862 21786 19918 21788
rect 19942 21786 19998 21788
rect 20022 21786 20078 21788
rect 20102 21786 20158 21788
rect 19862 21734 19908 21786
rect 19908 21734 19918 21786
rect 19942 21734 19972 21786
rect 19972 21734 19984 21786
rect 19984 21734 19998 21786
rect 20022 21734 20036 21786
rect 20036 21734 20048 21786
rect 20048 21734 20078 21786
rect 20102 21734 20112 21786
rect 20112 21734 20158 21786
rect 19862 21732 19918 21734
rect 19942 21732 19998 21734
rect 20022 21732 20078 21734
rect 20102 21732 20158 21734
rect 19862 20698 19918 20700
rect 19942 20698 19998 20700
rect 20022 20698 20078 20700
rect 20102 20698 20158 20700
rect 19862 20646 19908 20698
rect 19908 20646 19918 20698
rect 19942 20646 19972 20698
rect 19972 20646 19984 20698
rect 19984 20646 19998 20698
rect 20022 20646 20036 20698
rect 20036 20646 20048 20698
rect 20048 20646 20078 20698
rect 20102 20646 20112 20698
rect 20112 20646 20158 20698
rect 19862 20644 19918 20646
rect 19942 20644 19998 20646
rect 20022 20644 20078 20646
rect 20102 20644 20158 20646
rect 23013 26682 23069 26684
rect 23093 26682 23149 26684
rect 23173 26682 23229 26684
rect 23253 26682 23309 26684
rect 23013 26630 23059 26682
rect 23059 26630 23069 26682
rect 23093 26630 23123 26682
rect 23123 26630 23135 26682
rect 23135 26630 23149 26682
rect 23173 26630 23187 26682
rect 23187 26630 23199 26682
rect 23199 26630 23229 26682
rect 23253 26630 23263 26682
rect 23263 26630 23309 26682
rect 23013 26628 23069 26630
rect 23093 26628 23149 26630
rect 23173 26628 23229 26630
rect 23253 26628 23309 26630
rect 21270 23704 21326 23760
rect 21914 24656 21970 24712
rect 19862 19610 19918 19612
rect 19942 19610 19998 19612
rect 20022 19610 20078 19612
rect 20102 19610 20158 19612
rect 19862 19558 19908 19610
rect 19908 19558 19918 19610
rect 19942 19558 19972 19610
rect 19972 19558 19984 19610
rect 19984 19558 19998 19610
rect 20022 19558 20036 19610
rect 20036 19558 20048 19610
rect 20048 19558 20078 19610
rect 20102 19558 20112 19610
rect 20112 19558 20158 19610
rect 19862 19556 19918 19558
rect 19942 19556 19998 19558
rect 20022 19556 20078 19558
rect 20102 19556 20158 19558
rect 19862 18522 19918 18524
rect 19942 18522 19998 18524
rect 20022 18522 20078 18524
rect 20102 18522 20158 18524
rect 19862 18470 19908 18522
rect 19908 18470 19918 18522
rect 19942 18470 19972 18522
rect 19972 18470 19984 18522
rect 19984 18470 19998 18522
rect 20022 18470 20036 18522
rect 20036 18470 20048 18522
rect 20048 18470 20078 18522
rect 20102 18470 20112 18522
rect 20112 18470 20158 18522
rect 19862 18468 19918 18470
rect 19942 18468 19998 18470
rect 20022 18468 20078 18470
rect 20102 18468 20158 18470
rect 19862 17434 19918 17436
rect 19942 17434 19998 17436
rect 20022 17434 20078 17436
rect 20102 17434 20158 17436
rect 19862 17382 19908 17434
rect 19908 17382 19918 17434
rect 19942 17382 19972 17434
rect 19972 17382 19984 17434
rect 19984 17382 19998 17434
rect 20022 17382 20036 17434
rect 20036 17382 20048 17434
rect 20048 17382 20078 17434
rect 20102 17382 20112 17434
rect 20112 17382 20158 17434
rect 19862 17380 19918 17382
rect 19942 17380 19998 17382
rect 20022 17380 20078 17382
rect 20102 17380 20158 17382
rect 19862 16346 19918 16348
rect 19942 16346 19998 16348
rect 20022 16346 20078 16348
rect 20102 16346 20158 16348
rect 19862 16294 19908 16346
rect 19908 16294 19918 16346
rect 19942 16294 19972 16346
rect 19972 16294 19984 16346
rect 19984 16294 19998 16346
rect 20022 16294 20036 16346
rect 20036 16294 20048 16346
rect 20048 16294 20078 16346
rect 20102 16294 20112 16346
rect 20112 16294 20158 16346
rect 19862 16292 19918 16294
rect 19942 16292 19998 16294
rect 20022 16292 20078 16294
rect 20102 16292 20158 16294
rect 21546 21956 21602 21992
rect 21546 21936 21548 21956
rect 21548 21936 21600 21956
rect 21600 21936 21602 21956
rect 19862 15258 19918 15260
rect 19942 15258 19998 15260
rect 20022 15258 20078 15260
rect 20102 15258 20158 15260
rect 19862 15206 19908 15258
rect 19908 15206 19918 15258
rect 19942 15206 19972 15258
rect 19972 15206 19984 15258
rect 19984 15206 19998 15258
rect 20022 15206 20036 15258
rect 20036 15206 20048 15258
rect 20048 15206 20078 15258
rect 20102 15206 20112 15258
rect 20112 15206 20158 15258
rect 19862 15204 19918 15206
rect 19942 15204 19998 15206
rect 20022 15204 20078 15206
rect 20102 15204 20158 15206
rect 19862 14170 19918 14172
rect 19942 14170 19998 14172
rect 20022 14170 20078 14172
rect 20102 14170 20158 14172
rect 19862 14118 19908 14170
rect 19908 14118 19918 14170
rect 19942 14118 19972 14170
rect 19972 14118 19984 14170
rect 19984 14118 19998 14170
rect 20022 14118 20036 14170
rect 20036 14118 20048 14170
rect 20048 14118 20078 14170
rect 20102 14118 20112 14170
rect 20112 14118 20158 14170
rect 19862 14116 19918 14118
rect 19942 14116 19998 14118
rect 20022 14116 20078 14118
rect 20102 14116 20158 14118
rect 19862 13082 19918 13084
rect 19942 13082 19998 13084
rect 20022 13082 20078 13084
rect 20102 13082 20158 13084
rect 19862 13030 19908 13082
rect 19908 13030 19918 13082
rect 19942 13030 19972 13082
rect 19972 13030 19984 13082
rect 19984 13030 19998 13082
rect 20022 13030 20036 13082
rect 20036 13030 20048 13082
rect 20048 13030 20078 13082
rect 20102 13030 20112 13082
rect 20112 13030 20158 13082
rect 19862 13028 19918 13030
rect 19942 13028 19998 13030
rect 20022 13028 20078 13030
rect 20102 13028 20158 13030
rect 19522 10668 19578 10704
rect 19522 10648 19524 10668
rect 19524 10648 19576 10668
rect 19576 10648 19578 10668
rect 19862 11994 19918 11996
rect 19942 11994 19998 11996
rect 20022 11994 20078 11996
rect 20102 11994 20158 11996
rect 19862 11942 19908 11994
rect 19908 11942 19918 11994
rect 19942 11942 19972 11994
rect 19972 11942 19984 11994
rect 19984 11942 19998 11994
rect 20022 11942 20036 11994
rect 20036 11942 20048 11994
rect 20048 11942 20078 11994
rect 20102 11942 20112 11994
rect 20112 11942 20158 11994
rect 19862 11940 19918 11942
rect 19942 11940 19998 11942
rect 20022 11940 20078 11942
rect 20102 11940 20158 11942
rect 19862 10906 19918 10908
rect 19942 10906 19998 10908
rect 20022 10906 20078 10908
rect 20102 10906 20158 10908
rect 19862 10854 19908 10906
rect 19908 10854 19918 10906
rect 19942 10854 19972 10906
rect 19972 10854 19984 10906
rect 19984 10854 19998 10906
rect 20022 10854 20036 10906
rect 20036 10854 20048 10906
rect 20048 10854 20078 10906
rect 20102 10854 20112 10906
rect 20112 10854 20158 10906
rect 19862 10852 19918 10854
rect 19942 10852 19998 10854
rect 20022 10852 20078 10854
rect 20102 10852 20158 10854
rect 22742 23704 22798 23760
rect 26164 26138 26220 26140
rect 26244 26138 26300 26140
rect 26324 26138 26380 26140
rect 26404 26138 26460 26140
rect 26164 26086 26210 26138
rect 26210 26086 26220 26138
rect 26244 26086 26274 26138
rect 26274 26086 26286 26138
rect 26286 26086 26300 26138
rect 26324 26086 26338 26138
rect 26338 26086 26350 26138
rect 26350 26086 26380 26138
rect 26404 26086 26414 26138
rect 26414 26086 26460 26138
rect 26164 26084 26220 26086
rect 26244 26084 26300 26086
rect 26324 26084 26380 26086
rect 26404 26084 26460 26086
rect 23013 25594 23069 25596
rect 23093 25594 23149 25596
rect 23173 25594 23229 25596
rect 23253 25594 23309 25596
rect 23013 25542 23059 25594
rect 23059 25542 23069 25594
rect 23093 25542 23123 25594
rect 23123 25542 23135 25594
rect 23135 25542 23149 25594
rect 23173 25542 23187 25594
rect 23187 25542 23199 25594
rect 23199 25542 23229 25594
rect 23253 25542 23263 25594
rect 23263 25542 23309 25594
rect 23013 25540 23069 25542
rect 23093 25540 23149 25542
rect 23173 25540 23229 25542
rect 23253 25540 23309 25542
rect 23013 24506 23069 24508
rect 23093 24506 23149 24508
rect 23173 24506 23229 24508
rect 23253 24506 23309 24508
rect 23013 24454 23059 24506
rect 23059 24454 23069 24506
rect 23093 24454 23123 24506
rect 23123 24454 23135 24506
rect 23135 24454 23149 24506
rect 23173 24454 23187 24506
rect 23187 24454 23199 24506
rect 23199 24454 23229 24506
rect 23253 24454 23263 24506
rect 23263 24454 23309 24506
rect 23013 24452 23069 24454
rect 23093 24452 23149 24454
rect 23173 24452 23229 24454
rect 23253 24452 23309 24454
rect 23013 23418 23069 23420
rect 23093 23418 23149 23420
rect 23173 23418 23229 23420
rect 23253 23418 23309 23420
rect 23013 23366 23059 23418
rect 23059 23366 23069 23418
rect 23093 23366 23123 23418
rect 23123 23366 23135 23418
rect 23135 23366 23149 23418
rect 23173 23366 23187 23418
rect 23187 23366 23199 23418
rect 23199 23366 23229 23418
rect 23253 23366 23263 23418
rect 23263 23366 23309 23418
rect 23013 23364 23069 23366
rect 23093 23364 23149 23366
rect 23173 23364 23229 23366
rect 23253 23364 23309 23366
rect 23013 22330 23069 22332
rect 23093 22330 23149 22332
rect 23173 22330 23229 22332
rect 23253 22330 23309 22332
rect 23013 22278 23059 22330
rect 23059 22278 23069 22330
rect 23093 22278 23123 22330
rect 23123 22278 23135 22330
rect 23135 22278 23149 22330
rect 23173 22278 23187 22330
rect 23187 22278 23199 22330
rect 23199 22278 23229 22330
rect 23253 22278 23263 22330
rect 23263 22278 23309 22330
rect 23013 22276 23069 22278
rect 23093 22276 23149 22278
rect 23173 22276 23229 22278
rect 23253 22276 23309 22278
rect 26330 25200 26386 25256
rect 26164 25050 26220 25052
rect 26244 25050 26300 25052
rect 26324 25050 26380 25052
rect 26404 25050 26460 25052
rect 26164 24998 26210 25050
rect 26210 24998 26220 25050
rect 26244 24998 26274 25050
rect 26274 24998 26286 25050
rect 26286 24998 26300 25050
rect 26324 24998 26338 25050
rect 26338 24998 26350 25050
rect 26350 24998 26380 25050
rect 26404 24998 26414 25050
rect 26414 24998 26460 25050
rect 26164 24996 26220 24998
rect 26244 24996 26300 24998
rect 26324 24996 26380 24998
rect 26404 24996 26460 24998
rect 26164 23962 26220 23964
rect 26244 23962 26300 23964
rect 26324 23962 26380 23964
rect 26404 23962 26460 23964
rect 26164 23910 26210 23962
rect 26210 23910 26220 23962
rect 26244 23910 26274 23962
rect 26274 23910 26286 23962
rect 26286 23910 26300 23962
rect 26324 23910 26338 23962
rect 26338 23910 26350 23962
rect 26350 23910 26380 23962
rect 26404 23910 26414 23962
rect 26414 23910 26460 23962
rect 26164 23908 26220 23910
rect 26244 23908 26300 23910
rect 26324 23908 26380 23910
rect 26404 23908 26460 23910
rect 26164 22874 26220 22876
rect 26244 22874 26300 22876
rect 26324 22874 26380 22876
rect 26404 22874 26460 22876
rect 26164 22822 26210 22874
rect 26210 22822 26220 22874
rect 26244 22822 26274 22874
rect 26274 22822 26286 22874
rect 26286 22822 26300 22874
rect 26324 22822 26338 22874
rect 26338 22822 26350 22874
rect 26350 22822 26380 22874
rect 26404 22822 26414 22874
rect 26414 22822 26460 22874
rect 26164 22820 26220 22822
rect 26244 22820 26300 22822
rect 26324 22820 26380 22822
rect 26404 22820 26460 22822
rect 23013 21242 23069 21244
rect 23093 21242 23149 21244
rect 23173 21242 23229 21244
rect 23253 21242 23309 21244
rect 23013 21190 23059 21242
rect 23059 21190 23069 21242
rect 23093 21190 23123 21242
rect 23123 21190 23135 21242
rect 23135 21190 23149 21242
rect 23173 21190 23187 21242
rect 23187 21190 23199 21242
rect 23199 21190 23229 21242
rect 23253 21190 23263 21242
rect 23263 21190 23309 21242
rect 23013 21188 23069 21190
rect 23093 21188 23149 21190
rect 23173 21188 23229 21190
rect 23253 21188 23309 21190
rect 23013 20154 23069 20156
rect 23093 20154 23149 20156
rect 23173 20154 23229 20156
rect 23253 20154 23309 20156
rect 23013 20102 23059 20154
rect 23059 20102 23069 20154
rect 23093 20102 23123 20154
rect 23123 20102 23135 20154
rect 23135 20102 23149 20154
rect 23173 20102 23187 20154
rect 23187 20102 23199 20154
rect 23199 20102 23229 20154
rect 23253 20102 23263 20154
rect 23263 20102 23309 20154
rect 23013 20100 23069 20102
rect 23093 20100 23149 20102
rect 23173 20100 23229 20102
rect 23253 20100 23309 20102
rect 19862 9818 19918 9820
rect 19942 9818 19998 9820
rect 20022 9818 20078 9820
rect 20102 9818 20158 9820
rect 19862 9766 19908 9818
rect 19908 9766 19918 9818
rect 19942 9766 19972 9818
rect 19972 9766 19984 9818
rect 19984 9766 19998 9818
rect 20022 9766 20036 9818
rect 20036 9766 20048 9818
rect 20048 9766 20078 9818
rect 20102 9766 20112 9818
rect 20112 9766 20158 9818
rect 19862 9764 19918 9766
rect 19942 9764 19998 9766
rect 20022 9764 20078 9766
rect 20102 9764 20158 9766
rect 16711 7098 16767 7100
rect 16791 7098 16847 7100
rect 16871 7098 16927 7100
rect 16951 7098 17007 7100
rect 16711 7046 16757 7098
rect 16757 7046 16767 7098
rect 16791 7046 16821 7098
rect 16821 7046 16833 7098
rect 16833 7046 16847 7098
rect 16871 7046 16885 7098
rect 16885 7046 16897 7098
rect 16897 7046 16927 7098
rect 16951 7046 16961 7098
rect 16961 7046 17007 7098
rect 16711 7044 16767 7046
rect 16791 7044 16847 7046
rect 16871 7044 16927 7046
rect 16951 7044 17007 7046
rect 16711 6010 16767 6012
rect 16791 6010 16847 6012
rect 16871 6010 16927 6012
rect 16951 6010 17007 6012
rect 16711 5958 16757 6010
rect 16757 5958 16767 6010
rect 16791 5958 16821 6010
rect 16821 5958 16833 6010
rect 16833 5958 16847 6010
rect 16871 5958 16885 6010
rect 16885 5958 16897 6010
rect 16897 5958 16927 6010
rect 16951 5958 16961 6010
rect 16961 5958 17007 6010
rect 16711 5956 16767 5958
rect 16791 5956 16847 5958
rect 16871 5956 16927 5958
rect 16951 5956 17007 5958
rect 16711 4922 16767 4924
rect 16791 4922 16847 4924
rect 16871 4922 16927 4924
rect 16951 4922 17007 4924
rect 16711 4870 16757 4922
rect 16757 4870 16767 4922
rect 16791 4870 16821 4922
rect 16821 4870 16833 4922
rect 16833 4870 16847 4922
rect 16871 4870 16885 4922
rect 16885 4870 16897 4922
rect 16897 4870 16927 4922
rect 16951 4870 16961 4922
rect 16961 4870 17007 4922
rect 16711 4868 16767 4870
rect 16791 4868 16847 4870
rect 16871 4868 16927 4870
rect 16951 4868 17007 4870
rect 16711 3834 16767 3836
rect 16791 3834 16847 3836
rect 16871 3834 16927 3836
rect 16951 3834 17007 3836
rect 16711 3782 16757 3834
rect 16757 3782 16767 3834
rect 16791 3782 16821 3834
rect 16821 3782 16833 3834
rect 16833 3782 16847 3834
rect 16871 3782 16885 3834
rect 16885 3782 16897 3834
rect 16897 3782 16927 3834
rect 16951 3782 16961 3834
rect 16961 3782 17007 3834
rect 16711 3780 16767 3782
rect 16791 3780 16847 3782
rect 16871 3780 16927 3782
rect 16951 3780 17007 3782
rect 19862 8730 19918 8732
rect 19942 8730 19998 8732
rect 20022 8730 20078 8732
rect 20102 8730 20158 8732
rect 19862 8678 19908 8730
rect 19908 8678 19918 8730
rect 19942 8678 19972 8730
rect 19972 8678 19984 8730
rect 19984 8678 19998 8730
rect 20022 8678 20036 8730
rect 20036 8678 20048 8730
rect 20048 8678 20078 8730
rect 20102 8678 20112 8730
rect 20112 8678 20158 8730
rect 19862 8676 19918 8678
rect 19942 8676 19998 8678
rect 20022 8676 20078 8678
rect 20102 8676 20158 8678
rect 19862 7642 19918 7644
rect 19942 7642 19998 7644
rect 20022 7642 20078 7644
rect 20102 7642 20158 7644
rect 19862 7590 19908 7642
rect 19908 7590 19918 7642
rect 19942 7590 19972 7642
rect 19972 7590 19984 7642
rect 19984 7590 19998 7642
rect 20022 7590 20036 7642
rect 20036 7590 20048 7642
rect 20048 7590 20078 7642
rect 20102 7590 20112 7642
rect 20112 7590 20158 7642
rect 19862 7588 19918 7590
rect 19942 7588 19998 7590
rect 20022 7588 20078 7590
rect 20102 7588 20158 7590
rect 21270 10648 21326 10704
rect 19862 6554 19918 6556
rect 19942 6554 19998 6556
rect 20022 6554 20078 6556
rect 20102 6554 20158 6556
rect 19862 6502 19908 6554
rect 19908 6502 19918 6554
rect 19942 6502 19972 6554
rect 19972 6502 19984 6554
rect 19984 6502 19998 6554
rect 20022 6502 20036 6554
rect 20036 6502 20048 6554
rect 20048 6502 20078 6554
rect 20102 6502 20112 6554
rect 20112 6502 20158 6554
rect 19862 6500 19918 6502
rect 19942 6500 19998 6502
rect 20022 6500 20078 6502
rect 20102 6500 20158 6502
rect 23013 19066 23069 19068
rect 23093 19066 23149 19068
rect 23173 19066 23229 19068
rect 23253 19066 23309 19068
rect 23013 19014 23059 19066
rect 23059 19014 23069 19066
rect 23093 19014 23123 19066
rect 23123 19014 23135 19066
rect 23135 19014 23149 19066
rect 23173 19014 23187 19066
rect 23187 19014 23199 19066
rect 23199 19014 23229 19066
rect 23253 19014 23263 19066
rect 23263 19014 23309 19066
rect 23013 19012 23069 19014
rect 23093 19012 23149 19014
rect 23173 19012 23229 19014
rect 23253 19012 23309 19014
rect 23013 17978 23069 17980
rect 23093 17978 23149 17980
rect 23173 17978 23229 17980
rect 23253 17978 23309 17980
rect 23013 17926 23059 17978
rect 23059 17926 23069 17978
rect 23093 17926 23123 17978
rect 23123 17926 23135 17978
rect 23135 17926 23149 17978
rect 23173 17926 23187 17978
rect 23187 17926 23199 17978
rect 23199 17926 23229 17978
rect 23253 17926 23263 17978
rect 23263 17926 23309 17978
rect 23013 17924 23069 17926
rect 23093 17924 23149 17926
rect 23173 17924 23229 17926
rect 23253 17924 23309 17926
rect 23013 16890 23069 16892
rect 23093 16890 23149 16892
rect 23173 16890 23229 16892
rect 23253 16890 23309 16892
rect 23013 16838 23059 16890
rect 23059 16838 23069 16890
rect 23093 16838 23123 16890
rect 23123 16838 23135 16890
rect 23135 16838 23149 16890
rect 23173 16838 23187 16890
rect 23187 16838 23199 16890
rect 23199 16838 23229 16890
rect 23253 16838 23263 16890
rect 23263 16838 23309 16890
rect 23013 16836 23069 16838
rect 23093 16836 23149 16838
rect 23173 16836 23229 16838
rect 23253 16836 23309 16838
rect 23013 15802 23069 15804
rect 23093 15802 23149 15804
rect 23173 15802 23229 15804
rect 23253 15802 23309 15804
rect 23013 15750 23059 15802
rect 23059 15750 23069 15802
rect 23093 15750 23123 15802
rect 23123 15750 23135 15802
rect 23135 15750 23149 15802
rect 23173 15750 23187 15802
rect 23187 15750 23199 15802
rect 23199 15750 23229 15802
rect 23253 15750 23263 15802
rect 23263 15750 23309 15802
rect 23013 15748 23069 15750
rect 23093 15748 23149 15750
rect 23173 15748 23229 15750
rect 23253 15748 23309 15750
rect 23013 14714 23069 14716
rect 23093 14714 23149 14716
rect 23173 14714 23229 14716
rect 23253 14714 23309 14716
rect 23013 14662 23059 14714
rect 23059 14662 23069 14714
rect 23093 14662 23123 14714
rect 23123 14662 23135 14714
rect 23135 14662 23149 14714
rect 23173 14662 23187 14714
rect 23187 14662 23199 14714
rect 23199 14662 23229 14714
rect 23253 14662 23263 14714
rect 23263 14662 23309 14714
rect 23013 14660 23069 14662
rect 23093 14660 23149 14662
rect 23173 14660 23229 14662
rect 23253 14660 23309 14662
rect 23013 13626 23069 13628
rect 23093 13626 23149 13628
rect 23173 13626 23229 13628
rect 23253 13626 23309 13628
rect 23013 13574 23059 13626
rect 23059 13574 23069 13626
rect 23093 13574 23123 13626
rect 23123 13574 23135 13626
rect 23135 13574 23149 13626
rect 23173 13574 23187 13626
rect 23187 13574 23199 13626
rect 23199 13574 23229 13626
rect 23253 13574 23263 13626
rect 23263 13574 23309 13626
rect 23013 13572 23069 13574
rect 23093 13572 23149 13574
rect 23173 13572 23229 13574
rect 23253 13572 23309 13574
rect 23013 12538 23069 12540
rect 23093 12538 23149 12540
rect 23173 12538 23229 12540
rect 23253 12538 23309 12540
rect 23013 12486 23059 12538
rect 23059 12486 23069 12538
rect 23093 12486 23123 12538
rect 23123 12486 23135 12538
rect 23135 12486 23149 12538
rect 23173 12486 23187 12538
rect 23187 12486 23199 12538
rect 23199 12486 23229 12538
rect 23253 12486 23263 12538
rect 23263 12486 23309 12538
rect 23013 12484 23069 12486
rect 23093 12484 23149 12486
rect 23173 12484 23229 12486
rect 23253 12484 23309 12486
rect 23013 11450 23069 11452
rect 23093 11450 23149 11452
rect 23173 11450 23229 11452
rect 23253 11450 23309 11452
rect 23013 11398 23059 11450
rect 23059 11398 23069 11450
rect 23093 11398 23123 11450
rect 23123 11398 23135 11450
rect 23135 11398 23149 11450
rect 23173 11398 23187 11450
rect 23187 11398 23199 11450
rect 23199 11398 23229 11450
rect 23253 11398 23263 11450
rect 23263 11398 23309 11450
rect 23013 11396 23069 11398
rect 23093 11396 23149 11398
rect 23173 11396 23229 11398
rect 23253 11396 23309 11398
rect 23013 10362 23069 10364
rect 23093 10362 23149 10364
rect 23173 10362 23229 10364
rect 23253 10362 23309 10364
rect 23013 10310 23059 10362
rect 23059 10310 23069 10362
rect 23093 10310 23123 10362
rect 23123 10310 23135 10362
rect 23135 10310 23149 10362
rect 23173 10310 23187 10362
rect 23187 10310 23199 10362
rect 23199 10310 23229 10362
rect 23253 10310 23263 10362
rect 23263 10310 23309 10362
rect 23013 10308 23069 10310
rect 23093 10308 23149 10310
rect 23173 10308 23229 10310
rect 23253 10308 23309 10310
rect 23013 9274 23069 9276
rect 23093 9274 23149 9276
rect 23173 9274 23229 9276
rect 23253 9274 23309 9276
rect 23013 9222 23059 9274
rect 23059 9222 23069 9274
rect 23093 9222 23123 9274
rect 23123 9222 23135 9274
rect 23135 9222 23149 9274
rect 23173 9222 23187 9274
rect 23187 9222 23199 9274
rect 23199 9222 23229 9274
rect 23253 9222 23263 9274
rect 23263 9222 23309 9274
rect 23013 9220 23069 9222
rect 23093 9220 23149 9222
rect 23173 9220 23229 9222
rect 23253 9220 23309 9222
rect 26164 21786 26220 21788
rect 26244 21786 26300 21788
rect 26324 21786 26380 21788
rect 26404 21786 26460 21788
rect 26164 21734 26210 21786
rect 26210 21734 26220 21786
rect 26244 21734 26274 21786
rect 26274 21734 26286 21786
rect 26286 21734 26300 21786
rect 26324 21734 26338 21786
rect 26338 21734 26350 21786
rect 26350 21734 26380 21786
rect 26404 21734 26414 21786
rect 26414 21734 26460 21786
rect 26164 21732 26220 21734
rect 26244 21732 26300 21734
rect 26324 21732 26380 21734
rect 26404 21732 26460 21734
rect 25870 21120 25926 21176
rect 26164 20698 26220 20700
rect 26244 20698 26300 20700
rect 26324 20698 26380 20700
rect 26404 20698 26460 20700
rect 26164 20646 26210 20698
rect 26210 20646 26220 20698
rect 26244 20646 26274 20698
rect 26274 20646 26286 20698
rect 26286 20646 26300 20698
rect 26324 20646 26338 20698
rect 26338 20646 26350 20698
rect 26350 20646 26380 20698
rect 26404 20646 26414 20698
rect 26414 20646 26460 20698
rect 26164 20644 26220 20646
rect 26244 20644 26300 20646
rect 26324 20644 26380 20646
rect 26404 20644 26460 20646
rect 26164 19610 26220 19612
rect 26244 19610 26300 19612
rect 26324 19610 26380 19612
rect 26404 19610 26460 19612
rect 26164 19558 26210 19610
rect 26210 19558 26220 19610
rect 26244 19558 26274 19610
rect 26274 19558 26286 19610
rect 26286 19558 26300 19610
rect 26324 19558 26338 19610
rect 26338 19558 26350 19610
rect 26350 19558 26380 19610
rect 26404 19558 26414 19610
rect 26414 19558 26460 19610
rect 26164 19556 26220 19558
rect 26244 19556 26300 19558
rect 26324 19556 26380 19558
rect 26404 19556 26460 19558
rect 26164 18522 26220 18524
rect 26244 18522 26300 18524
rect 26324 18522 26380 18524
rect 26404 18522 26460 18524
rect 26164 18470 26210 18522
rect 26210 18470 26220 18522
rect 26244 18470 26274 18522
rect 26274 18470 26286 18522
rect 26286 18470 26300 18522
rect 26324 18470 26338 18522
rect 26338 18470 26350 18522
rect 26350 18470 26380 18522
rect 26404 18470 26414 18522
rect 26414 18470 26460 18522
rect 26164 18468 26220 18470
rect 26244 18468 26300 18470
rect 26324 18468 26380 18470
rect 26404 18468 26460 18470
rect 26164 17434 26220 17436
rect 26244 17434 26300 17436
rect 26324 17434 26380 17436
rect 26404 17434 26460 17436
rect 26164 17382 26210 17434
rect 26210 17382 26220 17434
rect 26244 17382 26274 17434
rect 26274 17382 26286 17434
rect 26286 17382 26300 17434
rect 26324 17382 26338 17434
rect 26338 17382 26350 17434
rect 26350 17382 26380 17434
rect 26404 17382 26414 17434
rect 26414 17382 26460 17434
rect 26164 17380 26220 17382
rect 26244 17380 26300 17382
rect 26324 17380 26380 17382
rect 26404 17380 26460 17382
rect 26330 17076 26332 17096
rect 26332 17076 26384 17096
rect 26384 17076 26386 17096
rect 26330 17040 26386 17076
rect 26164 16346 26220 16348
rect 26244 16346 26300 16348
rect 26324 16346 26380 16348
rect 26404 16346 26460 16348
rect 26164 16294 26210 16346
rect 26210 16294 26220 16346
rect 26244 16294 26274 16346
rect 26274 16294 26286 16346
rect 26286 16294 26300 16346
rect 26324 16294 26338 16346
rect 26338 16294 26350 16346
rect 26350 16294 26380 16346
rect 26404 16294 26414 16346
rect 26414 16294 26460 16346
rect 26164 16292 26220 16294
rect 26244 16292 26300 16294
rect 26324 16292 26380 16294
rect 26404 16292 26460 16294
rect 26164 15258 26220 15260
rect 26244 15258 26300 15260
rect 26324 15258 26380 15260
rect 26404 15258 26460 15260
rect 26164 15206 26210 15258
rect 26210 15206 26220 15258
rect 26244 15206 26274 15258
rect 26274 15206 26286 15258
rect 26286 15206 26300 15258
rect 26324 15206 26338 15258
rect 26338 15206 26350 15258
rect 26350 15206 26380 15258
rect 26404 15206 26414 15258
rect 26414 15206 26460 15258
rect 26164 15204 26220 15206
rect 26244 15204 26300 15206
rect 26324 15204 26380 15206
rect 26404 15204 26460 15206
rect 26164 14170 26220 14172
rect 26244 14170 26300 14172
rect 26324 14170 26380 14172
rect 26404 14170 26460 14172
rect 26164 14118 26210 14170
rect 26210 14118 26220 14170
rect 26244 14118 26274 14170
rect 26274 14118 26286 14170
rect 26286 14118 26300 14170
rect 26324 14118 26338 14170
rect 26338 14118 26350 14170
rect 26350 14118 26380 14170
rect 26404 14118 26414 14170
rect 26414 14118 26460 14170
rect 26164 14116 26220 14118
rect 26244 14116 26300 14118
rect 26324 14116 26380 14118
rect 26404 14116 26460 14118
rect 25410 12688 25466 12744
rect 25870 13232 25926 13288
rect 26164 13082 26220 13084
rect 26244 13082 26300 13084
rect 26324 13082 26380 13084
rect 26404 13082 26460 13084
rect 26164 13030 26210 13082
rect 26210 13030 26220 13082
rect 26244 13030 26274 13082
rect 26274 13030 26286 13082
rect 26286 13030 26300 13082
rect 26324 13030 26338 13082
rect 26338 13030 26350 13082
rect 26350 13030 26380 13082
rect 26404 13030 26414 13082
rect 26414 13030 26460 13082
rect 26164 13028 26220 13030
rect 26244 13028 26300 13030
rect 26324 13028 26380 13030
rect 26404 13028 26460 13030
rect 26164 11994 26220 11996
rect 26244 11994 26300 11996
rect 26324 11994 26380 11996
rect 26404 11994 26460 11996
rect 26164 11942 26210 11994
rect 26210 11942 26220 11994
rect 26244 11942 26274 11994
rect 26274 11942 26286 11994
rect 26286 11942 26300 11994
rect 26324 11942 26338 11994
rect 26338 11942 26350 11994
rect 26350 11942 26380 11994
rect 26404 11942 26414 11994
rect 26414 11942 26460 11994
rect 26164 11940 26220 11942
rect 26244 11940 26300 11942
rect 26324 11940 26380 11942
rect 26404 11940 26460 11942
rect 26164 10906 26220 10908
rect 26244 10906 26300 10908
rect 26324 10906 26380 10908
rect 26404 10906 26460 10908
rect 26164 10854 26210 10906
rect 26210 10854 26220 10906
rect 26244 10854 26274 10906
rect 26274 10854 26286 10906
rect 26286 10854 26300 10906
rect 26324 10854 26338 10906
rect 26338 10854 26350 10906
rect 26350 10854 26380 10906
rect 26404 10854 26414 10906
rect 26414 10854 26460 10906
rect 26164 10852 26220 10854
rect 26244 10852 26300 10854
rect 26324 10852 26380 10854
rect 26404 10852 26460 10854
rect 26164 9818 26220 9820
rect 26244 9818 26300 9820
rect 26324 9818 26380 9820
rect 26404 9818 26460 9820
rect 26164 9766 26210 9818
rect 26210 9766 26220 9818
rect 26244 9766 26274 9818
rect 26274 9766 26286 9818
rect 26286 9766 26300 9818
rect 26324 9766 26338 9818
rect 26338 9766 26350 9818
rect 26350 9766 26380 9818
rect 26404 9766 26414 9818
rect 26414 9766 26460 9818
rect 26164 9764 26220 9766
rect 26244 9764 26300 9766
rect 26324 9764 26380 9766
rect 26404 9764 26460 9766
rect 23013 8186 23069 8188
rect 23093 8186 23149 8188
rect 23173 8186 23229 8188
rect 23253 8186 23309 8188
rect 23013 8134 23059 8186
rect 23059 8134 23069 8186
rect 23093 8134 23123 8186
rect 23123 8134 23135 8186
rect 23135 8134 23149 8186
rect 23173 8134 23187 8186
rect 23187 8134 23199 8186
rect 23199 8134 23229 8186
rect 23253 8134 23263 8186
rect 23263 8134 23309 8186
rect 23013 8132 23069 8134
rect 23093 8132 23149 8134
rect 23173 8132 23229 8134
rect 23253 8132 23309 8134
rect 23013 7098 23069 7100
rect 23093 7098 23149 7100
rect 23173 7098 23229 7100
rect 23253 7098 23309 7100
rect 23013 7046 23059 7098
rect 23059 7046 23069 7098
rect 23093 7046 23123 7098
rect 23123 7046 23135 7098
rect 23135 7046 23149 7098
rect 23173 7046 23187 7098
rect 23187 7046 23199 7098
rect 23199 7046 23229 7098
rect 23253 7046 23263 7098
rect 23263 7046 23309 7098
rect 23013 7044 23069 7046
rect 23093 7044 23149 7046
rect 23173 7044 23229 7046
rect 23253 7044 23309 7046
rect 19862 5466 19918 5468
rect 19942 5466 19998 5468
rect 20022 5466 20078 5468
rect 20102 5466 20158 5468
rect 19862 5414 19908 5466
rect 19908 5414 19918 5466
rect 19942 5414 19972 5466
rect 19972 5414 19984 5466
rect 19984 5414 19998 5466
rect 20022 5414 20036 5466
rect 20036 5414 20048 5466
rect 20048 5414 20078 5466
rect 20102 5414 20112 5466
rect 20112 5414 20158 5466
rect 19862 5412 19918 5414
rect 19942 5412 19998 5414
rect 20022 5412 20078 5414
rect 20102 5412 20158 5414
rect 19862 4378 19918 4380
rect 19942 4378 19998 4380
rect 20022 4378 20078 4380
rect 20102 4378 20158 4380
rect 19862 4326 19908 4378
rect 19908 4326 19918 4378
rect 19942 4326 19972 4378
rect 19972 4326 19984 4378
rect 19984 4326 19998 4378
rect 20022 4326 20036 4378
rect 20036 4326 20048 4378
rect 20048 4326 20078 4378
rect 20102 4326 20112 4378
rect 20112 4326 20158 4378
rect 19862 4324 19918 4326
rect 19942 4324 19998 4326
rect 20022 4324 20078 4326
rect 20102 4324 20158 4326
rect 26164 8730 26220 8732
rect 26244 8730 26300 8732
rect 26324 8730 26380 8732
rect 26404 8730 26460 8732
rect 26164 8678 26210 8730
rect 26210 8678 26220 8730
rect 26244 8678 26274 8730
rect 26274 8678 26286 8730
rect 26286 8678 26300 8730
rect 26324 8678 26338 8730
rect 26338 8678 26350 8730
rect 26350 8678 26380 8730
rect 26404 8678 26414 8730
rect 26414 8678 26460 8730
rect 26164 8676 26220 8678
rect 26244 8676 26300 8678
rect 26324 8676 26380 8678
rect 26404 8676 26460 8678
rect 25962 8200 26018 8256
rect 26164 7642 26220 7644
rect 26244 7642 26300 7644
rect 26324 7642 26380 7644
rect 26404 7642 26460 7644
rect 26164 7590 26210 7642
rect 26210 7590 26220 7642
rect 26244 7590 26274 7642
rect 26274 7590 26286 7642
rect 26286 7590 26300 7642
rect 26324 7590 26338 7642
rect 26338 7590 26350 7642
rect 26350 7590 26380 7642
rect 26404 7590 26414 7642
rect 26414 7590 26460 7642
rect 26164 7588 26220 7590
rect 26244 7588 26300 7590
rect 26324 7588 26380 7590
rect 26404 7588 26460 7590
rect 26164 6554 26220 6556
rect 26244 6554 26300 6556
rect 26324 6554 26380 6556
rect 26404 6554 26460 6556
rect 26164 6502 26210 6554
rect 26210 6502 26220 6554
rect 26244 6502 26274 6554
rect 26274 6502 26286 6554
rect 26286 6502 26300 6554
rect 26324 6502 26338 6554
rect 26338 6502 26350 6554
rect 26350 6502 26380 6554
rect 26404 6502 26414 6554
rect 26414 6502 26460 6554
rect 26164 6500 26220 6502
rect 26244 6500 26300 6502
rect 26324 6500 26380 6502
rect 26404 6500 26460 6502
rect 23013 6010 23069 6012
rect 23093 6010 23149 6012
rect 23173 6010 23229 6012
rect 23253 6010 23309 6012
rect 23013 5958 23059 6010
rect 23059 5958 23069 6010
rect 23093 5958 23123 6010
rect 23123 5958 23135 6010
rect 23135 5958 23149 6010
rect 23173 5958 23187 6010
rect 23187 5958 23199 6010
rect 23199 5958 23229 6010
rect 23253 5958 23263 6010
rect 23263 5958 23309 6010
rect 23013 5956 23069 5958
rect 23093 5956 23149 5958
rect 23173 5956 23229 5958
rect 23253 5956 23309 5958
rect 23013 4922 23069 4924
rect 23093 4922 23149 4924
rect 23173 4922 23229 4924
rect 23253 4922 23309 4924
rect 23013 4870 23059 4922
rect 23059 4870 23069 4922
rect 23093 4870 23123 4922
rect 23123 4870 23135 4922
rect 23135 4870 23149 4922
rect 23173 4870 23187 4922
rect 23187 4870 23199 4922
rect 23199 4870 23229 4922
rect 23253 4870 23263 4922
rect 23263 4870 23309 4922
rect 23013 4868 23069 4870
rect 23093 4868 23149 4870
rect 23173 4868 23229 4870
rect 23253 4868 23309 4870
rect 23013 3834 23069 3836
rect 23093 3834 23149 3836
rect 23173 3834 23229 3836
rect 23253 3834 23309 3836
rect 23013 3782 23059 3834
rect 23059 3782 23069 3834
rect 23093 3782 23123 3834
rect 23123 3782 23135 3834
rect 23135 3782 23149 3834
rect 23173 3782 23187 3834
rect 23187 3782 23199 3834
rect 23199 3782 23229 3834
rect 23253 3782 23263 3834
rect 23263 3782 23309 3834
rect 23013 3780 23069 3782
rect 23093 3780 23149 3782
rect 23173 3780 23229 3782
rect 23253 3780 23309 3782
rect 19862 3290 19918 3292
rect 19942 3290 19998 3292
rect 20022 3290 20078 3292
rect 20102 3290 20158 3292
rect 19862 3238 19908 3290
rect 19908 3238 19918 3290
rect 19942 3238 19972 3290
rect 19972 3238 19984 3290
rect 19984 3238 19998 3290
rect 20022 3238 20036 3290
rect 20036 3238 20048 3290
rect 20048 3238 20078 3290
rect 20102 3238 20112 3290
rect 20112 3238 20158 3290
rect 19862 3236 19918 3238
rect 19942 3236 19998 3238
rect 20022 3236 20078 3238
rect 20102 3236 20158 3238
rect 16711 2746 16767 2748
rect 16791 2746 16847 2748
rect 16871 2746 16927 2748
rect 16951 2746 17007 2748
rect 16711 2694 16757 2746
rect 16757 2694 16767 2746
rect 16791 2694 16821 2746
rect 16821 2694 16833 2746
rect 16833 2694 16847 2746
rect 16871 2694 16885 2746
rect 16885 2694 16897 2746
rect 16897 2694 16927 2746
rect 16951 2694 16961 2746
rect 16961 2694 17007 2746
rect 16711 2692 16767 2694
rect 16791 2692 16847 2694
rect 16871 2692 16927 2694
rect 16951 2692 17007 2694
rect 23013 2746 23069 2748
rect 23093 2746 23149 2748
rect 23173 2746 23229 2748
rect 23253 2746 23309 2748
rect 23013 2694 23059 2746
rect 23059 2694 23069 2746
rect 23093 2694 23123 2746
rect 23123 2694 23135 2746
rect 23135 2694 23149 2746
rect 23173 2694 23187 2746
rect 23187 2694 23199 2746
rect 23199 2694 23229 2746
rect 23253 2694 23263 2746
rect 23263 2694 23309 2746
rect 23013 2692 23069 2694
rect 23093 2692 23149 2694
rect 23173 2692 23229 2694
rect 23253 2692 23309 2694
rect 26164 5466 26220 5468
rect 26244 5466 26300 5468
rect 26324 5466 26380 5468
rect 26404 5466 26460 5468
rect 26164 5414 26210 5466
rect 26210 5414 26220 5466
rect 26244 5414 26274 5466
rect 26274 5414 26286 5466
rect 26286 5414 26300 5466
rect 26324 5414 26338 5466
rect 26338 5414 26350 5466
rect 26350 5414 26380 5466
rect 26404 5414 26414 5466
rect 26414 5414 26460 5466
rect 26164 5412 26220 5414
rect 26244 5412 26300 5414
rect 26324 5412 26380 5414
rect 26404 5412 26460 5414
rect 26164 4378 26220 4380
rect 26244 4378 26300 4380
rect 26324 4378 26380 4380
rect 26404 4378 26460 4380
rect 26164 4326 26210 4378
rect 26210 4326 26220 4378
rect 26244 4326 26274 4378
rect 26274 4326 26286 4378
rect 26286 4326 26300 4378
rect 26324 4326 26338 4378
rect 26338 4326 26350 4378
rect 26350 4326 26380 4378
rect 26404 4326 26414 4378
rect 26414 4326 26460 4378
rect 26164 4324 26220 4326
rect 26244 4324 26300 4326
rect 26324 4324 26380 4326
rect 26404 4324 26460 4326
rect 25962 4120 26018 4176
rect 26164 3290 26220 3292
rect 26244 3290 26300 3292
rect 26324 3290 26380 3292
rect 26404 3290 26460 3292
rect 26164 3238 26210 3290
rect 26210 3238 26220 3290
rect 26244 3238 26274 3290
rect 26274 3238 26286 3290
rect 26286 3238 26300 3290
rect 26324 3238 26338 3290
rect 26338 3238 26350 3290
rect 26350 3238 26380 3290
rect 26404 3238 26414 3290
rect 26414 3238 26460 3290
rect 26164 3236 26220 3238
rect 26244 3236 26300 3238
rect 26324 3236 26380 3238
rect 26404 3236 26460 3238
rect 7258 2202 7314 2204
rect 7338 2202 7394 2204
rect 7418 2202 7474 2204
rect 7498 2202 7554 2204
rect 7258 2150 7304 2202
rect 7304 2150 7314 2202
rect 7338 2150 7368 2202
rect 7368 2150 7380 2202
rect 7380 2150 7394 2202
rect 7418 2150 7432 2202
rect 7432 2150 7444 2202
rect 7444 2150 7474 2202
rect 7498 2150 7508 2202
rect 7508 2150 7554 2202
rect 7258 2148 7314 2150
rect 7338 2148 7394 2150
rect 7418 2148 7474 2150
rect 7498 2148 7554 2150
rect 13560 2202 13616 2204
rect 13640 2202 13696 2204
rect 13720 2202 13776 2204
rect 13800 2202 13856 2204
rect 13560 2150 13606 2202
rect 13606 2150 13616 2202
rect 13640 2150 13670 2202
rect 13670 2150 13682 2202
rect 13682 2150 13696 2202
rect 13720 2150 13734 2202
rect 13734 2150 13746 2202
rect 13746 2150 13776 2202
rect 13800 2150 13810 2202
rect 13810 2150 13856 2202
rect 13560 2148 13616 2150
rect 13640 2148 13696 2150
rect 13720 2148 13776 2150
rect 13800 2148 13856 2150
rect 19862 2202 19918 2204
rect 19942 2202 19998 2204
rect 20022 2202 20078 2204
rect 20102 2202 20158 2204
rect 19862 2150 19908 2202
rect 19908 2150 19918 2202
rect 19942 2150 19972 2202
rect 19972 2150 19984 2202
rect 19984 2150 19998 2202
rect 20022 2150 20036 2202
rect 20036 2150 20048 2202
rect 20048 2150 20078 2202
rect 20102 2150 20112 2202
rect 20112 2150 20158 2202
rect 19862 2148 19918 2150
rect 19942 2148 19998 2150
rect 20022 2148 20078 2150
rect 20102 2148 20158 2150
rect 26164 2202 26220 2204
rect 26244 2202 26300 2204
rect 26324 2202 26380 2204
rect 26404 2202 26460 2204
rect 26164 2150 26210 2202
rect 26210 2150 26220 2202
rect 26244 2150 26274 2202
rect 26274 2150 26286 2202
rect 26286 2150 26300 2202
rect 26324 2150 26338 2202
rect 26338 2150 26350 2202
rect 26350 2150 26380 2202
rect 26404 2150 26414 2202
rect 26414 2150 26460 2202
rect 26164 2148 26220 2150
rect 26244 2148 26300 2150
rect 26324 2148 26380 2150
rect 26404 2148 26460 2150
rect 24766 40 24822 96
<< metal3 >>
rect 0 29338 800 29368
rect 2773 29338 2839 29341
rect 0 29336 2839 29338
rect 0 29280 2778 29336
rect 2834 29280 2839 29336
rect 0 29278 2839 29280
rect 0 29248 800 29278
rect 2773 29275 2839 29278
rect 7248 27232 7564 27233
rect 7248 27168 7254 27232
rect 7318 27168 7334 27232
rect 7398 27168 7414 27232
rect 7478 27168 7494 27232
rect 7558 27168 7564 27232
rect 7248 27167 7564 27168
rect 13550 27232 13866 27233
rect 13550 27168 13556 27232
rect 13620 27168 13636 27232
rect 13700 27168 13716 27232
rect 13780 27168 13796 27232
rect 13860 27168 13866 27232
rect 13550 27167 13866 27168
rect 19852 27232 20168 27233
rect 19852 27168 19858 27232
rect 19922 27168 19938 27232
rect 20002 27168 20018 27232
rect 20082 27168 20098 27232
rect 20162 27168 20168 27232
rect 19852 27167 20168 27168
rect 26154 27232 26470 27233
rect 26154 27168 26160 27232
rect 26224 27168 26240 27232
rect 26304 27168 26320 27232
rect 26384 27168 26400 27232
rect 26464 27168 26470 27232
rect 26154 27167 26470 27168
rect 4097 26688 4413 26689
rect 4097 26624 4103 26688
rect 4167 26624 4183 26688
rect 4247 26624 4263 26688
rect 4327 26624 4343 26688
rect 4407 26624 4413 26688
rect 4097 26623 4413 26624
rect 10399 26688 10715 26689
rect 10399 26624 10405 26688
rect 10469 26624 10485 26688
rect 10549 26624 10565 26688
rect 10629 26624 10645 26688
rect 10709 26624 10715 26688
rect 10399 26623 10715 26624
rect 16701 26688 17017 26689
rect 16701 26624 16707 26688
rect 16771 26624 16787 26688
rect 16851 26624 16867 26688
rect 16931 26624 16947 26688
rect 17011 26624 17017 26688
rect 16701 26623 17017 26624
rect 23003 26688 23319 26689
rect 23003 26624 23009 26688
rect 23073 26624 23089 26688
rect 23153 26624 23169 26688
rect 23233 26624 23249 26688
rect 23313 26624 23319 26688
rect 23003 26623 23319 26624
rect 10961 26482 11027 26485
rect 12893 26482 12959 26485
rect 14825 26482 14891 26485
rect 10961 26480 14891 26482
rect 10961 26424 10966 26480
rect 11022 26424 12898 26480
rect 12954 26424 14830 26480
rect 14886 26424 14891 26480
rect 10961 26422 14891 26424
rect 10961 26419 11027 26422
rect 12893 26419 12959 26422
rect 14825 26419 14891 26422
rect 7248 26144 7564 26145
rect 7248 26080 7254 26144
rect 7318 26080 7334 26144
rect 7398 26080 7414 26144
rect 7478 26080 7494 26144
rect 7558 26080 7564 26144
rect 7248 26079 7564 26080
rect 13550 26144 13866 26145
rect 13550 26080 13556 26144
rect 13620 26080 13636 26144
rect 13700 26080 13716 26144
rect 13780 26080 13796 26144
rect 13860 26080 13866 26144
rect 13550 26079 13866 26080
rect 19852 26144 20168 26145
rect 19852 26080 19858 26144
rect 19922 26080 19938 26144
rect 20002 26080 20018 26144
rect 20082 26080 20098 26144
rect 20162 26080 20168 26144
rect 19852 26079 20168 26080
rect 26154 26144 26470 26145
rect 26154 26080 26160 26144
rect 26224 26080 26240 26144
rect 26304 26080 26320 26144
rect 26384 26080 26400 26144
rect 26464 26080 26470 26144
rect 26154 26079 26470 26080
rect 4097 25600 4413 25601
rect 4097 25536 4103 25600
rect 4167 25536 4183 25600
rect 4247 25536 4263 25600
rect 4327 25536 4343 25600
rect 4407 25536 4413 25600
rect 4097 25535 4413 25536
rect 10399 25600 10715 25601
rect 10399 25536 10405 25600
rect 10469 25536 10485 25600
rect 10549 25536 10565 25600
rect 10629 25536 10645 25600
rect 10709 25536 10715 25600
rect 10399 25535 10715 25536
rect 16701 25600 17017 25601
rect 16701 25536 16707 25600
rect 16771 25536 16787 25600
rect 16851 25536 16867 25600
rect 16931 25536 16947 25600
rect 17011 25536 17017 25600
rect 16701 25535 17017 25536
rect 23003 25600 23319 25601
rect 23003 25536 23009 25600
rect 23073 25536 23089 25600
rect 23153 25536 23169 25600
rect 23233 25536 23249 25600
rect 23313 25536 23319 25600
rect 23003 25535 23319 25536
rect 0 25258 800 25288
rect 933 25258 999 25261
rect 0 25256 999 25258
rect 0 25200 938 25256
rect 994 25200 999 25256
rect 0 25198 999 25200
rect 0 25168 800 25198
rect 933 25195 999 25198
rect 26325 25258 26391 25261
rect 26665 25258 27465 25288
rect 26325 25256 27465 25258
rect 26325 25200 26330 25256
rect 26386 25200 27465 25256
rect 26325 25198 27465 25200
rect 26325 25195 26391 25198
rect 26665 25168 27465 25198
rect 7248 25056 7564 25057
rect 7248 24992 7254 25056
rect 7318 24992 7334 25056
rect 7398 24992 7414 25056
rect 7478 24992 7494 25056
rect 7558 24992 7564 25056
rect 7248 24991 7564 24992
rect 13550 25056 13866 25057
rect 13550 24992 13556 25056
rect 13620 24992 13636 25056
rect 13700 24992 13716 25056
rect 13780 24992 13796 25056
rect 13860 24992 13866 25056
rect 13550 24991 13866 24992
rect 19852 25056 20168 25057
rect 19852 24992 19858 25056
rect 19922 24992 19938 25056
rect 20002 24992 20018 25056
rect 20082 24992 20098 25056
rect 20162 24992 20168 25056
rect 19852 24991 20168 24992
rect 26154 25056 26470 25057
rect 26154 24992 26160 25056
rect 26224 24992 26240 25056
rect 26304 24992 26320 25056
rect 26384 24992 26400 25056
rect 26464 24992 26470 25056
rect 26154 24991 26470 24992
rect 6453 24716 6519 24717
rect 6453 24714 6500 24716
rect 6408 24712 6500 24714
rect 6408 24656 6458 24712
rect 6408 24654 6500 24656
rect 6453 24652 6500 24654
rect 6564 24652 6570 24716
rect 7557 24714 7623 24717
rect 21909 24714 21975 24717
rect 7557 24712 21975 24714
rect 7557 24656 7562 24712
rect 7618 24656 21914 24712
rect 21970 24656 21975 24712
rect 7557 24654 21975 24656
rect 6453 24651 6519 24652
rect 7557 24651 7623 24654
rect 21909 24651 21975 24654
rect 4097 24512 4413 24513
rect 4097 24448 4103 24512
rect 4167 24448 4183 24512
rect 4247 24448 4263 24512
rect 4327 24448 4343 24512
rect 4407 24448 4413 24512
rect 4097 24447 4413 24448
rect 10399 24512 10715 24513
rect 10399 24448 10405 24512
rect 10469 24448 10485 24512
rect 10549 24448 10565 24512
rect 10629 24448 10645 24512
rect 10709 24448 10715 24512
rect 10399 24447 10715 24448
rect 16701 24512 17017 24513
rect 16701 24448 16707 24512
rect 16771 24448 16787 24512
rect 16851 24448 16867 24512
rect 16931 24448 16947 24512
rect 17011 24448 17017 24512
rect 16701 24447 17017 24448
rect 23003 24512 23319 24513
rect 23003 24448 23009 24512
rect 23073 24448 23089 24512
rect 23153 24448 23169 24512
rect 23233 24448 23249 24512
rect 23313 24448 23319 24512
rect 23003 24447 23319 24448
rect 15837 24306 15903 24309
rect 18597 24306 18663 24309
rect 15837 24304 18663 24306
rect 15837 24248 15842 24304
rect 15898 24248 18602 24304
rect 18658 24248 18663 24304
rect 15837 24246 18663 24248
rect 15837 24243 15903 24246
rect 18597 24243 18663 24246
rect 7248 23968 7564 23969
rect 7248 23904 7254 23968
rect 7318 23904 7334 23968
rect 7398 23904 7414 23968
rect 7478 23904 7494 23968
rect 7558 23904 7564 23968
rect 7248 23903 7564 23904
rect 13550 23968 13866 23969
rect 13550 23904 13556 23968
rect 13620 23904 13636 23968
rect 13700 23904 13716 23968
rect 13780 23904 13796 23968
rect 13860 23904 13866 23968
rect 13550 23903 13866 23904
rect 19852 23968 20168 23969
rect 19852 23904 19858 23968
rect 19922 23904 19938 23968
rect 20002 23904 20018 23968
rect 20082 23904 20098 23968
rect 20162 23904 20168 23968
rect 19852 23903 20168 23904
rect 26154 23968 26470 23969
rect 26154 23904 26160 23968
rect 26224 23904 26240 23968
rect 26304 23904 26320 23968
rect 26384 23904 26400 23968
rect 26464 23904 26470 23968
rect 26154 23903 26470 23904
rect 21265 23762 21331 23765
rect 22737 23762 22803 23765
rect 21265 23760 22803 23762
rect 21265 23704 21270 23760
rect 21326 23704 22742 23760
rect 22798 23704 22803 23760
rect 21265 23702 22803 23704
rect 21265 23699 21331 23702
rect 22737 23699 22803 23702
rect 4097 23424 4413 23425
rect 4097 23360 4103 23424
rect 4167 23360 4183 23424
rect 4247 23360 4263 23424
rect 4327 23360 4343 23424
rect 4407 23360 4413 23424
rect 4097 23359 4413 23360
rect 10399 23424 10715 23425
rect 10399 23360 10405 23424
rect 10469 23360 10485 23424
rect 10549 23360 10565 23424
rect 10629 23360 10645 23424
rect 10709 23360 10715 23424
rect 10399 23359 10715 23360
rect 16701 23424 17017 23425
rect 16701 23360 16707 23424
rect 16771 23360 16787 23424
rect 16851 23360 16867 23424
rect 16931 23360 16947 23424
rect 17011 23360 17017 23424
rect 16701 23359 17017 23360
rect 23003 23424 23319 23425
rect 23003 23360 23009 23424
rect 23073 23360 23089 23424
rect 23153 23360 23169 23424
rect 23233 23360 23249 23424
rect 23313 23360 23319 23424
rect 23003 23359 23319 23360
rect 7248 22880 7564 22881
rect 7248 22816 7254 22880
rect 7318 22816 7334 22880
rect 7398 22816 7414 22880
rect 7478 22816 7494 22880
rect 7558 22816 7564 22880
rect 7248 22815 7564 22816
rect 13550 22880 13866 22881
rect 13550 22816 13556 22880
rect 13620 22816 13636 22880
rect 13700 22816 13716 22880
rect 13780 22816 13796 22880
rect 13860 22816 13866 22880
rect 13550 22815 13866 22816
rect 19852 22880 20168 22881
rect 19852 22816 19858 22880
rect 19922 22816 19938 22880
rect 20002 22816 20018 22880
rect 20082 22816 20098 22880
rect 20162 22816 20168 22880
rect 19852 22815 20168 22816
rect 26154 22880 26470 22881
rect 26154 22816 26160 22880
rect 26224 22816 26240 22880
rect 26304 22816 26320 22880
rect 26384 22816 26400 22880
rect 26464 22816 26470 22880
rect 26154 22815 26470 22816
rect 4097 22336 4413 22337
rect 4097 22272 4103 22336
rect 4167 22272 4183 22336
rect 4247 22272 4263 22336
rect 4327 22272 4343 22336
rect 4407 22272 4413 22336
rect 4097 22271 4413 22272
rect 10399 22336 10715 22337
rect 10399 22272 10405 22336
rect 10469 22272 10485 22336
rect 10549 22272 10565 22336
rect 10629 22272 10645 22336
rect 10709 22272 10715 22336
rect 10399 22271 10715 22272
rect 16701 22336 17017 22337
rect 16701 22272 16707 22336
rect 16771 22272 16787 22336
rect 16851 22272 16867 22336
rect 16931 22272 16947 22336
rect 17011 22272 17017 22336
rect 16701 22271 17017 22272
rect 23003 22336 23319 22337
rect 23003 22272 23009 22336
rect 23073 22272 23089 22336
rect 23153 22272 23169 22336
rect 23233 22272 23249 22336
rect 23313 22272 23319 22336
rect 23003 22271 23319 22272
rect 4981 21994 5047 21997
rect 21541 21994 21607 21997
rect 4981 21992 21607 21994
rect 4981 21936 4986 21992
rect 5042 21936 21546 21992
rect 21602 21936 21607 21992
rect 4981 21934 21607 21936
rect 4981 21931 5047 21934
rect 21541 21931 21607 21934
rect 7248 21792 7564 21793
rect 7248 21728 7254 21792
rect 7318 21728 7334 21792
rect 7398 21728 7414 21792
rect 7478 21728 7494 21792
rect 7558 21728 7564 21792
rect 7248 21727 7564 21728
rect 13550 21792 13866 21793
rect 13550 21728 13556 21792
rect 13620 21728 13636 21792
rect 13700 21728 13716 21792
rect 13780 21728 13796 21792
rect 13860 21728 13866 21792
rect 13550 21727 13866 21728
rect 19852 21792 20168 21793
rect 19852 21728 19858 21792
rect 19922 21728 19938 21792
rect 20002 21728 20018 21792
rect 20082 21728 20098 21792
rect 20162 21728 20168 21792
rect 19852 21727 20168 21728
rect 26154 21792 26470 21793
rect 26154 21728 26160 21792
rect 26224 21728 26240 21792
rect 26304 21728 26320 21792
rect 26384 21728 26400 21792
rect 26464 21728 26470 21792
rect 26154 21727 26470 21728
rect 4097 21248 4413 21249
rect 0 21178 800 21208
rect 4097 21184 4103 21248
rect 4167 21184 4183 21248
rect 4247 21184 4263 21248
rect 4327 21184 4343 21248
rect 4407 21184 4413 21248
rect 4097 21183 4413 21184
rect 10399 21248 10715 21249
rect 10399 21184 10405 21248
rect 10469 21184 10485 21248
rect 10549 21184 10565 21248
rect 10629 21184 10645 21248
rect 10709 21184 10715 21248
rect 10399 21183 10715 21184
rect 16701 21248 17017 21249
rect 16701 21184 16707 21248
rect 16771 21184 16787 21248
rect 16851 21184 16867 21248
rect 16931 21184 16947 21248
rect 17011 21184 17017 21248
rect 16701 21183 17017 21184
rect 23003 21248 23319 21249
rect 23003 21184 23009 21248
rect 23073 21184 23089 21248
rect 23153 21184 23169 21248
rect 23233 21184 23249 21248
rect 23313 21184 23319 21248
rect 23003 21183 23319 21184
rect 933 21178 999 21181
rect 0 21176 999 21178
rect 0 21120 938 21176
rect 994 21120 999 21176
rect 0 21118 999 21120
rect 0 21088 800 21118
rect 933 21115 999 21118
rect 25865 21178 25931 21181
rect 26665 21178 27465 21208
rect 25865 21176 27465 21178
rect 25865 21120 25870 21176
rect 25926 21120 27465 21176
rect 25865 21118 27465 21120
rect 25865 21115 25931 21118
rect 26665 21088 27465 21118
rect 6913 20906 6979 20909
rect 7189 20906 7255 20909
rect 6913 20904 7255 20906
rect 6913 20848 6918 20904
rect 6974 20848 7194 20904
rect 7250 20848 7255 20904
rect 6913 20846 7255 20848
rect 6913 20843 6979 20846
rect 7189 20843 7255 20846
rect 7248 20704 7564 20705
rect 7248 20640 7254 20704
rect 7318 20640 7334 20704
rect 7398 20640 7414 20704
rect 7478 20640 7494 20704
rect 7558 20640 7564 20704
rect 7248 20639 7564 20640
rect 13550 20704 13866 20705
rect 13550 20640 13556 20704
rect 13620 20640 13636 20704
rect 13700 20640 13716 20704
rect 13780 20640 13796 20704
rect 13860 20640 13866 20704
rect 13550 20639 13866 20640
rect 19852 20704 20168 20705
rect 19852 20640 19858 20704
rect 19922 20640 19938 20704
rect 20002 20640 20018 20704
rect 20082 20640 20098 20704
rect 20162 20640 20168 20704
rect 19852 20639 20168 20640
rect 26154 20704 26470 20705
rect 26154 20640 26160 20704
rect 26224 20640 26240 20704
rect 26304 20640 26320 20704
rect 26384 20640 26400 20704
rect 26464 20640 26470 20704
rect 26154 20639 26470 20640
rect 4097 20160 4413 20161
rect 4097 20096 4103 20160
rect 4167 20096 4183 20160
rect 4247 20096 4263 20160
rect 4327 20096 4343 20160
rect 4407 20096 4413 20160
rect 4097 20095 4413 20096
rect 10399 20160 10715 20161
rect 10399 20096 10405 20160
rect 10469 20096 10485 20160
rect 10549 20096 10565 20160
rect 10629 20096 10645 20160
rect 10709 20096 10715 20160
rect 10399 20095 10715 20096
rect 16701 20160 17017 20161
rect 16701 20096 16707 20160
rect 16771 20096 16787 20160
rect 16851 20096 16867 20160
rect 16931 20096 16947 20160
rect 17011 20096 17017 20160
rect 16701 20095 17017 20096
rect 23003 20160 23319 20161
rect 23003 20096 23009 20160
rect 23073 20096 23089 20160
rect 23153 20096 23169 20160
rect 23233 20096 23249 20160
rect 23313 20096 23319 20160
rect 23003 20095 23319 20096
rect 5257 19818 5323 19821
rect 6177 19818 6243 19821
rect 5257 19816 6243 19818
rect 5257 19760 5262 19816
rect 5318 19760 6182 19816
rect 6238 19760 6243 19816
rect 5257 19758 6243 19760
rect 5257 19755 5323 19758
rect 6177 19755 6243 19758
rect 7248 19616 7564 19617
rect 7248 19552 7254 19616
rect 7318 19552 7334 19616
rect 7398 19552 7414 19616
rect 7478 19552 7494 19616
rect 7558 19552 7564 19616
rect 7248 19551 7564 19552
rect 13550 19616 13866 19617
rect 13550 19552 13556 19616
rect 13620 19552 13636 19616
rect 13700 19552 13716 19616
rect 13780 19552 13796 19616
rect 13860 19552 13866 19616
rect 13550 19551 13866 19552
rect 19852 19616 20168 19617
rect 19852 19552 19858 19616
rect 19922 19552 19938 19616
rect 20002 19552 20018 19616
rect 20082 19552 20098 19616
rect 20162 19552 20168 19616
rect 19852 19551 20168 19552
rect 26154 19616 26470 19617
rect 26154 19552 26160 19616
rect 26224 19552 26240 19616
rect 26304 19552 26320 19616
rect 26384 19552 26400 19616
rect 26464 19552 26470 19616
rect 26154 19551 26470 19552
rect 6913 19274 6979 19277
rect 14457 19274 14523 19277
rect 6913 19272 14523 19274
rect 6913 19216 6918 19272
rect 6974 19216 14462 19272
rect 14518 19216 14523 19272
rect 6913 19214 14523 19216
rect 6913 19211 6979 19214
rect 14457 19211 14523 19214
rect 4097 19072 4413 19073
rect 4097 19008 4103 19072
rect 4167 19008 4183 19072
rect 4247 19008 4263 19072
rect 4327 19008 4343 19072
rect 4407 19008 4413 19072
rect 4097 19007 4413 19008
rect 10399 19072 10715 19073
rect 10399 19008 10405 19072
rect 10469 19008 10485 19072
rect 10549 19008 10565 19072
rect 10629 19008 10645 19072
rect 10709 19008 10715 19072
rect 10399 19007 10715 19008
rect 16701 19072 17017 19073
rect 16701 19008 16707 19072
rect 16771 19008 16787 19072
rect 16851 19008 16867 19072
rect 16931 19008 16947 19072
rect 17011 19008 17017 19072
rect 16701 19007 17017 19008
rect 23003 19072 23319 19073
rect 23003 19008 23009 19072
rect 23073 19008 23089 19072
rect 23153 19008 23169 19072
rect 23233 19008 23249 19072
rect 23313 19008 23319 19072
rect 23003 19007 23319 19008
rect 14641 18866 14707 18869
rect 16205 18866 16271 18869
rect 14641 18864 16271 18866
rect 14641 18808 14646 18864
rect 14702 18808 16210 18864
rect 16266 18808 16271 18864
rect 14641 18806 16271 18808
rect 14641 18803 14707 18806
rect 16205 18803 16271 18806
rect 16113 18730 16179 18733
rect 17677 18730 17743 18733
rect 16113 18728 17743 18730
rect 16113 18672 16118 18728
rect 16174 18672 17682 18728
rect 17738 18672 17743 18728
rect 16113 18670 17743 18672
rect 16113 18667 16179 18670
rect 17677 18667 17743 18670
rect 7248 18528 7564 18529
rect 7248 18464 7254 18528
rect 7318 18464 7334 18528
rect 7398 18464 7414 18528
rect 7478 18464 7494 18528
rect 7558 18464 7564 18528
rect 7248 18463 7564 18464
rect 13550 18528 13866 18529
rect 13550 18464 13556 18528
rect 13620 18464 13636 18528
rect 13700 18464 13716 18528
rect 13780 18464 13796 18528
rect 13860 18464 13866 18528
rect 13550 18463 13866 18464
rect 19852 18528 20168 18529
rect 19852 18464 19858 18528
rect 19922 18464 19938 18528
rect 20002 18464 20018 18528
rect 20082 18464 20098 18528
rect 20162 18464 20168 18528
rect 19852 18463 20168 18464
rect 26154 18528 26470 18529
rect 26154 18464 26160 18528
rect 26224 18464 26240 18528
rect 26304 18464 26320 18528
rect 26384 18464 26400 18528
rect 26464 18464 26470 18528
rect 26154 18463 26470 18464
rect 4097 17984 4413 17985
rect 4097 17920 4103 17984
rect 4167 17920 4183 17984
rect 4247 17920 4263 17984
rect 4327 17920 4343 17984
rect 4407 17920 4413 17984
rect 4097 17919 4413 17920
rect 10399 17984 10715 17985
rect 10399 17920 10405 17984
rect 10469 17920 10485 17984
rect 10549 17920 10565 17984
rect 10629 17920 10645 17984
rect 10709 17920 10715 17984
rect 10399 17919 10715 17920
rect 16701 17984 17017 17985
rect 16701 17920 16707 17984
rect 16771 17920 16787 17984
rect 16851 17920 16867 17984
rect 16931 17920 16947 17984
rect 17011 17920 17017 17984
rect 16701 17919 17017 17920
rect 23003 17984 23319 17985
rect 23003 17920 23009 17984
rect 23073 17920 23089 17984
rect 23153 17920 23169 17984
rect 23233 17920 23249 17984
rect 23313 17920 23319 17984
rect 23003 17919 23319 17920
rect 12709 17778 12775 17781
rect 17493 17778 17559 17781
rect 18689 17778 18755 17781
rect 12709 17776 18755 17778
rect 12709 17720 12714 17776
rect 12770 17720 17498 17776
rect 17554 17720 18694 17776
rect 18750 17720 18755 17776
rect 12709 17718 18755 17720
rect 12709 17715 12775 17718
rect 17493 17715 17559 17718
rect 18689 17715 18755 17718
rect 7248 17440 7564 17441
rect 7248 17376 7254 17440
rect 7318 17376 7334 17440
rect 7398 17376 7414 17440
rect 7478 17376 7494 17440
rect 7558 17376 7564 17440
rect 7248 17375 7564 17376
rect 13550 17440 13866 17441
rect 13550 17376 13556 17440
rect 13620 17376 13636 17440
rect 13700 17376 13716 17440
rect 13780 17376 13796 17440
rect 13860 17376 13866 17440
rect 13550 17375 13866 17376
rect 19852 17440 20168 17441
rect 19852 17376 19858 17440
rect 19922 17376 19938 17440
rect 20002 17376 20018 17440
rect 20082 17376 20098 17440
rect 20162 17376 20168 17440
rect 19852 17375 20168 17376
rect 26154 17440 26470 17441
rect 26154 17376 26160 17440
rect 26224 17376 26240 17440
rect 26304 17376 26320 17440
rect 26384 17376 26400 17440
rect 26464 17376 26470 17440
rect 26154 17375 26470 17376
rect 26325 17098 26391 17101
rect 26665 17098 27465 17128
rect 26325 17096 27465 17098
rect 26325 17040 26330 17096
rect 26386 17040 27465 17096
rect 26325 17038 27465 17040
rect 26325 17035 26391 17038
rect 26665 17008 27465 17038
rect 4097 16896 4413 16897
rect 4097 16832 4103 16896
rect 4167 16832 4183 16896
rect 4247 16832 4263 16896
rect 4327 16832 4343 16896
rect 4407 16832 4413 16896
rect 4097 16831 4413 16832
rect 10399 16896 10715 16897
rect 10399 16832 10405 16896
rect 10469 16832 10485 16896
rect 10549 16832 10565 16896
rect 10629 16832 10645 16896
rect 10709 16832 10715 16896
rect 10399 16831 10715 16832
rect 16701 16896 17017 16897
rect 16701 16832 16707 16896
rect 16771 16832 16787 16896
rect 16851 16832 16867 16896
rect 16931 16832 16947 16896
rect 17011 16832 17017 16896
rect 16701 16831 17017 16832
rect 23003 16896 23319 16897
rect 23003 16832 23009 16896
rect 23073 16832 23089 16896
rect 23153 16832 23169 16896
rect 23233 16832 23249 16896
rect 23313 16832 23319 16896
rect 23003 16831 23319 16832
rect 1485 16554 1551 16557
rect 798 16552 1551 16554
rect 798 16496 1490 16552
rect 1546 16496 1551 16552
rect 798 16494 1551 16496
rect 798 16448 858 16494
rect 1485 16491 1551 16494
rect 0 16358 858 16448
rect 0 16328 800 16358
rect 7248 16352 7564 16353
rect 7248 16288 7254 16352
rect 7318 16288 7334 16352
rect 7398 16288 7414 16352
rect 7478 16288 7494 16352
rect 7558 16288 7564 16352
rect 7248 16287 7564 16288
rect 13550 16352 13866 16353
rect 13550 16288 13556 16352
rect 13620 16288 13636 16352
rect 13700 16288 13716 16352
rect 13780 16288 13796 16352
rect 13860 16288 13866 16352
rect 13550 16287 13866 16288
rect 19852 16352 20168 16353
rect 19852 16288 19858 16352
rect 19922 16288 19938 16352
rect 20002 16288 20018 16352
rect 20082 16288 20098 16352
rect 20162 16288 20168 16352
rect 19852 16287 20168 16288
rect 26154 16352 26470 16353
rect 26154 16288 26160 16352
rect 26224 16288 26240 16352
rect 26304 16288 26320 16352
rect 26384 16288 26400 16352
rect 26464 16288 26470 16352
rect 26154 16287 26470 16288
rect 4097 15808 4413 15809
rect 4097 15744 4103 15808
rect 4167 15744 4183 15808
rect 4247 15744 4263 15808
rect 4327 15744 4343 15808
rect 4407 15744 4413 15808
rect 4097 15743 4413 15744
rect 10399 15808 10715 15809
rect 10399 15744 10405 15808
rect 10469 15744 10485 15808
rect 10549 15744 10565 15808
rect 10629 15744 10645 15808
rect 10709 15744 10715 15808
rect 10399 15743 10715 15744
rect 16701 15808 17017 15809
rect 16701 15744 16707 15808
rect 16771 15744 16787 15808
rect 16851 15744 16867 15808
rect 16931 15744 16947 15808
rect 17011 15744 17017 15808
rect 16701 15743 17017 15744
rect 23003 15808 23319 15809
rect 23003 15744 23009 15808
rect 23073 15744 23089 15808
rect 23153 15744 23169 15808
rect 23233 15744 23249 15808
rect 23313 15744 23319 15808
rect 23003 15743 23319 15744
rect 3233 15466 3299 15469
rect 5901 15466 5967 15469
rect 3233 15464 5967 15466
rect 3233 15408 3238 15464
rect 3294 15408 5906 15464
rect 5962 15408 5967 15464
rect 3233 15406 5967 15408
rect 3233 15403 3299 15406
rect 5901 15403 5967 15406
rect 7248 15264 7564 15265
rect 7248 15200 7254 15264
rect 7318 15200 7334 15264
rect 7398 15200 7414 15264
rect 7478 15200 7494 15264
rect 7558 15200 7564 15264
rect 7248 15199 7564 15200
rect 13550 15264 13866 15265
rect 13550 15200 13556 15264
rect 13620 15200 13636 15264
rect 13700 15200 13716 15264
rect 13780 15200 13796 15264
rect 13860 15200 13866 15264
rect 13550 15199 13866 15200
rect 19852 15264 20168 15265
rect 19852 15200 19858 15264
rect 19922 15200 19938 15264
rect 20002 15200 20018 15264
rect 20082 15200 20098 15264
rect 20162 15200 20168 15264
rect 19852 15199 20168 15200
rect 26154 15264 26470 15265
rect 26154 15200 26160 15264
rect 26224 15200 26240 15264
rect 26304 15200 26320 15264
rect 26384 15200 26400 15264
rect 26464 15200 26470 15264
rect 26154 15199 26470 15200
rect 9949 15058 10015 15061
rect 16757 15058 16823 15061
rect 9949 15056 16823 15058
rect 9949 15000 9954 15056
rect 10010 15000 16762 15056
rect 16818 15000 16823 15056
rect 9949 14998 16823 15000
rect 9949 14995 10015 14998
rect 16757 14995 16823 14998
rect 3141 14922 3207 14925
rect 6494 14922 6500 14924
rect 3141 14920 6500 14922
rect 3141 14864 3146 14920
rect 3202 14864 6500 14920
rect 3141 14862 6500 14864
rect 3141 14859 3207 14862
rect 6494 14860 6500 14862
rect 6564 14860 6570 14924
rect 4097 14720 4413 14721
rect 4097 14656 4103 14720
rect 4167 14656 4183 14720
rect 4247 14656 4263 14720
rect 4327 14656 4343 14720
rect 4407 14656 4413 14720
rect 4097 14655 4413 14656
rect 10399 14720 10715 14721
rect 10399 14656 10405 14720
rect 10469 14656 10485 14720
rect 10549 14656 10565 14720
rect 10629 14656 10645 14720
rect 10709 14656 10715 14720
rect 10399 14655 10715 14656
rect 16701 14720 17017 14721
rect 16701 14656 16707 14720
rect 16771 14656 16787 14720
rect 16851 14656 16867 14720
rect 16931 14656 16947 14720
rect 17011 14656 17017 14720
rect 16701 14655 17017 14656
rect 23003 14720 23319 14721
rect 23003 14656 23009 14720
rect 23073 14656 23089 14720
rect 23153 14656 23169 14720
rect 23233 14656 23249 14720
rect 23313 14656 23319 14720
rect 23003 14655 23319 14656
rect 7248 14176 7564 14177
rect 7248 14112 7254 14176
rect 7318 14112 7334 14176
rect 7398 14112 7414 14176
rect 7478 14112 7494 14176
rect 7558 14112 7564 14176
rect 7248 14111 7564 14112
rect 13550 14176 13866 14177
rect 13550 14112 13556 14176
rect 13620 14112 13636 14176
rect 13700 14112 13716 14176
rect 13780 14112 13796 14176
rect 13860 14112 13866 14176
rect 13550 14111 13866 14112
rect 19852 14176 20168 14177
rect 19852 14112 19858 14176
rect 19922 14112 19938 14176
rect 20002 14112 20018 14176
rect 20082 14112 20098 14176
rect 20162 14112 20168 14176
rect 19852 14111 20168 14112
rect 26154 14176 26470 14177
rect 26154 14112 26160 14176
rect 26224 14112 26240 14176
rect 26304 14112 26320 14176
rect 26384 14112 26400 14176
rect 26464 14112 26470 14176
rect 26154 14111 26470 14112
rect 4097 13632 4413 13633
rect 4097 13568 4103 13632
rect 4167 13568 4183 13632
rect 4247 13568 4263 13632
rect 4327 13568 4343 13632
rect 4407 13568 4413 13632
rect 4097 13567 4413 13568
rect 10399 13632 10715 13633
rect 10399 13568 10405 13632
rect 10469 13568 10485 13632
rect 10549 13568 10565 13632
rect 10629 13568 10645 13632
rect 10709 13568 10715 13632
rect 10399 13567 10715 13568
rect 16701 13632 17017 13633
rect 16701 13568 16707 13632
rect 16771 13568 16787 13632
rect 16851 13568 16867 13632
rect 16931 13568 16947 13632
rect 17011 13568 17017 13632
rect 16701 13567 17017 13568
rect 23003 13632 23319 13633
rect 23003 13568 23009 13632
rect 23073 13568 23089 13632
rect 23153 13568 23169 13632
rect 23233 13568 23249 13632
rect 23313 13568 23319 13632
rect 23003 13567 23319 13568
rect 25865 13290 25931 13293
rect 25865 13288 26802 13290
rect 25865 13232 25870 13288
rect 25926 13232 26802 13288
rect 25865 13230 26802 13232
rect 25865 13227 25931 13230
rect 7248 13088 7564 13089
rect 7248 13024 7254 13088
rect 7318 13024 7334 13088
rect 7398 13024 7414 13088
rect 7478 13024 7494 13088
rect 7558 13024 7564 13088
rect 7248 13023 7564 13024
rect 13550 13088 13866 13089
rect 13550 13024 13556 13088
rect 13620 13024 13636 13088
rect 13700 13024 13716 13088
rect 13780 13024 13796 13088
rect 13860 13024 13866 13088
rect 13550 13023 13866 13024
rect 19852 13088 20168 13089
rect 19852 13024 19858 13088
rect 19922 13024 19938 13088
rect 20002 13024 20018 13088
rect 20082 13024 20098 13088
rect 20162 13024 20168 13088
rect 19852 13023 20168 13024
rect 26154 13088 26470 13089
rect 26154 13024 26160 13088
rect 26224 13024 26240 13088
rect 26304 13024 26320 13088
rect 26384 13024 26400 13088
rect 26464 13024 26470 13088
rect 26742 13048 26802 13230
rect 26154 13023 26470 13024
rect 26665 12928 27465 13048
rect 13905 12882 13971 12885
rect 14181 12882 14247 12885
rect 15009 12882 15075 12885
rect 13905 12880 15075 12882
rect 13905 12824 13910 12880
rect 13966 12824 14186 12880
rect 14242 12824 15014 12880
rect 15070 12824 15075 12880
rect 13905 12822 15075 12824
rect 13905 12819 13971 12822
rect 14181 12819 14247 12822
rect 15009 12819 15075 12822
rect 15929 12746 15995 12749
rect 25405 12746 25471 12749
rect 15929 12744 25471 12746
rect 15929 12688 15934 12744
rect 15990 12688 25410 12744
rect 25466 12688 25471 12744
rect 15929 12686 25471 12688
rect 15929 12683 15995 12686
rect 25405 12683 25471 12686
rect 4097 12544 4413 12545
rect 4097 12480 4103 12544
rect 4167 12480 4183 12544
rect 4247 12480 4263 12544
rect 4327 12480 4343 12544
rect 4407 12480 4413 12544
rect 4097 12479 4413 12480
rect 10399 12544 10715 12545
rect 10399 12480 10405 12544
rect 10469 12480 10485 12544
rect 10549 12480 10565 12544
rect 10629 12480 10645 12544
rect 10709 12480 10715 12544
rect 10399 12479 10715 12480
rect 16701 12544 17017 12545
rect 16701 12480 16707 12544
rect 16771 12480 16787 12544
rect 16851 12480 16867 12544
rect 16931 12480 16947 12544
rect 17011 12480 17017 12544
rect 16701 12479 17017 12480
rect 23003 12544 23319 12545
rect 23003 12480 23009 12544
rect 23073 12480 23089 12544
rect 23153 12480 23169 12544
rect 23233 12480 23249 12544
rect 23313 12480 23319 12544
rect 23003 12479 23319 12480
rect 0 12338 800 12368
rect 933 12338 999 12341
rect 0 12336 999 12338
rect 0 12280 938 12336
rect 994 12280 999 12336
rect 0 12278 999 12280
rect 0 12248 800 12278
rect 933 12275 999 12278
rect 14457 12338 14523 12341
rect 15653 12338 15719 12341
rect 14457 12336 15719 12338
rect 14457 12280 14462 12336
rect 14518 12280 15658 12336
rect 15714 12280 15719 12336
rect 14457 12278 15719 12280
rect 14457 12275 14523 12278
rect 15653 12275 15719 12278
rect 7248 12000 7564 12001
rect 7248 11936 7254 12000
rect 7318 11936 7334 12000
rect 7398 11936 7414 12000
rect 7478 11936 7494 12000
rect 7558 11936 7564 12000
rect 7248 11935 7564 11936
rect 13550 12000 13866 12001
rect 13550 11936 13556 12000
rect 13620 11936 13636 12000
rect 13700 11936 13716 12000
rect 13780 11936 13796 12000
rect 13860 11936 13866 12000
rect 13550 11935 13866 11936
rect 19852 12000 20168 12001
rect 19852 11936 19858 12000
rect 19922 11936 19938 12000
rect 20002 11936 20018 12000
rect 20082 11936 20098 12000
rect 20162 11936 20168 12000
rect 19852 11935 20168 11936
rect 26154 12000 26470 12001
rect 26154 11936 26160 12000
rect 26224 11936 26240 12000
rect 26304 11936 26320 12000
rect 26384 11936 26400 12000
rect 26464 11936 26470 12000
rect 26154 11935 26470 11936
rect 13629 11794 13695 11797
rect 14733 11794 14799 11797
rect 15561 11794 15627 11797
rect 13629 11792 15627 11794
rect 13629 11736 13634 11792
rect 13690 11736 14738 11792
rect 14794 11736 15566 11792
rect 15622 11736 15627 11792
rect 13629 11734 15627 11736
rect 13629 11731 13695 11734
rect 14733 11731 14799 11734
rect 15561 11731 15627 11734
rect 4097 11456 4413 11457
rect 4097 11392 4103 11456
rect 4167 11392 4183 11456
rect 4247 11392 4263 11456
rect 4327 11392 4343 11456
rect 4407 11392 4413 11456
rect 4097 11391 4413 11392
rect 10399 11456 10715 11457
rect 10399 11392 10405 11456
rect 10469 11392 10485 11456
rect 10549 11392 10565 11456
rect 10629 11392 10645 11456
rect 10709 11392 10715 11456
rect 10399 11391 10715 11392
rect 16701 11456 17017 11457
rect 16701 11392 16707 11456
rect 16771 11392 16787 11456
rect 16851 11392 16867 11456
rect 16931 11392 16947 11456
rect 17011 11392 17017 11456
rect 16701 11391 17017 11392
rect 23003 11456 23319 11457
rect 23003 11392 23009 11456
rect 23073 11392 23089 11456
rect 23153 11392 23169 11456
rect 23233 11392 23249 11456
rect 23313 11392 23319 11456
rect 23003 11391 23319 11392
rect 7248 10912 7564 10913
rect 7248 10848 7254 10912
rect 7318 10848 7334 10912
rect 7398 10848 7414 10912
rect 7478 10848 7494 10912
rect 7558 10848 7564 10912
rect 7248 10847 7564 10848
rect 13550 10912 13866 10913
rect 13550 10848 13556 10912
rect 13620 10848 13636 10912
rect 13700 10848 13716 10912
rect 13780 10848 13796 10912
rect 13860 10848 13866 10912
rect 13550 10847 13866 10848
rect 19852 10912 20168 10913
rect 19852 10848 19858 10912
rect 19922 10848 19938 10912
rect 20002 10848 20018 10912
rect 20082 10848 20098 10912
rect 20162 10848 20168 10912
rect 19852 10847 20168 10848
rect 26154 10912 26470 10913
rect 26154 10848 26160 10912
rect 26224 10848 26240 10912
rect 26304 10848 26320 10912
rect 26384 10848 26400 10912
rect 26464 10848 26470 10912
rect 26154 10847 26470 10848
rect 5625 10706 5691 10709
rect 6729 10706 6795 10709
rect 5625 10704 6795 10706
rect 5625 10648 5630 10704
rect 5686 10648 6734 10704
rect 6790 10648 6795 10704
rect 5625 10646 6795 10648
rect 5625 10643 5691 10646
rect 6729 10643 6795 10646
rect 19517 10706 19583 10709
rect 21265 10706 21331 10709
rect 19517 10704 21331 10706
rect 19517 10648 19522 10704
rect 19578 10648 21270 10704
rect 21326 10648 21331 10704
rect 19517 10646 21331 10648
rect 19517 10643 19583 10646
rect 21265 10643 21331 10646
rect 9857 10570 9923 10573
rect 10685 10570 10751 10573
rect 9857 10568 10751 10570
rect 9857 10512 9862 10568
rect 9918 10512 10690 10568
rect 10746 10512 10751 10568
rect 9857 10510 10751 10512
rect 9857 10507 9923 10510
rect 10685 10507 10751 10510
rect 4097 10368 4413 10369
rect 4097 10304 4103 10368
rect 4167 10304 4183 10368
rect 4247 10304 4263 10368
rect 4327 10304 4343 10368
rect 4407 10304 4413 10368
rect 4097 10303 4413 10304
rect 10399 10368 10715 10369
rect 10399 10304 10405 10368
rect 10469 10304 10485 10368
rect 10549 10304 10565 10368
rect 10629 10304 10645 10368
rect 10709 10304 10715 10368
rect 10399 10303 10715 10304
rect 16701 10368 17017 10369
rect 16701 10304 16707 10368
rect 16771 10304 16787 10368
rect 16851 10304 16867 10368
rect 16931 10304 16947 10368
rect 17011 10304 17017 10368
rect 16701 10303 17017 10304
rect 23003 10368 23319 10369
rect 23003 10304 23009 10368
rect 23073 10304 23089 10368
rect 23153 10304 23169 10368
rect 23233 10304 23249 10368
rect 23313 10304 23319 10368
rect 23003 10303 23319 10304
rect 7248 9824 7564 9825
rect 7248 9760 7254 9824
rect 7318 9760 7334 9824
rect 7398 9760 7414 9824
rect 7478 9760 7494 9824
rect 7558 9760 7564 9824
rect 7248 9759 7564 9760
rect 13550 9824 13866 9825
rect 13550 9760 13556 9824
rect 13620 9760 13636 9824
rect 13700 9760 13716 9824
rect 13780 9760 13796 9824
rect 13860 9760 13866 9824
rect 13550 9759 13866 9760
rect 19852 9824 20168 9825
rect 19852 9760 19858 9824
rect 19922 9760 19938 9824
rect 20002 9760 20018 9824
rect 20082 9760 20098 9824
rect 20162 9760 20168 9824
rect 19852 9759 20168 9760
rect 26154 9824 26470 9825
rect 26154 9760 26160 9824
rect 26224 9760 26240 9824
rect 26304 9760 26320 9824
rect 26384 9760 26400 9824
rect 26464 9760 26470 9824
rect 26154 9759 26470 9760
rect 3877 9618 3943 9621
rect 4797 9618 4863 9621
rect 3877 9616 4863 9618
rect 3877 9560 3882 9616
rect 3938 9560 4802 9616
rect 4858 9560 4863 9616
rect 3877 9558 4863 9560
rect 3877 9555 3943 9558
rect 4797 9555 4863 9558
rect 4097 9280 4413 9281
rect 4097 9216 4103 9280
rect 4167 9216 4183 9280
rect 4247 9216 4263 9280
rect 4327 9216 4343 9280
rect 4407 9216 4413 9280
rect 4097 9215 4413 9216
rect 10399 9280 10715 9281
rect 10399 9216 10405 9280
rect 10469 9216 10485 9280
rect 10549 9216 10565 9280
rect 10629 9216 10645 9280
rect 10709 9216 10715 9280
rect 10399 9215 10715 9216
rect 16701 9280 17017 9281
rect 16701 9216 16707 9280
rect 16771 9216 16787 9280
rect 16851 9216 16867 9280
rect 16931 9216 16947 9280
rect 17011 9216 17017 9280
rect 16701 9215 17017 9216
rect 23003 9280 23319 9281
rect 23003 9216 23009 9280
rect 23073 9216 23089 9280
rect 23153 9216 23169 9280
rect 23233 9216 23249 9280
rect 23313 9216 23319 9280
rect 23003 9215 23319 9216
rect 7248 8736 7564 8737
rect 7248 8672 7254 8736
rect 7318 8672 7334 8736
rect 7398 8672 7414 8736
rect 7478 8672 7494 8736
rect 7558 8672 7564 8736
rect 7248 8671 7564 8672
rect 13550 8736 13866 8737
rect 13550 8672 13556 8736
rect 13620 8672 13636 8736
rect 13700 8672 13716 8736
rect 13780 8672 13796 8736
rect 13860 8672 13866 8736
rect 13550 8671 13866 8672
rect 19852 8736 20168 8737
rect 19852 8672 19858 8736
rect 19922 8672 19938 8736
rect 20002 8672 20018 8736
rect 20082 8672 20098 8736
rect 20162 8672 20168 8736
rect 19852 8671 20168 8672
rect 26154 8736 26470 8737
rect 26154 8672 26160 8736
rect 26224 8672 26240 8736
rect 26304 8672 26320 8736
rect 26384 8672 26400 8736
rect 26464 8672 26470 8736
rect 26154 8671 26470 8672
rect 6453 8530 6519 8533
rect 8385 8530 8451 8533
rect 6453 8528 8451 8530
rect 6453 8472 6458 8528
rect 6514 8472 8390 8528
rect 8446 8472 8451 8528
rect 6453 8470 8451 8472
rect 6453 8467 6519 8470
rect 8385 8467 8451 8470
rect 0 8258 800 8288
rect 1301 8258 1367 8261
rect 0 8256 1367 8258
rect 0 8200 1306 8256
rect 1362 8200 1367 8256
rect 0 8198 1367 8200
rect 0 8168 800 8198
rect 1301 8195 1367 8198
rect 25957 8258 26023 8261
rect 26665 8258 27465 8288
rect 25957 8256 27465 8258
rect 25957 8200 25962 8256
rect 26018 8200 27465 8256
rect 25957 8198 27465 8200
rect 25957 8195 26023 8198
rect 4097 8192 4413 8193
rect 4097 8128 4103 8192
rect 4167 8128 4183 8192
rect 4247 8128 4263 8192
rect 4327 8128 4343 8192
rect 4407 8128 4413 8192
rect 4097 8127 4413 8128
rect 10399 8192 10715 8193
rect 10399 8128 10405 8192
rect 10469 8128 10485 8192
rect 10549 8128 10565 8192
rect 10629 8128 10645 8192
rect 10709 8128 10715 8192
rect 10399 8127 10715 8128
rect 16701 8192 17017 8193
rect 16701 8128 16707 8192
rect 16771 8128 16787 8192
rect 16851 8128 16867 8192
rect 16931 8128 16947 8192
rect 17011 8128 17017 8192
rect 16701 8127 17017 8128
rect 23003 8192 23319 8193
rect 23003 8128 23009 8192
rect 23073 8128 23089 8192
rect 23153 8128 23169 8192
rect 23233 8128 23249 8192
rect 23313 8128 23319 8192
rect 26665 8168 27465 8198
rect 23003 8127 23319 8128
rect 7248 7648 7564 7649
rect 7248 7584 7254 7648
rect 7318 7584 7334 7648
rect 7398 7584 7414 7648
rect 7478 7584 7494 7648
rect 7558 7584 7564 7648
rect 7248 7583 7564 7584
rect 13550 7648 13866 7649
rect 13550 7584 13556 7648
rect 13620 7584 13636 7648
rect 13700 7584 13716 7648
rect 13780 7584 13796 7648
rect 13860 7584 13866 7648
rect 13550 7583 13866 7584
rect 19852 7648 20168 7649
rect 19852 7584 19858 7648
rect 19922 7584 19938 7648
rect 20002 7584 20018 7648
rect 20082 7584 20098 7648
rect 20162 7584 20168 7648
rect 19852 7583 20168 7584
rect 26154 7648 26470 7649
rect 26154 7584 26160 7648
rect 26224 7584 26240 7648
rect 26304 7584 26320 7648
rect 26384 7584 26400 7648
rect 26464 7584 26470 7648
rect 26154 7583 26470 7584
rect 4097 7104 4413 7105
rect 4097 7040 4103 7104
rect 4167 7040 4183 7104
rect 4247 7040 4263 7104
rect 4327 7040 4343 7104
rect 4407 7040 4413 7104
rect 4097 7039 4413 7040
rect 10399 7104 10715 7105
rect 10399 7040 10405 7104
rect 10469 7040 10485 7104
rect 10549 7040 10565 7104
rect 10629 7040 10645 7104
rect 10709 7040 10715 7104
rect 10399 7039 10715 7040
rect 16701 7104 17017 7105
rect 16701 7040 16707 7104
rect 16771 7040 16787 7104
rect 16851 7040 16867 7104
rect 16931 7040 16947 7104
rect 17011 7040 17017 7104
rect 16701 7039 17017 7040
rect 23003 7104 23319 7105
rect 23003 7040 23009 7104
rect 23073 7040 23089 7104
rect 23153 7040 23169 7104
rect 23233 7040 23249 7104
rect 23313 7040 23319 7104
rect 23003 7039 23319 7040
rect 7248 6560 7564 6561
rect 7248 6496 7254 6560
rect 7318 6496 7334 6560
rect 7398 6496 7414 6560
rect 7478 6496 7494 6560
rect 7558 6496 7564 6560
rect 7248 6495 7564 6496
rect 13550 6560 13866 6561
rect 13550 6496 13556 6560
rect 13620 6496 13636 6560
rect 13700 6496 13716 6560
rect 13780 6496 13796 6560
rect 13860 6496 13866 6560
rect 13550 6495 13866 6496
rect 19852 6560 20168 6561
rect 19852 6496 19858 6560
rect 19922 6496 19938 6560
rect 20002 6496 20018 6560
rect 20082 6496 20098 6560
rect 20162 6496 20168 6560
rect 19852 6495 20168 6496
rect 26154 6560 26470 6561
rect 26154 6496 26160 6560
rect 26224 6496 26240 6560
rect 26304 6496 26320 6560
rect 26384 6496 26400 6560
rect 26464 6496 26470 6560
rect 26154 6495 26470 6496
rect 4097 6016 4413 6017
rect 4097 5952 4103 6016
rect 4167 5952 4183 6016
rect 4247 5952 4263 6016
rect 4327 5952 4343 6016
rect 4407 5952 4413 6016
rect 4097 5951 4413 5952
rect 10399 6016 10715 6017
rect 10399 5952 10405 6016
rect 10469 5952 10485 6016
rect 10549 5952 10565 6016
rect 10629 5952 10645 6016
rect 10709 5952 10715 6016
rect 10399 5951 10715 5952
rect 16701 6016 17017 6017
rect 16701 5952 16707 6016
rect 16771 5952 16787 6016
rect 16851 5952 16867 6016
rect 16931 5952 16947 6016
rect 17011 5952 17017 6016
rect 16701 5951 17017 5952
rect 23003 6016 23319 6017
rect 23003 5952 23009 6016
rect 23073 5952 23089 6016
rect 23153 5952 23169 6016
rect 23233 5952 23249 6016
rect 23313 5952 23319 6016
rect 23003 5951 23319 5952
rect 7248 5472 7564 5473
rect 7248 5408 7254 5472
rect 7318 5408 7334 5472
rect 7398 5408 7414 5472
rect 7478 5408 7494 5472
rect 7558 5408 7564 5472
rect 7248 5407 7564 5408
rect 13550 5472 13866 5473
rect 13550 5408 13556 5472
rect 13620 5408 13636 5472
rect 13700 5408 13716 5472
rect 13780 5408 13796 5472
rect 13860 5408 13866 5472
rect 13550 5407 13866 5408
rect 19852 5472 20168 5473
rect 19852 5408 19858 5472
rect 19922 5408 19938 5472
rect 20002 5408 20018 5472
rect 20082 5408 20098 5472
rect 20162 5408 20168 5472
rect 19852 5407 20168 5408
rect 26154 5472 26470 5473
rect 26154 5408 26160 5472
rect 26224 5408 26240 5472
rect 26304 5408 26320 5472
rect 26384 5408 26400 5472
rect 26464 5408 26470 5472
rect 26154 5407 26470 5408
rect 4097 4928 4413 4929
rect 4097 4864 4103 4928
rect 4167 4864 4183 4928
rect 4247 4864 4263 4928
rect 4327 4864 4343 4928
rect 4407 4864 4413 4928
rect 4097 4863 4413 4864
rect 10399 4928 10715 4929
rect 10399 4864 10405 4928
rect 10469 4864 10485 4928
rect 10549 4864 10565 4928
rect 10629 4864 10645 4928
rect 10709 4864 10715 4928
rect 10399 4863 10715 4864
rect 16701 4928 17017 4929
rect 16701 4864 16707 4928
rect 16771 4864 16787 4928
rect 16851 4864 16867 4928
rect 16931 4864 16947 4928
rect 17011 4864 17017 4928
rect 16701 4863 17017 4864
rect 23003 4928 23319 4929
rect 23003 4864 23009 4928
rect 23073 4864 23089 4928
rect 23153 4864 23169 4928
rect 23233 4864 23249 4928
rect 23313 4864 23319 4928
rect 23003 4863 23319 4864
rect 7248 4384 7564 4385
rect 7248 4320 7254 4384
rect 7318 4320 7334 4384
rect 7398 4320 7414 4384
rect 7478 4320 7494 4384
rect 7558 4320 7564 4384
rect 7248 4319 7564 4320
rect 13550 4384 13866 4385
rect 13550 4320 13556 4384
rect 13620 4320 13636 4384
rect 13700 4320 13716 4384
rect 13780 4320 13796 4384
rect 13860 4320 13866 4384
rect 13550 4319 13866 4320
rect 19852 4384 20168 4385
rect 19852 4320 19858 4384
rect 19922 4320 19938 4384
rect 20002 4320 20018 4384
rect 20082 4320 20098 4384
rect 20162 4320 20168 4384
rect 19852 4319 20168 4320
rect 26154 4384 26470 4385
rect 26154 4320 26160 4384
rect 26224 4320 26240 4384
rect 26304 4320 26320 4384
rect 26384 4320 26400 4384
rect 26464 4320 26470 4384
rect 26154 4319 26470 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 25957 4178 26023 4181
rect 26665 4178 27465 4208
rect 25957 4176 27465 4178
rect 25957 4120 25962 4176
rect 26018 4120 27465 4176
rect 25957 4118 27465 4120
rect 25957 4115 26023 4118
rect 26665 4088 27465 4118
rect 4097 3840 4413 3841
rect 4097 3776 4103 3840
rect 4167 3776 4183 3840
rect 4247 3776 4263 3840
rect 4327 3776 4343 3840
rect 4407 3776 4413 3840
rect 4097 3775 4413 3776
rect 10399 3840 10715 3841
rect 10399 3776 10405 3840
rect 10469 3776 10485 3840
rect 10549 3776 10565 3840
rect 10629 3776 10645 3840
rect 10709 3776 10715 3840
rect 10399 3775 10715 3776
rect 16701 3840 17017 3841
rect 16701 3776 16707 3840
rect 16771 3776 16787 3840
rect 16851 3776 16867 3840
rect 16931 3776 16947 3840
rect 17011 3776 17017 3840
rect 16701 3775 17017 3776
rect 23003 3840 23319 3841
rect 23003 3776 23009 3840
rect 23073 3776 23089 3840
rect 23153 3776 23169 3840
rect 23233 3776 23249 3840
rect 23313 3776 23319 3840
rect 23003 3775 23319 3776
rect 7248 3296 7564 3297
rect 7248 3232 7254 3296
rect 7318 3232 7334 3296
rect 7398 3232 7414 3296
rect 7478 3232 7494 3296
rect 7558 3232 7564 3296
rect 7248 3231 7564 3232
rect 13550 3296 13866 3297
rect 13550 3232 13556 3296
rect 13620 3232 13636 3296
rect 13700 3232 13716 3296
rect 13780 3232 13796 3296
rect 13860 3232 13866 3296
rect 13550 3231 13866 3232
rect 19852 3296 20168 3297
rect 19852 3232 19858 3296
rect 19922 3232 19938 3296
rect 20002 3232 20018 3296
rect 20082 3232 20098 3296
rect 20162 3232 20168 3296
rect 19852 3231 20168 3232
rect 26154 3296 26470 3297
rect 26154 3232 26160 3296
rect 26224 3232 26240 3296
rect 26304 3232 26320 3296
rect 26384 3232 26400 3296
rect 26464 3232 26470 3296
rect 26154 3231 26470 3232
rect 4097 2752 4413 2753
rect 4097 2688 4103 2752
rect 4167 2688 4183 2752
rect 4247 2688 4263 2752
rect 4327 2688 4343 2752
rect 4407 2688 4413 2752
rect 4097 2687 4413 2688
rect 10399 2752 10715 2753
rect 10399 2688 10405 2752
rect 10469 2688 10485 2752
rect 10549 2688 10565 2752
rect 10629 2688 10645 2752
rect 10709 2688 10715 2752
rect 10399 2687 10715 2688
rect 16701 2752 17017 2753
rect 16701 2688 16707 2752
rect 16771 2688 16787 2752
rect 16851 2688 16867 2752
rect 16931 2688 16947 2752
rect 17011 2688 17017 2752
rect 16701 2687 17017 2688
rect 23003 2752 23319 2753
rect 23003 2688 23009 2752
rect 23073 2688 23089 2752
rect 23153 2688 23169 2752
rect 23233 2688 23249 2752
rect 23313 2688 23319 2752
rect 23003 2687 23319 2688
rect 7248 2208 7564 2209
rect 7248 2144 7254 2208
rect 7318 2144 7334 2208
rect 7398 2144 7414 2208
rect 7478 2144 7494 2208
rect 7558 2144 7564 2208
rect 7248 2143 7564 2144
rect 13550 2208 13866 2209
rect 13550 2144 13556 2208
rect 13620 2144 13636 2208
rect 13700 2144 13716 2208
rect 13780 2144 13796 2208
rect 13860 2144 13866 2208
rect 13550 2143 13866 2144
rect 19852 2208 20168 2209
rect 19852 2144 19858 2208
rect 19922 2144 19938 2208
rect 20002 2144 20018 2208
rect 20082 2144 20098 2208
rect 20162 2144 20168 2208
rect 19852 2143 20168 2144
rect 26154 2208 26470 2209
rect 26154 2144 26160 2208
rect 26224 2144 26240 2208
rect 26304 2144 26320 2208
rect 26384 2144 26400 2208
rect 26464 2144 26470 2208
rect 26154 2143 26470 2144
rect 24761 98 24827 101
rect 26665 98 27465 128
rect 24761 96 27465 98
rect 24761 40 24766 96
rect 24822 40 27465 96
rect 24761 38 27465 40
rect 24761 35 24827 38
rect 26665 8 27465 38
<< via3 >>
rect 7254 27228 7318 27232
rect 7254 27172 7258 27228
rect 7258 27172 7314 27228
rect 7314 27172 7318 27228
rect 7254 27168 7318 27172
rect 7334 27228 7398 27232
rect 7334 27172 7338 27228
rect 7338 27172 7394 27228
rect 7394 27172 7398 27228
rect 7334 27168 7398 27172
rect 7414 27228 7478 27232
rect 7414 27172 7418 27228
rect 7418 27172 7474 27228
rect 7474 27172 7478 27228
rect 7414 27168 7478 27172
rect 7494 27228 7558 27232
rect 7494 27172 7498 27228
rect 7498 27172 7554 27228
rect 7554 27172 7558 27228
rect 7494 27168 7558 27172
rect 13556 27228 13620 27232
rect 13556 27172 13560 27228
rect 13560 27172 13616 27228
rect 13616 27172 13620 27228
rect 13556 27168 13620 27172
rect 13636 27228 13700 27232
rect 13636 27172 13640 27228
rect 13640 27172 13696 27228
rect 13696 27172 13700 27228
rect 13636 27168 13700 27172
rect 13716 27228 13780 27232
rect 13716 27172 13720 27228
rect 13720 27172 13776 27228
rect 13776 27172 13780 27228
rect 13716 27168 13780 27172
rect 13796 27228 13860 27232
rect 13796 27172 13800 27228
rect 13800 27172 13856 27228
rect 13856 27172 13860 27228
rect 13796 27168 13860 27172
rect 19858 27228 19922 27232
rect 19858 27172 19862 27228
rect 19862 27172 19918 27228
rect 19918 27172 19922 27228
rect 19858 27168 19922 27172
rect 19938 27228 20002 27232
rect 19938 27172 19942 27228
rect 19942 27172 19998 27228
rect 19998 27172 20002 27228
rect 19938 27168 20002 27172
rect 20018 27228 20082 27232
rect 20018 27172 20022 27228
rect 20022 27172 20078 27228
rect 20078 27172 20082 27228
rect 20018 27168 20082 27172
rect 20098 27228 20162 27232
rect 20098 27172 20102 27228
rect 20102 27172 20158 27228
rect 20158 27172 20162 27228
rect 20098 27168 20162 27172
rect 26160 27228 26224 27232
rect 26160 27172 26164 27228
rect 26164 27172 26220 27228
rect 26220 27172 26224 27228
rect 26160 27168 26224 27172
rect 26240 27228 26304 27232
rect 26240 27172 26244 27228
rect 26244 27172 26300 27228
rect 26300 27172 26304 27228
rect 26240 27168 26304 27172
rect 26320 27228 26384 27232
rect 26320 27172 26324 27228
rect 26324 27172 26380 27228
rect 26380 27172 26384 27228
rect 26320 27168 26384 27172
rect 26400 27228 26464 27232
rect 26400 27172 26404 27228
rect 26404 27172 26460 27228
rect 26460 27172 26464 27228
rect 26400 27168 26464 27172
rect 4103 26684 4167 26688
rect 4103 26628 4107 26684
rect 4107 26628 4163 26684
rect 4163 26628 4167 26684
rect 4103 26624 4167 26628
rect 4183 26684 4247 26688
rect 4183 26628 4187 26684
rect 4187 26628 4243 26684
rect 4243 26628 4247 26684
rect 4183 26624 4247 26628
rect 4263 26684 4327 26688
rect 4263 26628 4267 26684
rect 4267 26628 4323 26684
rect 4323 26628 4327 26684
rect 4263 26624 4327 26628
rect 4343 26684 4407 26688
rect 4343 26628 4347 26684
rect 4347 26628 4403 26684
rect 4403 26628 4407 26684
rect 4343 26624 4407 26628
rect 10405 26684 10469 26688
rect 10405 26628 10409 26684
rect 10409 26628 10465 26684
rect 10465 26628 10469 26684
rect 10405 26624 10469 26628
rect 10485 26684 10549 26688
rect 10485 26628 10489 26684
rect 10489 26628 10545 26684
rect 10545 26628 10549 26684
rect 10485 26624 10549 26628
rect 10565 26684 10629 26688
rect 10565 26628 10569 26684
rect 10569 26628 10625 26684
rect 10625 26628 10629 26684
rect 10565 26624 10629 26628
rect 10645 26684 10709 26688
rect 10645 26628 10649 26684
rect 10649 26628 10705 26684
rect 10705 26628 10709 26684
rect 10645 26624 10709 26628
rect 16707 26684 16771 26688
rect 16707 26628 16711 26684
rect 16711 26628 16767 26684
rect 16767 26628 16771 26684
rect 16707 26624 16771 26628
rect 16787 26684 16851 26688
rect 16787 26628 16791 26684
rect 16791 26628 16847 26684
rect 16847 26628 16851 26684
rect 16787 26624 16851 26628
rect 16867 26684 16931 26688
rect 16867 26628 16871 26684
rect 16871 26628 16927 26684
rect 16927 26628 16931 26684
rect 16867 26624 16931 26628
rect 16947 26684 17011 26688
rect 16947 26628 16951 26684
rect 16951 26628 17007 26684
rect 17007 26628 17011 26684
rect 16947 26624 17011 26628
rect 23009 26684 23073 26688
rect 23009 26628 23013 26684
rect 23013 26628 23069 26684
rect 23069 26628 23073 26684
rect 23009 26624 23073 26628
rect 23089 26684 23153 26688
rect 23089 26628 23093 26684
rect 23093 26628 23149 26684
rect 23149 26628 23153 26684
rect 23089 26624 23153 26628
rect 23169 26684 23233 26688
rect 23169 26628 23173 26684
rect 23173 26628 23229 26684
rect 23229 26628 23233 26684
rect 23169 26624 23233 26628
rect 23249 26684 23313 26688
rect 23249 26628 23253 26684
rect 23253 26628 23309 26684
rect 23309 26628 23313 26684
rect 23249 26624 23313 26628
rect 7254 26140 7318 26144
rect 7254 26084 7258 26140
rect 7258 26084 7314 26140
rect 7314 26084 7318 26140
rect 7254 26080 7318 26084
rect 7334 26140 7398 26144
rect 7334 26084 7338 26140
rect 7338 26084 7394 26140
rect 7394 26084 7398 26140
rect 7334 26080 7398 26084
rect 7414 26140 7478 26144
rect 7414 26084 7418 26140
rect 7418 26084 7474 26140
rect 7474 26084 7478 26140
rect 7414 26080 7478 26084
rect 7494 26140 7558 26144
rect 7494 26084 7498 26140
rect 7498 26084 7554 26140
rect 7554 26084 7558 26140
rect 7494 26080 7558 26084
rect 13556 26140 13620 26144
rect 13556 26084 13560 26140
rect 13560 26084 13616 26140
rect 13616 26084 13620 26140
rect 13556 26080 13620 26084
rect 13636 26140 13700 26144
rect 13636 26084 13640 26140
rect 13640 26084 13696 26140
rect 13696 26084 13700 26140
rect 13636 26080 13700 26084
rect 13716 26140 13780 26144
rect 13716 26084 13720 26140
rect 13720 26084 13776 26140
rect 13776 26084 13780 26140
rect 13716 26080 13780 26084
rect 13796 26140 13860 26144
rect 13796 26084 13800 26140
rect 13800 26084 13856 26140
rect 13856 26084 13860 26140
rect 13796 26080 13860 26084
rect 19858 26140 19922 26144
rect 19858 26084 19862 26140
rect 19862 26084 19918 26140
rect 19918 26084 19922 26140
rect 19858 26080 19922 26084
rect 19938 26140 20002 26144
rect 19938 26084 19942 26140
rect 19942 26084 19998 26140
rect 19998 26084 20002 26140
rect 19938 26080 20002 26084
rect 20018 26140 20082 26144
rect 20018 26084 20022 26140
rect 20022 26084 20078 26140
rect 20078 26084 20082 26140
rect 20018 26080 20082 26084
rect 20098 26140 20162 26144
rect 20098 26084 20102 26140
rect 20102 26084 20158 26140
rect 20158 26084 20162 26140
rect 20098 26080 20162 26084
rect 26160 26140 26224 26144
rect 26160 26084 26164 26140
rect 26164 26084 26220 26140
rect 26220 26084 26224 26140
rect 26160 26080 26224 26084
rect 26240 26140 26304 26144
rect 26240 26084 26244 26140
rect 26244 26084 26300 26140
rect 26300 26084 26304 26140
rect 26240 26080 26304 26084
rect 26320 26140 26384 26144
rect 26320 26084 26324 26140
rect 26324 26084 26380 26140
rect 26380 26084 26384 26140
rect 26320 26080 26384 26084
rect 26400 26140 26464 26144
rect 26400 26084 26404 26140
rect 26404 26084 26460 26140
rect 26460 26084 26464 26140
rect 26400 26080 26464 26084
rect 4103 25596 4167 25600
rect 4103 25540 4107 25596
rect 4107 25540 4163 25596
rect 4163 25540 4167 25596
rect 4103 25536 4167 25540
rect 4183 25596 4247 25600
rect 4183 25540 4187 25596
rect 4187 25540 4243 25596
rect 4243 25540 4247 25596
rect 4183 25536 4247 25540
rect 4263 25596 4327 25600
rect 4263 25540 4267 25596
rect 4267 25540 4323 25596
rect 4323 25540 4327 25596
rect 4263 25536 4327 25540
rect 4343 25596 4407 25600
rect 4343 25540 4347 25596
rect 4347 25540 4403 25596
rect 4403 25540 4407 25596
rect 4343 25536 4407 25540
rect 10405 25596 10469 25600
rect 10405 25540 10409 25596
rect 10409 25540 10465 25596
rect 10465 25540 10469 25596
rect 10405 25536 10469 25540
rect 10485 25596 10549 25600
rect 10485 25540 10489 25596
rect 10489 25540 10545 25596
rect 10545 25540 10549 25596
rect 10485 25536 10549 25540
rect 10565 25596 10629 25600
rect 10565 25540 10569 25596
rect 10569 25540 10625 25596
rect 10625 25540 10629 25596
rect 10565 25536 10629 25540
rect 10645 25596 10709 25600
rect 10645 25540 10649 25596
rect 10649 25540 10705 25596
rect 10705 25540 10709 25596
rect 10645 25536 10709 25540
rect 16707 25596 16771 25600
rect 16707 25540 16711 25596
rect 16711 25540 16767 25596
rect 16767 25540 16771 25596
rect 16707 25536 16771 25540
rect 16787 25596 16851 25600
rect 16787 25540 16791 25596
rect 16791 25540 16847 25596
rect 16847 25540 16851 25596
rect 16787 25536 16851 25540
rect 16867 25596 16931 25600
rect 16867 25540 16871 25596
rect 16871 25540 16927 25596
rect 16927 25540 16931 25596
rect 16867 25536 16931 25540
rect 16947 25596 17011 25600
rect 16947 25540 16951 25596
rect 16951 25540 17007 25596
rect 17007 25540 17011 25596
rect 16947 25536 17011 25540
rect 23009 25596 23073 25600
rect 23009 25540 23013 25596
rect 23013 25540 23069 25596
rect 23069 25540 23073 25596
rect 23009 25536 23073 25540
rect 23089 25596 23153 25600
rect 23089 25540 23093 25596
rect 23093 25540 23149 25596
rect 23149 25540 23153 25596
rect 23089 25536 23153 25540
rect 23169 25596 23233 25600
rect 23169 25540 23173 25596
rect 23173 25540 23229 25596
rect 23229 25540 23233 25596
rect 23169 25536 23233 25540
rect 23249 25596 23313 25600
rect 23249 25540 23253 25596
rect 23253 25540 23309 25596
rect 23309 25540 23313 25596
rect 23249 25536 23313 25540
rect 7254 25052 7318 25056
rect 7254 24996 7258 25052
rect 7258 24996 7314 25052
rect 7314 24996 7318 25052
rect 7254 24992 7318 24996
rect 7334 25052 7398 25056
rect 7334 24996 7338 25052
rect 7338 24996 7394 25052
rect 7394 24996 7398 25052
rect 7334 24992 7398 24996
rect 7414 25052 7478 25056
rect 7414 24996 7418 25052
rect 7418 24996 7474 25052
rect 7474 24996 7478 25052
rect 7414 24992 7478 24996
rect 7494 25052 7558 25056
rect 7494 24996 7498 25052
rect 7498 24996 7554 25052
rect 7554 24996 7558 25052
rect 7494 24992 7558 24996
rect 13556 25052 13620 25056
rect 13556 24996 13560 25052
rect 13560 24996 13616 25052
rect 13616 24996 13620 25052
rect 13556 24992 13620 24996
rect 13636 25052 13700 25056
rect 13636 24996 13640 25052
rect 13640 24996 13696 25052
rect 13696 24996 13700 25052
rect 13636 24992 13700 24996
rect 13716 25052 13780 25056
rect 13716 24996 13720 25052
rect 13720 24996 13776 25052
rect 13776 24996 13780 25052
rect 13716 24992 13780 24996
rect 13796 25052 13860 25056
rect 13796 24996 13800 25052
rect 13800 24996 13856 25052
rect 13856 24996 13860 25052
rect 13796 24992 13860 24996
rect 19858 25052 19922 25056
rect 19858 24996 19862 25052
rect 19862 24996 19918 25052
rect 19918 24996 19922 25052
rect 19858 24992 19922 24996
rect 19938 25052 20002 25056
rect 19938 24996 19942 25052
rect 19942 24996 19998 25052
rect 19998 24996 20002 25052
rect 19938 24992 20002 24996
rect 20018 25052 20082 25056
rect 20018 24996 20022 25052
rect 20022 24996 20078 25052
rect 20078 24996 20082 25052
rect 20018 24992 20082 24996
rect 20098 25052 20162 25056
rect 20098 24996 20102 25052
rect 20102 24996 20158 25052
rect 20158 24996 20162 25052
rect 20098 24992 20162 24996
rect 26160 25052 26224 25056
rect 26160 24996 26164 25052
rect 26164 24996 26220 25052
rect 26220 24996 26224 25052
rect 26160 24992 26224 24996
rect 26240 25052 26304 25056
rect 26240 24996 26244 25052
rect 26244 24996 26300 25052
rect 26300 24996 26304 25052
rect 26240 24992 26304 24996
rect 26320 25052 26384 25056
rect 26320 24996 26324 25052
rect 26324 24996 26380 25052
rect 26380 24996 26384 25052
rect 26320 24992 26384 24996
rect 26400 25052 26464 25056
rect 26400 24996 26404 25052
rect 26404 24996 26460 25052
rect 26460 24996 26464 25052
rect 26400 24992 26464 24996
rect 6500 24712 6564 24716
rect 6500 24656 6514 24712
rect 6514 24656 6564 24712
rect 6500 24652 6564 24656
rect 4103 24508 4167 24512
rect 4103 24452 4107 24508
rect 4107 24452 4163 24508
rect 4163 24452 4167 24508
rect 4103 24448 4167 24452
rect 4183 24508 4247 24512
rect 4183 24452 4187 24508
rect 4187 24452 4243 24508
rect 4243 24452 4247 24508
rect 4183 24448 4247 24452
rect 4263 24508 4327 24512
rect 4263 24452 4267 24508
rect 4267 24452 4323 24508
rect 4323 24452 4327 24508
rect 4263 24448 4327 24452
rect 4343 24508 4407 24512
rect 4343 24452 4347 24508
rect 4347 24452 4403 24508
rect 4403 24452 4407 24508
rect 4343 24448 4407 24452
rect 10405 24508 10469 24512
rect 10405 24452 10409 24508
rect 10409 24452 10465 24508
rect 10465 24452 10469 24508
rect 10405 24448 10469 24452
rect 10485 24508 10549 24512
rect 10485 24452 10489 24508
rect 10489 24452 10545 24508
rect 10545 24452 10549 24508
rect 10485 24448 10549 24452
rect 10565 24508 10629 24512
rect 10565 24452 10569 24508
rect 10569 24452 10625 24508
rect 10625 24452 10629 24508
rect 10565 24448 10629 24452
rect 10645 24508 10709 24512
rect 10645 24452 10649 24508
rect 10649 24452 10705 24508
rect 10705 24452 10709 24508
rect 10645 24448 10709 24452
rect 16707 24508 16771 24512
rect 16707 24452 16711 24508
rect 16711 24452 16767 24508
rect 16767 24452 16771 24508
rect 16707 24448 16771 24452
rect 16787 24508 16851 24512
rect 16787 24452 16791 24508
rect 16791 24452 16847 24508
rect 16847 24452 16851 24508
rect 16787 24448 16851 24452
rect 16867 24508 16931 24512
rect 16867 24452 16871 24508
rect 16871 24452 16927 24508
rect 16927 24452 16931 24508
rect 16867 24448 16931 24452
rect 16947 24508 17011 24512
rect 16947 24452 16951 24508
rect 16951 24452 17007 24508
rect 17007 24452 17011 24508
rect 16947 24448 17011 24452
rect 23009 24508 23073 24512
rect 23009 24452 23013 24508
rect 23013 24452 23069 24508
rect 23069 24452 23073 24508
rect 23009 24448 23073 24452
rect 23089 24508 23153 24512
rect 23089 24452 23093 24508
rect 23093 24452 23149 24508
rect 23149 24452 23153 24508
rect 23089 24448 23153 24452
rect 23169 24508 23233 24512
rect 23169 24452 23173 24508
rect 23173 24452 23229 24508
rect 23229 24452 23233 24508
rect 23169 24448 23233 24452
rect 23249 24508 23313 24512
rect 23249 24452 23253 24508
rect 23253 24452 23309 24508
rect 23309 24452 23313 24508
rect 23249 24448 23313 24452
rect 7254 23964 7318 23968
rect 7254 23908 7258 23964
rect 7258 23908 7314 23964
rect 7314 23908 7318 23964
rect 7254 23904 7318 23908
rect 7334 23964 7398 23968
rect 7334 23908 7338 23964
rect 7338 23908 7394 23964
rect 7394 23908 7398 23964
rect 7334 23904 7398 23908
rect 7414 23964 7478 23968
rect 7414 23908 7418 23964
rect 7418 23908 7474 23964
rect 7474 23908 7478 23964
rect 7414 23904 7478 23908
rect 7494 23964 7558 23968
rect 7494 23908 7498 23964
rect 7498 23908 7554 23964
rect 7554 23908 7558 23964
rect 7494 23904 7558 23908
rect 13556 23964 13620 23968
rect 13556 23908 13560 23964
rect 13560 23908 13616 23964
rect 13616 23908 13620 23964
rect 13556 23904 13620 23908
rect 13636 23964 13700 23968
rect 13636 23908 13640 23964
rect 13640 23908 13696 23964
rect 13696 23908 13700 23964
rect 13636 23904 13700 23908
rect 13716 23964 13780 23968
rect 13716 23908 13720 23964
rect 13720 23908 13776 23964
rect 13776 23908 13780 23964
rect 13716 23904 13780 23908
rect 13796 23964 13860 23968
rect 13796 23908 13800 23964
rect 13800 23908 13856 23964
rect 13856 23908 13860 23964
rect 13796 23904 13860 23908
rect 19858 23964 19922 23968
rect 19858 23908 19862 23964
rect 19862 23908 19918 23964
rect 19918 23908 19922 23964
rect 19858 23904 19922 23908
rect 19938 23964 20002 23968
rect 19938 23908 19942 23964
rect 19942 23908 19998 23964
rect 19998 23908 20002 23964
rect 19938 23904 20002 23908
rect 20018 23964 20082 23968
rect 20018 23908 20022 23964
rect 20022 23908 20078 23964
rect 20078 23908 20082 23964
rect 20018 23904 20082 23908
rect 20098 23964 20162 23968
rect 20098 23908 20102 23964
rect 20102 23908 20158 23964
rect 20158 23908 20162 23964
rect 20098 23904 20162 23908
rect 26160 23964 26224 23968
rect 26160 23908 26164 23964
rect 26164 23908 26220 23964
rect 26220 23908 26224 23964
rect 26160 23904 26224 23908
rect 26240 23964 26304 23968
rect 26240 23908 26244 23964
rect 26244 23908 26300 23964
rect 26300 23908 26304 23964
rect 26240 23904 26304 23908
rect 26320 23964 26384 23968
rect 26320 23908 26324 23964
rect 26324 23908 26380 23964
rect 26380 23908 26384 23964
rect 26320 23904 26384 23908
rect 26400 23964 26464 23968
rect 26400 23908 26404 23964
rect 26404 23908 26460 23964
rect 26460 23908 26464 23964
rect 26400 23904 26464 23908
rect 4103 23420 4167 23424
rect 4103 23364 4107 23420
rect 4107 23364 4163 23420
rect 4163 23364 4167 23420
rect 4103 23360 4167 23364
rect 4183 23420 4247 23424
rect 4183 23364 4187 23420
rect 4187 23364 4243 23420
rect 4243 23364 4247 23420
rect 4183 23360 4247 23364
rect 4263 23420 4327 23424
rect 4263 23364 4267 23420
rect 4267 23364 4323 23420
rect 4323 23364 4327 23420
rect 4263 23360 4327 23364
rect 4343 23420 4407 23424
rect 4343 23364 4347 23420
rect 4347 23364 4403 23420
rect 4403 23364 4407 23420
rect 4343 23360 4407 23364
rect 10405 23420 10469 23424
rect 10405 23364 10409 23420
rect 10409 23364 10465 23420
rect 10465 23364 10469 23420
rect 10405 23360 10469 23364
rect 10485 23420 10549 23424
rect 10485 23364 10489 23420
rect 10489 23364 10545 23420
rect 10545 23364 10549 23420
rect 10485 23360 10549 23364
rect 10565 23420 10629 23424
rect 10565 23364 10569 23420
rect 10569 23364 10625 23420
rect 10625 23364 10629 23420
rect 10565 23360 10629 23364
rect 10645 23420 10709 23424
rect 10645 23364 10649 23420
rect 10649 23364 10705 23420
rect 10705 23364 10709 23420
rect 10645 23360 10709 23364
rect 16707 23420 16771 23424
rect 16707 23364 16711 23420
rect 16711 23364 16767 23420
rect 16767 23364 16771 23420
rect 16707 23360 16771 23364
rect 16787 23420 16851 23424
rect 16787 23364 16791 23420
rect 16791 23364 16847 23420
rect 16847 23364 16851 23420
rect 16787 23360 16851 23364
rect 16867 23420 16931 23424
rect 16867 23364 16871 23420
rect 16871 23364 16927 23420
rect 16927 23364 16931 23420
rect 16867 23360 16931 23364
rect 16947 23420 17011 23424
rect 16947 23364 16951 23420
rect 16951 23364 17007 23420
rect 17007 23364 17011 23420
rect 16947 23360 17011 23364
rect 23009 23420 23073 23424
rect 23009 23364 23013 23420
rect 23013 23364 23069 23420
rect 23069 23364 23073 23420
rect 23009 23360 23073 23364
rect 23089 23420 23153 23424
rect 23089 23364 23093 23420
rect 23093 23364 23149 23420
rect 23149 23364 23153 23420
rect 23089 23360 23153 23364
rect 23169 23420 23233 23424
rect 23169 23364 23173 23420
rect 23173 23364 23229 23420
rect 23229 23364 23233 23420
rect 23169 23360 23233 23364
rect 23249 23420 23313 23424
rect 23249 23364 23253 23420
rect 23253 23364 23309 23420
rect 23309 23364 23313 23420
rect 23249 23360 23313 23364
rect 7254 22876 7318 22880
rect 7254 22820 7258 22876
rect 7258 22820 7314 22876
rect 7314 22820 7318 22876
rect 7254 22816 7318 22820
rect 7334 22876 7398 22880
rect 7334 22820 7338 22876
rect 7338 22820 7394 22876
rect 7394 22820 7398 22876
rect 7334 22816 7398 22820
rect 7414 22876 7478 22880
rect 7414 22820 7418 22876
rect 7418 22820 7474 22876
rect 7474 22820 7478 22876
rect 7414 22816 7478 22820
rect 7494 22876 7558 22880
rect 7494 22820 7498 22876
rect 7498 22820 7554 22876
rect 7554 22820 7558 22876
rect 7494 22816 7558 22820
rect 13556 22876 13620 22880
rect 13556 22820 13560 22876
rect 13560 22820 13616 22876
rect 13616 22820 13620 22876
rect 13556 22816 13620 22820
rect 13636 22876 13700 22880
rect 13636 22820 13640 22876
rect 13640 22820 13696 22876
rect 13696 22820 13700 22876
rect 13636 22816 13700 22820
rect 13716 22876 13780 22880
rect 13716 22820 13720 22876
rect 13720 22820 13776 22876
rect 13776 22820 13780 22876
rect 13716 22816 13780 22820
rect 13796 22876 13860 22880
rect 13796 22820 13800 22876
rect 13800 22820 13856 22876
rect 13856 22820 13860 22876
rect 13796 22816 13860 22820
rect 19858 22876 19922 22880
rect 19858 22820 19862 22876
rect 19862 22820 19918 22876
rect 19918 22820 19922 22876
rect 19858 22816 19922 22820
rect 19938 22876 20002 22880
rect 19938 22820 19942 22876
rect 19942 22820 19998 22876
rect 19998 22820 20002 22876
rect 19938 22816 20002 22820
rect 20018 22876 20082 22880
rect 20018 22820 20022 22876
rect 20022 22820 20078 22876
rect 20078 22820 20082 22876
rect 20018 22816 20082 22820
rect 20098 22876 20162 22880
rect 20098 22820 20102 22876
rect 20102 22820 20158 22876
rect 20158 22820 20162 22876
rect 20098 22816 20162 22820
rect 26160 22876 26224 22880
rect 26160 22820 26164 22876
rect 26164 22820 26220 22876
rect 26220 22820 26224 22876
rect 26160 22816 26224 22820
rect 26240 22876 26304 22880
rect 26240 22820 26244 22876
rect 26244 22820 26300 22876
rect 26300 22820 26304 22876
rect 26240 22816 26304 22820
rect 26320 22876 26384 22880
rect 26320 22820 26324 22876
rect 26324 22820 26380 22876
rect 26380 22820 26384 22876
rect 26320 22816 26384 22820
rect 26400 22876 26464 22880
rect 26400 22820 26404 22876
rect 26404 22820 26460 22876
rect 26460 22820 26464 22876
rect 26400 22816 26464 22820
rect 4103 22332 4167 22336
rect 4103 22276 4107 22332
rect 4107 22276 4163 22332
rect 4163 22276 4167 22332
rect 4103 22272 4167 22276
rect 4183 22332 4247 22336
rect 4183 22276 4187 22332
rect 4187 22276 4243 22332
rect 4243 22276 4247 22332
rect 4183 22272 4247 22276
rect 4263 22332 4327 22336
rect 4263 22276 4267 22332
rect 4267 22276 4323 22332
rect 4323 22276 4327 22332
rect 4263 22272 4327 22276
rect 4343 22332 4407 22336
rect 4343 22276 4347 22332
rect 4347 22276 4403 22332
rect 4403 22276 4407 22332
rect 4343 22272 4407 22276
rect 10405 22332 10469 22336
rect 10405 22276 10409 22332
rect 10409 22276 10465 22332
rect 10465 22276 10469 22332
rect 10405 22272 10469 22276
rect 10485 22332 10549 22336
rect 10485 22276 10489 22332
rect 10489 22276 10545 22332
rect 10545 22276 10549 22332
rect 10485 22272 10549 22276
rect 10565 22332 10629 22336
rect 10565 22276 10569 22332
rect 10569 22276 10625 22332
rect 10625 22276 10629 22332
rect 10565 22272 10629 22276
rect 10645 22332 10709 22336
rect 10645 22276 10649 22332
rect 10649 22276 10705 22332
rect 10705 22276 10709 22332
rect 10645 22272 10709 22276
rect 16707 22332 16771 22336
rect 16707 22276 16711 22332
rect 16711 22276 16767 22332
rect 16767 22276 16771 22332
rect 16707 22272 16771 22276
rect 16787 22332 16851 22336
rect 16787 22276 16791 22332
rect 16791 22276 16847 22332
rect 16847 22276 16851 22332
rect 16787 22272 16851 22276
rect 16867 22332 16931 22336
rect 16867 22276 16871 22332
rect 16871 22276 16927 22332
rect 16927 22276 16931 22332
rect 16867 22272 16931 22276
rect 16947 22332 17011 22336
rect 16947 22276 16951 22332
rect 16951 22276 17007 22332
rect 17007 22276 17011 22332
rect 16947 22272 17011 22276
rect 23009 22332 23073 22336
rect 23009 22276 23013 22332
rect 23013 22276 23069 22332
rect 23069 22276 23073 22332
rect 23009 22272 23073 22276
rect 23089 22332 23153 22336
rect 23089 22276 23093 22332
rect 23093 22276 23149 22332
rect 23149 22276 23153 22332
rect 23089 22272 23153 22276
rect 23169 22332 23233 22336
rect 23169 22276 23173 22332
rect 23173 22276 23229 22332
rect 23229 22276 23233 22332
rect 23169 22272 23233 22276
rect 23249 22332 23313 22336
rect 23249 22276 23253 22332
rect 23253 22276 23309 22332
rect 23309 22276 23313 22332
rect 23249 22272 23313 22276
rect 7254 21788 7318 21792
rect 7254 21732 7258 21788
rect 7258 21732 7314 21788
rect 7314 21732 7318 21788
rect 7254 21728 7318 21732
rect 7334 21788 7398 21792
rect 7334 21732 7338 21788
rect 7338 21732 7394 21788
rect 7394 21732 7398 21788
rect 7334 21728 7398 21732
rect 7414 21788 7478 21792
rect 7414 21732 7418 21788
rect 7418 21732 7474 21788
rect 7474 21732 7478 21788
rect 7414 21728 7478 21732
rect 7494 21788 7558 21792
rect 7494 21732 7498 21788
rect 7498 21732 7554 21788
rect 7554 21732 7558 21788
rect 7494 21728 7558 21732
rect 13556 21788 13620 21792
rect 13556 21732 13560 21788
rect 13560 21732 13616 21788
rect 13616 21732 13620 21788
rect 13556 21728 13620 21732
rect 13636 21788 13700 21792
rect 13636 21732 13640 21788
rect 13640 21732 13696 21788
rect 13696 21732 13700 21788
rect 13636 21728 13700 21732
rect 13716 21788 13780 21792
rect 13716 21732 13720 21788
rect 13720 21732 13776 21788
rect 13776 21732 13780 21788
rect 13716 21728 13780 21732
rect 13796 21788 13860 21792
rect 13796 21732 13800 21788
rect 13800 21732 13856 21788
rect 13856 21732 13860 21788
rect 13796 21728 13860 21732
rect 19858 21788 19922 21792
rect 19858 21732 19862 21788
rect 19862 21732 19918 21788
rect 19918 21732 19922 21788
rect 19858 21728 19922 21732
rect 19938 21788 20002 21792
rect 19938 21732 19942 21788
rect 19942 21732 19998 21788
rect 19998 21732 20002 21788
rect 19938 21728 20002 21732
rect 20018 21788 20082 21792
rect 20018 21732 20022 21788
rect 20022 21732 20078 21788
rect 20078 21732 20082 21788
rect 20018 21728 20082 21732
rect 20098 21788 20162 21792
rect 20098 21732 20102 21788
rect 20102 21732 20158 21788
rect 20158 21732 20162 21788
rect 20098 21728 20162 21732
rect 26160 21788 26224 21792
rect 26160 21732 26164 21788
rect 26164 21732 26220 21788
rect 26220 21732 26224 21788
rect 26160 21728 26224 21732
rect 26240 21788 26304 21792
rect 26240 21732 26244 21788
rect 26244 21732 26300 21788
rect 26300 21732 26304 21788
rect 26240 21728 26304 21732
rect 26320 21788 26384 21792
rect 26320 21732 26324 21788
rect 26324 21732 26380 21788
rect 26380 21732 26384 21788
rect 26320 21728 26384 21732
rect 26400 21788 26464 21792
rect 26400 21732 26404 21788
rect 26404 21732 26460 21788
rect 26460 21732 26464 21788
rect 26400 21728 26464 21732
rect 4103 21244 4167 21248
rect 4103 21188 4107 21244
rect 4107 21188 4163 21244
rect 4163 21188 4167 21244
rect 4103 21184 4167 21188
rect 4183 21244 4247 21248
rect 4183 21188 4187 21244
rect 4187 21188 4243 21244
rect 4243 21188 4247 21244
rect 4183 21184 4247 21188
rect 4263 21244 4327 21248
rect 4263 21188 4267 21244
rect 4267 21188 4323 21244
rect 4323 21188 4327 21244
rect 4263 21184 4327 21188
rect 4343 21244 4407 21248
rect 4343 21188 4347 21244
rect 4347 21188 4403 21244
rect 4403 21188 4407 21244
rect 4343 21184 4407 21188
rect 10405 21244 10469 21248
rect 10405 21188 10409 21244
rect 10409 21188 10465 21244
rect 10465 21188 10469 21244
rect 10405 21184 10469 21188
rect 10485 21244 10549 21248
rect 10485 21188 10489 21244
rect 10489 21188 10545 21244
rect 10545 21188 10549 21244
rect 10485 21184 10549 21188
rect 10565 21244 10629 21248
rect 10565 21188 10569 21244
rect 10569 21188 10625 21244
rect 10625 21188 10629 21244
rect 10565 21184 10629 21188
rect 10645 21244 10709 21248
rect 10645 21188 10649 21244
rect 10649 21188 10705 21244
rect 10705 21188 10709 21244
rect 10645 21184 10709 21188
rect 16707 21244 16771 21248
rect 16707 21188 16711 21244
rect 16711 21188 16767 21244
rect 16767 21188 16771 21244
rect 16707 21184 16771 21188
rect 16787 21244 16851 21248
rect 16787 21188 16791 21244
rect 16791 21188 16847 21244
rect 16847 21188 16851 21244
rect 16787 21184 16851 21188
rect 16867 21244 16931 21248
rect 16867 21188 16871 21244
rect 16871 21188 16927 21244
rect 16927 21188 16931 21244
rect 16867 21184 16931 21188
rect 16947 21244 17011 21248
rect 16947 21188 16951 21244
rect 16951 21188 17007 21244
rect 17007 21188 17011 21244
rect 16947 21184 17011 21188
rect 23009 21244 23073 21248
rect 23009 21188 23013 21244
rect 23013 21188 23069 21244
rect 23069 21188 23073 21244
rect 23009 21184 23073 21188
rect 23089 21244 23153 21248
rect 23089 21188 23093 21244
rect 23093 21188 23149 21244
rect 23149 21188 23153 21244
rect 23089 21184 23153 21188
rect 23169 21244 23233 21248
rect 23169 21188 23173 21244
rect 23173 21188 23229 21244
rect 23229 21188 23233 21244
rect 23169 21184 23233 21188
rect 23249 21244 23313 21248
rect 23249 21188 23253 21244
rect 23253 21188 23309 21244
rect 23309 21188 23313 21244
rect 23249 21184 23313 21188
rect 7254 20700 7318 20704
rect 7254 20644 7258 20700
rect 7258 20644 7314 20700
rect 7314 20644 7318 20700
rect 7254 20640 7318 20644
rect 7334 20700 7398 20704
rect 7334 20644 7338 20700
rect 7338 20644 7394 20700
rect 7394 20644 7398 20700
rect 7334 20640 7398 20644
rect 7414 20700 7478 20704
rect 7414 20644 7418 20700
rect 7418 20644 7474 20700
rect 7474 20644 7478 20700
rect 7414 20640 7478 20644
rect 7494 20700 7558 20704
rect 7494 20644 7498 20700
rect 7498 20644 7554 20700
rect 7554 20644 7558 20700
rect 7494 20640 7558 20644
rect 13556 20700 13620 20704
rect 13556 20644 13560 20700
rect 13560 20644 13616 20700
rect 13616 20644 13620 20700
rect 13556 20640 13620 20644
rect 13636 20700 13700 20704
rect 13636 20644 13640 20700
rect 13640 20644 13696 20700
rect 13696 20644 13700 20700
rect 13636 20640 13700 20644
rect 13716 20700 13780 20704
rect 13716 20644 13720 20700
rect 13720 20644 13776 20700
rect 13776 20644 13780 20700
rect 13716 20640 13780 20644
rect 13796 20700 13860 20704
rect 13796 20644 13800 20700
rect 13800 20644 13856 20700
rect 13856 20644 13860 20700
rect 13796 20640 13860 20644
rect 19858 20700 19922 20704
rect 19858 20644 19862 20700
rect 19862 20644 19918 20700
rect 19918 20644 19922 20700
rect 19858 20640 19922 20644
rect 19938 20700 20002 20704
rect 19938 20644 19942 20700
rect 19942 20644 19998 20700
rect 19998 20644 20002 20700
rect 19938 20640 20002 20644
rect 20018 20700 20082 20704
rect 20018 20644 20022 20700
rect 20022 20644 20078 20700
rect 20078 20644 20082 20700
rect 20018 20640 20082 20644
rect 20098 20700 20162 20704
rect 20098 20644 20102 20700
rect 20102 20644 20158 20700
rect 20158 20644 20162 20700
rect 20098 20640 20162 20644
rect 26160 20700 26224 20704
rect 26160 20644 26164 20700
rect 26164 20644 26220 20700
rect 26220 20644 26224 20700
rect 26160 20640 26224 20644
rect 26240 20700 26304 20704
rect 26240 20644 26244 20700
rect 26244 20644 26300 20700
rect 26300 20644 26304 20700
rect 26240 20640 26304 20644
rect 26320 20700 26384 20704
rect 26320 20644 26324 20700
rect 26324 20644 26380 20700
rect 26380 20644 26384 20700
rect 26320 20640 26384 20644
rect 26400 20700 26464 20704
rect 26400 20644 26404 20700
rect 26404 20644 26460 20700
rect 26460 20644 26464 20700
rect 26400 20640 26464 20644
rect 4103 20156 4167 20160
rect 4103 20100 4107 20156
rect 4107 20100 4163 20156
rect 4163 20100 4167 20156
rect 4103 20096 4167 20100
rect 4183 20156 4247 20160
rect 4183 20100 4187 20156
rect 4187 20100 4243 20156
rect 4243 20100 4247 20156
rect 4183 20096 4247 20100
rect 4263 20156 4327 20160
rect 4263 20100 4267 20156
rect 4267 20100 4323 20156
rect 4323 20100 4327 20156
rect 4263 20096 4327 20100
rect 4343 20156 4407 20160
rect 4343 20100 4347 20156
rect 4347 20100 4403 20156
rect 4403 20100 4407 20156
rect 4343 20096 4407 20100
rect 10405 20156 10469 20160
rect 10405 20100 10409 20156
rect 10409 20100 10465 20156
rect 10465 20100 10469 20156
rect 10405 20096 10469 20100
rect 10485 20156 10549 20160
rect 10485 20100 10489 20156
rect 10489 20100 10545 20156
rect 10545 20100 10549 20156
rect 10485 20096 10549 20100
rect 10565 20156 10629 20160
rect 10565 20100 10569 20156
rect 10569 20100 10625 20156
rect 10625 20100 10629 20156
rect 10565 20096 10629 20100
rect 10645 20156 10709 20160
rect 10645 20100 10649 20156
rect 10649 20100 10705 20156
rect 10705 20100 10709 20156
rect 10645 20096 10709 20100
rect 16707 20156 16771 20160
rect 16707 20100 16711 20156
rect 16711 20100 16767 20156
rect 16767 20100 16771 20156
rect 16707 20096 16771 20100
rect 16787 20156 16851 20160
rect 16787 20100 16791 20156
rect 16791 20100 16847 20156
rect 16847 20100 16851 20156
rect 16787 20096 16851 20100
rect 16867 20156 16931 20160
rect 16867 20100 16871 20156
rect 16871 20100 16927 20156
rect 16927 20100 16931 20156
rect 16867 20096 16931 20100
rect 16947 20156 17011 20160
rect 16947 20100 16951 20156
rect 16951 20100 17007 20156
rect 17007 20100 17011 20156
rect 16947 20096 17011 20100
rect 23009 20156 23073 20160
rect 23009 20100 23013 20156
rect 23013 20100 23069 20156
rect 23069 20100 23073 20156
rect 23009 20096 23073 20100
rect 23089 20156 23153 20160
rect 23089 20100 23093 20156
rect 23093 20100 23149 20156
rect 23149 20100 23153 20156
rect 23089 20096 23153 20100
rect 23169 20156 23233 20160
rect 23169 20100 23173 20156
rect 23173 20100 23229 20156
rect 23229 20100 23233 20156
rect 23169 20096 23233 20100
rect 23249 20156 23313 20160
rect 23249 20100 23253 20156
rect 23253 20100 23309 20156
rect 23309 20100 23313 20156
rect 23249 20096 23313 20100
rect 7254 19612 7318 19616
rect 7254 19556 7258 19612
rect 7258 19556 7314 19612
rect 7314 19556 7318 19612
rect 7254 19552 7318 19556
rect 7334 19612 7398 19616
rect 7334 19556 7338 19612
rect 7338 19556 7394 19612
rect 7394 19556 7398 19612
rect 7334 19552 7398 19556
rect 7414 19612 7478 19616
rect 7414 19556 7418 19612
rect 7418 19556 7474 19612
rect 7474 19556 7478 19612
rect 7414 19552 7478 19556
rect 7494 19612 7558 19616
rect 7494 19556 7498 19612
rect 7498 19556 7554 19612
rect 7554 19556 7558 19612
rect 7494 19552 7558 19556
rect 13556 19612 13620 19616
rect 13556 19556 13560 19612
rect 13560 19556 13616 19612
rect 13616 19556 13620 19612
rect 13556 19552 13620 19556
rect 13636 19612 13700 19616
rect 13636 19556 13640 19612
rect 13640 19556 13696 19612
rect 13696 19556 13700 19612
rect 13636 19552 13700 19556
rect 13716 19612 13780 19616
rect 13716 19556 13720 19612
rect 13720 19556 13776 19612
rect 13776 19556 13780 19612
rect 13716 19552 13780 19556
rect 13796 19612 13860 19616
rect 13796 19556 13800 19612
rect 13800 19556 13856 19612
rect 13856 19556 13860 19612
rect 13796 19552 13860 19556
rect 19858 19612 19922 19616
rect 19858 19556 19862 19612
rect 19862 19556 19918 19612
rect 19918 19556 19922 19612
rect 19858 19552 19922 19556
rect 19938 19612 20002 19616
rect 19938 19556 19942 19612
rect 19942 19556 19998 19612
rect 19998 19556 20002 19612
rect 19938 19552 20002 19556
rect 20018 19612 20082 19616
rect 20018 19556 20022 19612
rect 20022 19556 20078 19612
rect 20078 19556 20082 19612
rect 20018 19552 20082 19556
rect 20098 19612 20162 19616
rect 20098 19556 20102 19612
rect 20102 19556 20158 19612
rect 20158 19556 20162 19612
rect 20098 19552 20162 19556
rect 26160 19612 26224 19616
rect 26160 19556 26164 19612
rect 26164 19556 26220 19612
rect 26220 19556 26224 19612
rect 26160 19552 26224 19556
rect 26240 19612 26304 19616
rect 26240 19556 26244 19612
rect 26244 19556 26300 19612
rect 26300 19556 26304 19612
rect 26240 19552 26304 19556
rect 26320 19612 26384 19616
rect 26320 19556 26324 19612
rect 26324 19556 26380 19612
rect 26380 19556 26384 19612
rect 26320 19552 26384 19556
rect 26400 19612 26464 19616
rect 26400 19556 26404 19612
rect 26404 19556 26460 19612
rect 26460 19556 26464 19612
rect 26400 19552 26464 19556
rect 4103 19068 4167 19072
rect 4103 19012 4107 19068
rect 4107 19012 4163 19068
rect 4163 19012 4167 19068
rect 4103 19008 4167 19012
rect 4183 19068 4247 19072
rect 4183 19012 4187 19068
rect 4187 19012 4243 19068
rect 4243 19012 4247 19068
rect 4183 19008 4247 19012
rect 4263 19068 4327 19072
rect 4263 19012 4267 19068
rect 4267 19012 4323 19068
rect 4323 19012 4327 19068
rect 4263 19008 4327 19012
rect 4343 19068 4407 19072
rect 4343 19012 4347 19068
rect 4347 19012 4403 19068
rect 4403 19012 4407 19068
rect 4343 19008 4407 19012
rect 10405 19068 10469 19072
rect 10405 19012 10409 19068
rect 10409 19012 10465 19068
rect 10465 19012 10469 19068
rect 10405 19008 10469 19012
rect 10485 19068 10549 19072
rect 10485 19012 10489 19068
rect 10489 19012 10545 19068
rect 10545 19012 10549 19068
rect 10485 19008 10549 19012
rect 10565 19068 10629 19072
rect 10565 19012 10569 19068
rect 10569 19012 10625 19068
rect 10625 19012 10629 19068
rect 10565 19008 10629 19012
rect 10645 19068 10709 19072
rect 10645 19012 10649 19068
rect 10649 19012 10705 19068
rect 10705 19012 10709 19068
rect 10645 19008 10709 19012
rect 16707 19068 16771 19072
rect 16707 19012 16711 19068
rect 16711 19012 16767 19068
rect 16767 19012 16771 19068
rect 16707 19008 16771 19012
rect 16787 19068 16851 19072
rect 16787 19012 16791 19068
rect 16791 19012 16847 19068
rect 16847 19012 16851 19068
rect 16787 19008 16851 19012
rect 16867 19068 16931 19072
rect 16867 19012 16871 19068
rect 16871 19012 16927 19068
rect 16927 19012 16931 19068
rect 16867 19008 16931 19012
rect 16947 19068 17011 19072
rect 16947 19012 16951 19068
rect 16951 19012 17007 19068
rect 17007 19012 17011 19068
rect 16947 19008 17011 19012
rect 23009 19068 23073 19072
rect 23009 19012 23013 19068
rect 23013 19012 23069 19068
rect 23069 19012 23073 19068
rect 23009 19008 23073 19012
rect 23089 19068 23153 19072
rect 23089 19012 23093 19068
rect 23093 19012 23149 19068
rect 23149 19012 23153 19068
rect 23089 19008 23153 19012
rect 23169 19068 23233 19072
rect 23169 19012 23173 19068
rect 23173 19012 23229 19068
rect 23229 19012 23233 19068
rect 23169 19008 23233 19012
rect 23249 19068 23313 19072
rect 23249 19012 23253 19068
rect 23253 19012 23309 19068
rect 23309 19012 23313 19068
rect 23249 19008 23313 19012
rect 7254 18524 7318 18528
rect 7254 18468 7258 18524
rect 7258 18468 7314 18524
rect 7314 18468 7318 18524
rect 7254 18464 7318 18468
rect 7334 18524 7398 18528
rect 7334 18468 7338 18524
rect 7338 18468 7394 18524
rect 7394 18468 7398 18524
rect 7334 18464 7398 18468
rect 7414 18524 7478 18528
rect 7414 18468 7418 18524
rect 7418 18468 7474 18524
rect 7474 18468 7478 18524
rect 7414 18464 7478 18468
rect 7494 18524 7558 18528
rect 7494 18468 7498 18524
rect 7498 18468 7554 18524
rect 7554 18468 7558 18524
rect 7494 18464 7558 18468
rect 13556 18524 13620 18528
rect 13556 18468 13560 18524
rect 13560 18468 13616 18524
rect 13616 18468 13620 18524
rect 13556 18464 13620 18468
rect 13636 18524 13700 18528
rect 13636 18468 13640 18524
rect 13640 18468 13696 18524
rect 13696 18468 13700 18524
rect 13636 18464 13700 18468
rect 13716 18524 13780 18528
rect 13716 18468 13720 18524
rect 13720 18468 13776 18524
rect 13776 18468 13780 18524
rect 13716 18464 13780 18468
rect 13796 18524 13860 18528
rect 13796 18468 13800 18524
rect 13800 18468 13856 18524
rect 13856 18468 13860 18524
rect 13796 18464 13860 18468
rect 19858 18524 19922 18528
rect 19858 18468 19862 18524
rect 19862 18468 19918 18524
rect 19918 18468 19922 18524
rect 19858 18464 19922 18468
rect 19938 18524 20002 18528
rect 19938 18468 19942 18524
rect 19942 18468 19998 18524
rect 19998 18468 20002 18524
rect 19938 18464 20002 18468
rect 20018 18524 20082 18528
rect 20018 18468 20022 18524
rect 20022 18468 20078 18524
rect 20078 18468 20082 18524
rect 20018 18464 20082 18468
rect 20098 18524 20162 18528
rect 20098 18468 20102 18524
rect 20102 18468 20158 18524
rect 20158 18468 20162 18524
rect 20098 18464 20162 18468
rect 26160 18524 26224 18528
rect 26160 18468 26164 18524
rect 26164 18468 26220 18524
rect 26220 18468 26224 18524
rect 26160 18464 26224 18468
rect 26240 18524 26304 18528
rect 26240 18468 26244 18524
rect 26244 18468 26300 18524
rect 26300 18468 26304 18524
rect 26240 18464 26304 18468
rect 26320 18524 26384 18528
rect 26320 18468 26324 18524
rect 26324 18468 26380 18524
rect 26380 18468 26384 18524
rect 26320 18464 26384 18468
rect 26400 18524 26464 18528
rect 26400 18468 26404 18524
rect 26404 18468 26460 18524
rect 26460 18468 26464 18524
rect 26400 18464 26464 18468
rect 4103 17980 4167 17984
rect 4103 17924 4107 17980
rect 4107 17924 4163 17980
rect 4163 17924 4167 17980
rect 4103 17920 4167 17924
rect 4183 17980 4247 17984
rect 4183 17924 4187 17980
rect 4187 17924 4243 17980
rect 4243 17924 4247 17980
rect 4183 17920 4247 17924
rect 4263 17980 4327 17984
rect 4263 17924 4267 17980
rect 4267 17924 4323 17980
rect 4323 17924 4327 17980
rect 4263 17920 4327 17924
rect 4343 17980 4407 17984
rect 4343 17924 4347 17980
rect 4347 17924 4403 17980
rect 4403 17924 4407 17980
rect 4343 17920 4407 17924
rect 10405 17980 10469 17984
rect 10405 17924 10409 17980
rect 10409 17924 10465 17980
rect 10465 17924 10469 17980
rect 10405 17920 10469 17924
rect 10485 17980 10549 17984
rect 10485 17924 10489 17980
rect 10489 17924 10545 17980
rect 10545 17924 10549 17980
rect 10485 17920 10549 17924
rect 10565 17980 10629 17984
rect 10565 17924 10569 17980
rect 10569 17924 10625 17980
rect 10625 17924 10629 17980
rect 10565 17920 10629 17924
rect 10645 17980 10709 17984
rect 10645 17924 10649 17980
rect 10649 17924 10705 17980
rect 10705 17924 10709 17980
rect 10645 17920 10709 17924
rect 16707 17980 16771 17984
rect 16707 17924 16711 17980
rect 16711 17924 16767 17980
rect 16767 17924 16771 17980
rect 16707 17920 16771 17924
rect 16787 17980 16851 17984
rect 16787 17924 16791 17980
rect 16791 17924 16847 17980
rect 16847 17924 16851 17980
rect 16787 17920 16851 17924
rect 16867 17980 16931 17984
rect 16867 17924 16871 17980
rect 16871 17924 16927 17980
rect 16927 17924 16931 17980
rect 16867 17920 16931 17924
rect 16947 17980 17011 17984
rect 16947 17924 16951 17980
rect 16951 17924 17007 17980
rect 17007 17924 17011 17980
rect 16947 17920 17011 17924
rect 23009 17980 23073 17984
rect 23009 17924 23013 17980
rect 23013 17924 23069 17980
rect 23069 17924 23073 17980
rect 23009 17920 23073 17924
rect 23089 17980 23153 17984
rect 23089 17924 23093 17980
rect 23093 17924 23149 17980
rect 23149 17924 23153 17980
rect 23089 17920 23153 17924
rect 23169 17980 23233 17984
rect 23169 17924 23173 17980
rect 23173 17924 23229 17980
rect 23229 17924 23233 17980
rect 23169 17920 23233 17924
rect 23249 17980 23313 17984
rect 23249 17924 23253 17980
rect 23253 17924 23309 17980
rect 23309 17924 23313 17980
rect 23249 17920 23313 17924
rect 7254 17436 7318 17440
rect 7254 17380 7258 17436
rect 7258 17380 7314 17436
rect 7314 17380 7318 17436
rect 7254 17376 7318 17380
rect 7334 17436 7398 17440
rect 7334 17380 7338 17436
rect 7338 17380 7394 17436
rect 7394 17380 7398 17436
rect 7334 17376 7398 17380
rect 7414 17436 7478 17440
rect 7414 17380 7418 17436
rect 7418 17380 7474 17436
rect 7474 17380 7478 17436
rect 7414 17376 7478 17380
rect 7494 17436 7558 17440
rect 7494 17380 7498 17436
rect 7498 17380 7554 17436
rect 7554 17380 7558 17436
rect 7494 17376 7558 17380
rect 13556 17436 13620 17440
rect 13556 17380 13560 17436
rect 13560 17380 13616 17436
rect 13616 17380 13620 17436
rect 13556 17376 13620 17380
rect 13636 17436 13700 17440
rect 13636 17380 13640 17436
rect 13640 17380 13696 17436
rect 13696 17380 13700 17436
rect 13636 17376 13700 17380
rect 13716 17436 13780 17440
rect 13716 17380 13720 17436
rect 13720 17380 13776 17436
rect 13776 17380 13780 17436
rect 13716 17376 13780 17380
rect 13796 17436 13860 17440
rect 13796 17380 13800 17436
rect 13800 17380 13856 17436
rect 13856 17380 13860 17436
rect 13796 17376 13860 17380
rect 19858 17436 19922 17440
rect 19858 17380 19862 17436
rect 19862 17380 19918 17436
rect 19918 17380 19922 17436
rect 19858 17376 19922 17380
rect 19938 17436 20002 17440
rect 19938 17380 19942 17436
rect 19942 17380 19998 17436
rect 19998 17380 20002 17436
rect 19938 17376 20002 17380
rect 20018 17436 20082 17440
rect 20018 17380 20022 17436
rect 20022 17380 20078 17436
rect 20078 17380 20082 17436
rect 20018 17376 20082 17380
rect 20098 17436 20162 17440
rect 20098 17380 20102 17436
rect 20102 17380 20158 17436
rect 20158 17380 20162 17436
rect 20098 17376 20162 17380
rect 26160 17436 26224 17440
rect 26160 17380 26164 17436
rect 26164 17380 26220 17436
rect 26220 17380 26224 17436
rect 26160 17376 26224 17380
rect 26240 17436 26304 17440
rect 26240 17380 26244 17436
rect 26244 17380 26300 17436
rect 26300 17380 26304 17436
rect 26240 17376 26304 17380
rect 26320 17436 26384 17440
rect 26320 17380 26324 17436
rect 26324 17380 26380 17436
rect 26380 17380 26384 17436
rect 26320 17376 26384 17380
rect 26400 17436 26464 17440
rect 26400 17380 26404 17436
rect 26404 17380 26460 17436
rect 26460 17380 26464 17436
rect 26400 17376 26464 17380
rect 4103 16892 4167 16896
rect 4103 16836 4107 16892
rect 4107 16836 4163 16892
rect 4163 16836 4167 16892
rect 4103 16832 4167 16836
rect 4183 16892 4247 16896
rect 4183 16836 4187 16892
rect 4187 16836 4243 16892
rect 4243 16836 4247 16892
rect 4183 16832 4247 16836
rect 4263 16892 4327 16896
rect 4263 16836 4267 16892
rect 4267 16836 4323 16892
rect 4323 16836 4327 16892
rect 4263 16832 4327 16836
rect 4343 16892 4407 16896
rect 4343 16836 4347 16892
rect 4347 16836 4403 16892
rect 4403 16836 4407 16892
rect 4343 16832 4407 16836
rect 10405 16892 10469 16896
rect 10405 16836 10409 16892
rect 10409 16836 10465 16892
rect 10465 16836 10469 16892
rect 10405 16832 10469 16836
rect 10485 16892 10549 16896
rect 10485 16836 10489 16892
rect 10489 16836 10545 16892
rect 10545 16836 10549 16892
rect 10485 16832 10549 16836
rect 10565 16892 10629 16896
rect 10565 16836 10569 16892
rect 10569 16836 10625 16892
rect 10625 16836 10629 16892
rect 10565 16832 10629 16836
rect 10645 16892 10709 16896
rect 10645 16836 10649 16892
rect 10649 16836 10705 16892
rect 10705 16836 10709 16892
rect 10645 16832 10709 16836
rect 16707 16892 16771 16896
rect 16707 16836 16711 16892
rect 16711 16836 16767 16892
rect 16767 16836 16771 16892
rect 16707 16832 16771 16836
rect 16787 16892 16851 16896
rect 16787 16836 16791 16892
rect 16791 16836 16847 16892
rect 16847 16836 16851 16892
rect 16787 16832 16851 16836
rect 16867 16892 16931 16896
rect 16867 16836 16871 16892
rect 16871 16836 16927 16892
rect 16927 16836 16931 16892
rect 16867 16832 16931 16836
rect 16947 16892 17011 16896
rect 16947 16836 16951 16892
rect 16951 16836 17007 16892
rect 17007 16836 17011 16892
rect 16947 16832 17011 16836
rect 23009 16892 23073 16896
rect 23009 16836 23013 16892
rect 23013 16836 23069 16892
rect 23069 16836 23073 16892
rect 23009 16832 23073 16836
rect 23089 16892 23153 16896
rect 23089 16836 23093 16892
rect 23093 16836 23149 16892
rect 23149 16836 23153 16892
rect 23089 16832 23153 16836
rect 23169 16892 23233 16896
rect 23169 16836 23173 16892
rect 23173 16836 23229 16892
rect 23229 16836 23233 16892
rect 23169 16832 23233 16836
rect 23249 16892 23313 16896
rect 23249 16836 23253 16892
rect 23253 16836 23309 16892
rect 23309 16836 23313 16892
rect 23249 16832 23313 16836
rect 7254 16348 7318 16352
rect 7254 16292 7258 16348
rect 7258 16292 7314 16348
rect 7314 16292 7318 16348
rect 7254 16288 7318 16292
rect 7334 16348 7398 16352
rect 7334 16292 7338 16348
rect 7338 16292 7394 16348
rect 7394 16292 7398 16348
rect 7334 16288 7398 16292
rect 7414 16348 7478 16352
rect 7414 16292 7418 16348
rect 7418 16292 7474 16348
rect 7474 16292 7478 16348
rect 7414 16288 7478 16292
rect 7494 16348 7558 16352
rect 7494 16292 7498 16348
rect 7498 16292 7554 16348
rect 7554 16292 7558 16348
rect 7494 16288 7558 16292
rect 13556 16348 13620 16352
rect 13556 16292 13560 16348
rect 13560 16292 13616 16348
rect 13616 16292 13620 16348
rect 13556 16288 13620 16292
rect 13636 16348 13700 16352
rect 13636 16292 13640 16348
rect 13640 16292 13696 16348
rect 13696 16292 13700 16348
rect 13636 16288 13700 16292
rect 13716 16348 13780 16352
rect 13716 16292 13720 16348
rect 13720 16292 13776 16348
rect 13776 16292 13780 16348
rect 13716 16288 13780 16292
rect 13796 16348 13860 16352
rect 13796 16292 13800 16348
rect 13800 16292 13856 16348
rect 13856 16292 13860 16348
rect 13796 16288 13860 16292
rect 19858 16348 19922 16352
rect 19858 16292 19862 16348
rect 19862 16292 19918 16348
rect 19918 16292 19922 16348
rect 19858 16288 19922 16292
rect 19938 16348 20002 16352
rect 19938 16292 19942 16348
rect 19942 16292 19998 16348
rect 19998 16292 20002 16348
rect 19938 16288 20002 16292
rect 20018 16348 20082 16352
rect 20018 16292 20022 16348
rect 20022 16292 20078 16348
rect 20078 16292 20082 16348
rect 20018 16288 20082 16292
rect 20098 16348 20162 16352
rect 20098 16292 20102 16348
rect 20102 16292 20158 16348
rect 20158 16292 20162 16348
rect 20098 16288 20162 16292
rect 26160 16348 26224 16352
rect 26160 16292 26164 16348
rect 26164 16292 26220 16348
rect 26220 16292 26224 16348
rect 26160 16288 26224 16292
rect 26240 16348 26304 16352
rect 26240 16292 26244 16348
rect 26244 16292 26300 16348
rect 26300 16292 26304 16348
rect 26240 16288 26304 16292
rect 26320 16348 26384 16352
rect 26320 16292 26324 16348
rect 26324 16292 26380 16348
rect 26380 16292 26384 16348
rect 26320 16288 26384 16292
rect 26400 16348 26464 16352
rect 26400 16292 26404 16348
rect 26404 16292 26460 16348
rect 26460 16292 26464 16348
rect 26400 16288 26464 16292
rect 4103 15804 4167 15808
rect 4103 15748 4107 15804
rect 4107 15748 4163 15804
rect 4163 15748 4167 15804
rect 4103 15744 4167 15748
rect 4183 15804 4247 15808
rect 4183 15748 4187 15804
rect 4187 15748 4243 15804
rect 4243 15748 4247 15804
rect 4183 15744 4247 15748
rect 4263 15804 4327 15808
rect 4263 15748 4267 15804
rect 4267 15748 4323 15804
rect 4323 15748 4327 15804
rect 4263 15744 4327 15748
rect 4343 15804 4407 15808
rect 4343 15748 4347 15804
rect 4347 15748 4403 15804
rect 4403 15748 4407 15804
rect 4343 15744 4407 15748
rect 10405 15804 10469 15808
rect 10405 15748 10409 15804
rect 10409 15748 10465 15804
rect 10465 15748 10469 15804
rect 10405 15744 10469 15748
rect 10485 15804 10549 15808
rect 10485 15748 10489 15804
rect 10489 15748 10545 15804
rect 10545 15748 10549 15804
rect 10485 15744 10549 15748
rect 10565 15804 10629 15808
rect 10565 15748 10569 15804
rect 10569 15748 10625 15804
rect 10625 15748 10629 15804
rect 10565 15744 10629 15748
rect 10645 15804 10709 15808
rect 10645 15748 10649 15804
rect 10649 15748 10705 15804
rect 10705 15748 10709 15804
rect 10645 15744 10709 15748
rect 16707 15804 16771 15808
rect 16707 15748 16711 15804
rect 16711 15748 16767 15804
rect 16767 15748 16771 15804
rect 16707 15744 16771 15748
rect 16787 15804 16851 15808
rect 16787 15748 16791 15804
rect 16791 15748 16847 15804
rect 16847 15748 16851 15804
rect 16787 15744 16851 15748
rect 16867 15804 16931 15808
rect 16867 15748 16871 15804
rect 16871 15748 16927 15804
rect 16927 15748 16931 15804
rect 16867 15744 16931 15748
rect 16947 15804 17011 15808
rect 16947 15748 16951 15804
rect 16951 15748 17007 15804
rect 17007 15748 17011 15804
rect 16947 15744 17011 15748
rect 23009 15804 23073 15808
rect 23009 15748 23013 15804
rect 23013 15748 23069 15804
rect 23069 15748 23073 15804
rect 23009 15744 23073 15748
rect 23089 15804 23153 15808
rect 23089 15748 23093 15804
rect 23093 15748 23149 15804
rect 23149 15748 23153 15804
rect 23089 15744 23153 15748
rect 23169 15804 23233 15808
rect 23169 15748 23173 15804
rect 23173 15748 23229 15804
rect 23229 15748 23233 15804
rect 23169 15744 23233 15748
rect 23249 15804 23313 15808
rect 23249 15748 23253 15804
rect 23253 15748 23309 15804
rect 23309 15748 23313 15804
rect 23249 15744 23313 15748
rect 7254 15260 7318 15264
rect 7254 15204 7258 15260
rect 7258 15204 7314 15260
rect 7314 15204 7318 15260
rect 7254 15200 7318 15204
rect 7334 15260 7398 15264
rect 7334 15204 7338 15260
rect 7338 15204 7394 15260
rect 7394 15204 7398 15260
rect 7334 15200 7398 15204
rect 7414 15260 7478 15264
rect 7414 15204 7418 15260
rect 7418 15204 7474 15260
rect 7474 15204 7478 15260
rect 7414 15200 7478 15204
rect 7494 15260 7558 15264
rect 7494 15204 7498 15260
rect 7498 15204 7554 15260
rect 7554 15204 7558 15260
rect 7494 15200 7558 15204
rect 13556 15260 13620 15264
rect 13556 15204 13560 15260
rect 13560 15204 13616 15260
rect 13616 15204 13620 15260
rect 13556 15200 13620 15204
rect 13636 15260 13700 15264
rect 13636 15204 13640 15260
rect 13640 15204 13696 15260
rect 13696 15204 13700 15260
rect 13636 15200 13700 15204
rect 13716 15260 13780 15264
rect 13716 15204 13720 15260
rect 13720 15204 13776 15260
rect 13776 15204 13780 15260
rect 13716 15200 13780 15204
rect 13796 15260 13860 15264
rect 13796 15204 13800 15260
rect 13800 15204 13856 15260
rect 13856 15204 13860 15260
rect 13796 15200 13860 15204
rect 19858 15260 19922 15264
rect 19858 15204 19862 15260
rect 19862 15204 19918 15260
rect 19918 15204 19922 15260
rect 19858 15200 19922 15204
rect 19938 15260 20002 15264
rect 19938 15204 19942 15260
rect 19942 15204 19998 15260
rect 19998 15204 20002 15260
rect 19938 15200 20002 15204
rect 20018 15260 20082 15264
rect 20018 15204 20022 15260
rect 20022 15204 20078 15260
rect 20078 15204 20082 15260
rect 20018 15200 20082 15204
rect 20098 15260 20162 15264
rect 20098 15204 20102 15260
rect 20102 15204 20158 15260
rect 20158 15204 20162 15260
rect 20098 15200 20162 15204
rect 26160 15260 26224 15264
rect 26160 15204 26164 15260
rect 26164 15204 26220 15260
rect 26220 15204 26224 15260
rect 26160 15200 26224 15204
rect 26240 15260 26304 15264
rect 26240 15204 26244 15260
rect 26244 15204 26300 15260
rect 26300 15204 26304 15260
rect 26240 15200 26304 15204
rect 26320 15260 26384 15264
rect 26320 15204 26324 15260
rect 26324 15204 26380 15260
rect 26380 15204 26384 15260
rect 26320 15200 26384 15204
rect 26400 15260 26464 15264
rect 26400 15204 26404 15260
rect 26404 15204 26460 15260
rect 26460 15204 26464 15260
rect 26400 15200 26464 15204
rect 6500 14860 6564 14924
rect 4103 14716 4167 14720
rect 4103 14660 4107 14716
rect 4107 14660 4163 14716
rect 4163 14660 4167 14716
rect 4103 14656 4167 14660
rect 4183 14716 4247 14720
rect 4183 14660 4187 14716
rect 4187 14660 4243 14716
rect 4243 14660 4247 14716
rect 4183 14656 4247 14660
rect 4263 14716 4327 14720
rect 4263 14660 4267 14716
rect 4267 14660 4323 14716
rect 4323 14660 4327 14716
rect 4263 14656 4327 14660
rect 4343 14716 4407 14720
rect 4343 14660 4347 14716
rect 4347 14660 4403 14716
rect 4403 14660 4407 14716
rect 4343 14656 4407 14660
rect 10405 14716 10469 14720
rect 10405 14660 10409 14716
rect 10409 14660 10465 14716
rect 10465 14660 10469 14716
rect 10405 14656 10469 14660
rect 10485 14716 10549 14720
rect 10485 14660 10489 14716
rect 10489 14660 10545 14716
rect 10545 14660 10549 14716
rect 10485 14656 10549 14660
rect 10565 14716 10629 14720
rect 10565 14660 10569 14716
rect 10569 14660 10625 14716
rect 10625 14660 10629 14716
rect 10565 14656 10629 14660
rect 10645 14716 10709 14720
rect 10645 14660 10649 14716
rect 10649 14660 10705 14716
rect 10705 14660 10709 14716
rect 10645 14656 10709 14660
rect 16707 14716 16771 14720
rect 16707 14660 16711 14716
rect 16711 14660 16767 14716
rect 16767 14660 16771 14716
rect 16707 14656 16771 14660
rect 16787 14716 16851 14720
rect 16787 14660 16791 14716
rect 16791 14660 16847 14716
rect 16847 14660 16851 14716
rect 16787 14656 16851 14660
rect 16867 14716 16931 14720
rect 16867 14660 16871 14716
rect 16871 14660 16927 14716
rect 16927 14660 16931 14716
rect 16867 14656 16931 14660
rect 16947 14716 17011 14720
rect 16947 14660 16951 14716
rect 16951 14660 17007 14716
rect 17007 14660 17011 14716
rect 16947 14656 17011 14660
rect 23009 14716 23073 14720
rect 23009 14660 23013 14716
rect 23013 14660 23069 14716
rect 23069 14660 23073 14716
rect 23009 14656 23073 14660
rect 23089 14716 23153 14720
rect 23089 14660 23093 14716
rect 23093 14660 23149 14716
rect 23149 14660 23153 14716
rect 23089 14656 23153 14660
rect 23169 14716 23233 14720
rect 23169 14660 23173 14716
rect 23173 14660 23229 14716
rect 23229 14660 23233 14716
rect 23169 14656 23233 14660
rect 23249 14716 23313 14720
rect 23249 14660 23253 14716
rect 23253 14660 23309 14716
rect 23309 14660 23313 14716
rect 23249 14656 23313 14660
rect 7254 14172 7318 14176
rect 7254 14116 7258 14172
rect 7258 14116 7314 14172
rect 7314 14116 7318 14172
rect 7254 14112 7318 14116
rect 7334 14172 7398 14176
rect 7334 14116 7338 14172
rect 7338 14116 7394 14172
rect 7394 14116 7398 14172
rect 7334 14112 7398 14116
rect 7414 14172 7478 14176
rect 7414 14116 7418 14172
rect 7418 14116 7474 14172
rect 7474 14116 7478 14172
rect 7414 14112 7478 14116
rect 7494 14172 7558 14176
rect 7494 14116 7498 14172
rect 7498 14116 7554 14172
rect 7554 14116 7558 14172
rect 7494 14112 7558 14116
rect 13556 14172 13620 14176
rect 13556 14116 13560 14172
rect 13560 14116 13616 14172
rect 13616 14116 13620 14172
rect 13556 14112 13620 14116
rect 13636 14172 13700 14176
rect 13636 14116 13640 14172
rect 13640 14116 13696 14172
rect 13696 14116 13700 14172
rect 13636 14112 13700 14116
rect 13716 14172 13780 14176
rect 13716 14116 13720 14172
rect 13720 14116 13776 14172
rect 13776 14116 13780 14172
rect 13716 14112 13780 14116
rect 13796 14172 13860 14176
rect 13796 14116 13800 14172
rect 13800 14116 13856 14172
rect 13856 14116 13860 14172
rect 13796 14112 13860 14116
rect 19858 14172 19922 14176
rect 19858 14116 19862 14172
rect 19862 14116 19918 14172
rect 19918 14116 19922 14172
rect 19858 14112 19922 14116
rect 19938 14172 20002 14176
rect 19938 14116 19942 14172
rect 19942 14116 19998 14172
rect 19998 14116 20002 14172
rect 19938 14112 20002 14116
rect 20018 14172 20082 14176
rect 20018 14116 20022 14172
rect 20022 14116 20078 14172
rect 20078 14116 20082 14172
rect 20018 14112 20082 14116
rect 20098 14172 20162 14176
rect 20098 14116 20102 14172
rect 20102 14116 20158 14172
rect 20158 14116 20162 14172
rect 20098 14112 20162 14116
rect 26160 14172 26224 14176
rect 26160 14116 26164 14172
rect 26164 14116 26220 14172
rect 26220 14116 26224 14172
rect 26160 14112 26224 14116
rect 26240 14172 26304 14176
rect 26240 14116 26244 14172
rect 26244 14116 26300 14172
rect 26300 14116 26304 14172
rect 26240 14112 26304 14116
rect 26320 14172 26384 14176
rect 26320 14116 26324 14172
rect 26324 14116 26380 14172
rect 26380 14116 26384 14172
rect 26320 14112 26384 14116
rect 26400 14172 26464 14176
rect 26400 14116 26404 14172
rect 26404 14116 26460 14172
rect 26460 14116 26464 14172
rect 26400 14112 26464 14116
rect 4103 13628 4167 13632
rect 4103 13572 4107 13628
rect 4107 13572 4163 13628
rect 4163 13572 4167 13628
rect 4103 13568 4167 13572
rect 4183 13628 4247 13632
rect 4183 13572 4187 13628
rect 4187 13572 4243 13628
rect 4243 13572 4247 13628
rect 4183 13568 4247 13572
rect 4263 13628 4327 13632
rect 4263 13572 4267 13628
rect 4267 13572 4323 13628
rect 4323 13572 4327 13628
rect 4263 13568 4327 13572
rect 4343 13628 4407 13632
rect 4343 13572 4347 13628
rect 4347 13572 4403 13628
rect 4403 13572 4407 13628
rect 4343 13568 4407 13572
rect 10405 13628 10469 13632
rect 10405 13572 10409 13628
rect 10409 13572 10465 13628
rect 10465 13572 10469 13628
rect 10405 13568 10469 13572
rect 10485 13628 10549 13632
rect 10485 13572 10489 13628
rect 10489 13572 10545 13628
rect 10545 13572 10549 13628
rect 10485 13568 10549 13572
rect 10565 13628 10629 13632
rect 10565 13572 10569 13628
rect 10569 13572 10625 13628
rect 10625 13572 10629 13628
rect 10565 13568 10629 13572
rect 10645 13628 10709 13632
rect 10645 13572 10649 13628
rect 10649 13572 10705 13628
rect 10705 13572 10709 13628
rect 10645 13568 10709 13572
rect 16707 13628 16771 13632
rect 16707 13572 16711 13628
rect 16711 13572 16767 13628
rect 16767 13572 16771 13628
rect 16707 13568 16771 13572
rect 16787 13628 16851 13632
rect 16787 13572 16791 13628
rect 16791 13572 16847 13628
rect 16847 13572 16851 13628
rect 16787 13568 16851 13572
rect 16867 13628 16931 13632
rect 16867 13572 16871 13628
rect 16871 13572 16927 13628
rect 16927 13572 16931 13628
rect 16867 13568 16931 13572
rect 16947 13628 17011 13632
rect 16947 13572 16951 13628
rect 16951 13572 17007 13628
rect 17007 13572 17011 13628
rect 16947 13568 17011 13572
rect 23009 13628 23073 13632
rect 23009 13572 23013 13628
rect 23013 13572 23069 13628
rect 23069 13572 23073 13628
rect 23009 13568 23073 13572
rect 23089 13628 23153 13632
rect 23089 13572 23093 13628
rect 23093 13572 23149 13628
rect 23149 13572 23153 13628
rect 23089 13568 23153 13572
rect 23169 13628 23233 13632
rect 23169 13572 23173 13628
rect 23173 13572 23229 13628
rect 23229 13572 23233 13628
rect 23169 13568 23233 13572
rect 23249 13628 23313 13632
rect 23249 13572 23253 13628
rect 23253 13572 23309 13628
rect 23309 13572 23313 13628
rect 23249 13568 23313 13572
rect 7254 13084 7318 13088
rect 7254 13028 7258 13084
rect 7258 13028 7314 13084
rect 7314 13028 7318 13084
rect 7254 13024 7318 13028
rect 7334 13084 7398 13088
rect 7334 13028 7338 13084
rect 7338 13028 7394 13084
rect 7394 13028 7398 13084
rect 7334 13024 7398 13028
rect 7414 13084 7478 13088
rect 7414 13028 7418 13084
rect 7418 13028 7474 13084
rect 7474 13028 7478 13084
rect 7414 13024 7478 13028
rect 7494 13084 7558 13088
rect 7494 13028 7498 13084
rect 7498 13028 7554 13084
rect 7554 13028 7558 13084
rect 7494 13024 7558 13028
rect 13556 13084 13620 13088
rect 13556 13028 13560 13084
rect 13560 13028 13616 13084
rect 13616 13028 13620 13084
rect 13556 13024 13620 13028
rect 13636 13084 13700 13088
rect 13636 13028 13640 13084
rect 13640 13028 13696 13084
rect 13696 13028 13700 13084
rect 13636 13024 13700 13028
rect 13716 13084 13780 13088
rect 13716 13028 13720 13084
rect 13720 13028 13776 13084
rect 13776 13028 13780 13084
rect 13716 13024 13780 13028
rect 13796 13084 13860 13088
rect 13796 13028 13800 13084
rect 13800 13028 13856 13084
rect 13856 13028 13860 13084
rect 13796 13024 13860 13028
rect 19858 13084 19922 13088
rect 19858 13028 19862 13084
rect 19862 13028 19918 13084
rect 19918 13028 19922 13084
rect 19858 13024 19922 13028
rect 19938 13084 20002 13088
rect 19938 13028 19942 13084
rect 19942 13028 19998 13084
rect 19998 13028 20002 13084
rect 19938 13024 20002 13028
rect 20018 13084 20082 13088
rect 20018 13028 20022 13084
rect 20022 13028 20078 13084
rect 20078 13028 20082 13084
rect 20018 13024 20082 13028
rect 20098 13084 20162 13088
rect 20098 13028 20102 13084
rect 20102 13028 20158 13084
rect 20158 13028 20162 13084
rect 20098 13024 20162 13028
rect 26160 13084 26224 13088
rect 26160 13028 26164 13084
rect 26164 13028 26220 13084
rect 26220 13028 26224 13084
rect 26160 13024 26224 13028
rect 26240 13084 26304 13088
rect 26240 13028 26244 13084
rect 26244 13028 26300 13084
rect 26300 13028 26304 13084
rect 26240 13024 26304 13028
rect 26320 13084 26384 13088
rect 26320 13028 26324 13084
rect 26324 13028 26380 13084
rect 26380 13028 26384 13084
rect 26320 13024 26384 13028
rect 26400 13084 26464 13088
rect 26400 13028 26404 13084
rect 26404 13028 26460 13084
rect 26460 13028 26464 13084
rect 26400 13024 26464 13028
rect 4103 12540 4167 12544
rect 4103 12484 4107 12540
rect 4107 12484 4163 12540
rect 4163 12484 4167 12540
rect 4103 12480 4167 12484
rect 4183 12540 4247 12544
rect 4183 12484 4187 12540
rect 4187 12484 4243 12540
rect 4243 12484 4247 12540
rect 4183 12480 4247 12484
rect 4263 12540 4327 12544
rect 4263 12484 4267 12540
rect 4267 12484 4323 12540
rect 4323 12484 4327 12540
rect 4263 12480 4327 12484
rect 4343 12540 4407 12544
rect 4343 12484 4347 12540
rect 4347 12484 4403 12540
rect 4403 12484 4407 12540
rect 4343 12480 4407 12484
rect 10405 12540 10469 12544
rect 10405 12484 10409 12540
rect 10409 12484 10465 12540
rect 10465 12484 10469 12540
rect 10405 12480 10469 12484
rect 10485 12540 10549 12544
rect 10485 12484 10489 12540
rect 10489 12484 10545 12540
rect 10545 12484 10549 12540
rect 10485 12480 10549 12484
rect 10565 12540 10629 12544
rect 10565 12484 10569 12540
rect 10569 12484 10625 12540
rect 10625 12484 10629 12540
rect 10565 12480 10629 12484
rect 10645 12540 10709 12544
rect 10645 12484 10649 12540
rect 10649 12484 10705 12540
rect 10705 12484 10709 12540
rect 10645 12480 10709 12484
rect 16707 12540 16771 12544
rect 16707 12484 16711 12540
rect 16711 12484 16767 12540
rect 16767 12484 16771 12540
rect 16707 12480 16771 12484
rect 16787 12540 16851 12544
rect 16787 12484 16791 12540
rect 16791 12484 16847 12540
rect 16847 12484 16851 12540
rect 16787 12480 16851 12484
rect 16867 12540 16931 12544
rect 16867 12484 16871 12540
rect 16871 12484 16927 12540
rect 16927 12484 16931 12540
rect 16867 12480 16931 12484
rect 16947 12540 17011 12544
rect 16947 12484 16951 12540
rect 16951 12484 17007 12540
rect 17007 12484 17011 12540
rect 16947 12480 17011 12484
rect 23009 12540 23073 12544
rect 23009 12484 23013 12540
rect 23013 12484 23069 12540
rect 23069 12484 23073 12540
rect 23009 12480 23073 12484
rect 23089 12540 23153 12544
rect 23089 12484 23093 12540
rect 23093 12484 23149 12540
rect 23149 12484 23153 12540
rect 23089 12480 23153 12484
rect 23169 12540 23233 12544
rect 23169 12484 23173 12540
rect 23173 12484 23229 12540
rect 23229 12484 23233 12540
rect 23169 12480 23233 12484
rect 23249 12540 23313 12544
rect 23249 12484 23253 12540
rect 23253 12484 23309 12540
rect 23309 12484 23313 12540
rect 23249 12480 23313 12484
rect 7254 11996 7318 12000
rect 7254 11940 7258 11996
rect 7258 11940 7314 11996
rect 7314 11940 7318 11996
rect 7254 11936 7318 11940
rect 7334 11996 7398 12000
rect 7334 11940 7338 11996
rect 7338 11940 7394 11996
rect 7394 11940 7398 11996
rect 7334 11936 7398 11940
rect 7414 11996 7478 12000
rect 7414 11940 7418 11996
rect 7418 11940 7474 11996
rect 7474 11940 7478 11996
rect 7414 11936 7478 11940
rect 7494 11996 7558 12000
rect 7494 11940 7498 11996
rect 7498 11940 7554 11996
rect 7554 11940 7558 11996
rect 7494 11936 7558 11940
rect 13556 11996 13620 12000
rect 13556 11940 13560 11996
rect 13560 11940 13616 11996
rect 13616 11940 13620 11996
rect 13556 11936 13620 11940
rect 13636 11996 13700 12000
rect 13636 11940 13640 11996
rect 13640 11940 13696 11996
rect 13696 11940 13700 11996
rect 13636 11936 13700 11940
rect 13716 11996 13780 12000
rect 13716 11940 13720 11996
rect 13720 11940 13776 11996
rect 13776 11940 13780 11996
rect 13716 11936 13780 11940
rect 13796 11996 13860 12000
rect 13796 11940 13800 11996
rect 13800 11940 13856 11996
rect 13856 11940 13860 11996
rect 13796 11936 13860 11940
rect 19858 11996 19922 12000
rect 19858 11940 19862 11996
rect 19862 11940 19918 11996
rect 19918 11940 19922 11996
rect 19858 11936 19922 11940
rect 19938 11996 20002 12000
rect 19938 11940 19942 11996
rect 19942 11940 19998 11996
rect 19998 11940 20002 11996
rect 19938 11936 20002 11940
rect 20018 11996 20082 12000
rect 20018 11940 20022 11996
rect 20022 11940 20078 11996
rect 20078 11940 20082 11996
rect 20018 11936 20082 11940
rect 20098 11996 20162 12000
rect 20098 11940 20102 11996
rect 20102 11940 20158 11996
rect 20158 11940 20162 11996
rect 20098 11936 20162 11940
rect 26160 11996 26224 12000
rect 26160 11940 26164 11996
rect 26164 11940 26220 11996
rect 26220 11940 26224 11996
rect 26160 11936 26224 11940
rect 26240 11996 26304 12000
rect 26240 11940 26244 11996
rect 26244 11940 26300 11996
rect 26300 11940 26304 11996
rect 26240 11936 26304 11940
rect 26320 11996 26384 12000
rect 26320 11940 26324 11996
rect 26324 11940 26380 11996
rect 26380 11940 26384 11996
rect 26320 11936 26384 11940
rect 26400 11996 26464 12000
rect 26400 11940 26404 11996
rect 26404 11940 26460 11996
rect 26460 11940 26464 11996
rect 26400 11936 26464 11940
rect 4103 11452 4167 11456
rect 4103 11396 4107 11452
rect 4107 11396 4163 11452
rect 4163 11396 4167 11452
rect 4103 11392 4167 11396
rect 4183 11452 4247 11456
rect 4183 11396 4187 11452
rect 4187 11396 4243 11452
rect 4243 11396 4247 11452
rect 4183 11392 4247 11396
rect 4263 11452 4327 11456
rect 4263 11396 4267 11452
rect 4267 11396 4323 11452
rect 4323 11396 4327 11452
rect 4263 11392 4327 11396
rect 4343 11452 4407 11456
rect 4343 11396 4347 11452
rect 4347 11396 4403 11452
rect 4403 11396 4407 11452
rect 4343 11392 4407 11396
rect 10405 11452 10469 11456
rect 10405 11396 10409 11452
rect 10409 11396 10465 11452
rect 10465 11396 10469 11452
rect 10405 11392 10469 11396
rect 10485 11452 10549 11456
rect 10485 11396 10489 11452
rect 10489 11396 10545 11452
rect 10545 11396 10549 11452
rect 10485 11392 10549 11396
rect 10565 11452 10629 11456
rect 10565 11396 10569 11452
rect 10569 11396 10625 11452
rect 10625 11396 10629 11452
rect 10565 11392 10629 11396
rect 10645 11452 10709 11456
rect 10645 11396 10649 11452
rect 10649 11396 10705 11452
rect 10705 11396 10709 11452
rect 10645 11392 10709 11396
rect 16707 11452 16771 11456
rect 16707 11396 16711 11452
rect 16711 11396 16767 11452
rect 16767 11396 16771 11452
rect 16707 11392 16771 11396
rect 16787 11452 16851 11456
rect 16787 11396 16791 11452
rect 16791 11396 16847 11452
rect 16847 11396 16851 11452
rect 16787 11392 16851 11396
rect 16867 11452 16931 11456
rect 16867 11396 16871 11452
rect 16871 11396 16927 11452
rect 16927 11396 16931 11452
rect 16867 11392 16931 11396
rect 16947 11452 17011 11456
rect 16947 11396 16951 11452
rect 16951 11396 17007 11452
rect 17007 11396 17011 11452
rect 16947 11392 17011 11396
rect 23009 11452 23073 11456
rect 23009 11396 23013 11452
rect 23013 11396 23069 11452
rect 23069 11396 23073 11452
rect 23009 11392 23073 11396
rect 23089 11452 23153 11456
rect 23089 11396 23093 11452
rect 23093 11396 23149 11452
rect 23149 11396 23153 11452
rect 23089 11392 23153 11396
rect 23169 11452 23233 11456
rect 23169 11396 23173 11452
rect 23173 11396 23229 11452
rect 23229 11396 23233 11452
rect 23169 11392 23233 11396
rect 23249 11452 23313 11456
rect 23249 11396 23253 11452
rect 23253 11396 23309 11452
rect 23309 11396 23313 11452
rect 23249 11392 23313 11396
rect 7254 10908 7318 10912
rect 7254 10852 7258 10908
rect 7258 10852 7314 10908
rect 7314 10852 7318 10908
rect 7254 10848 7318 10852
rect 7334 10908 7398 10912
rect 7334 10852 7338 10908
rect 7338 10852 7394 10908
rect 7394 10852 7398 10908
rect 7334 10848 7398 10852
rect 7414 10908 7478 10912
rect 7414 10852 7418 10908
rect 7418 10852 7474 10908
rect 7474 10852 7478 10908
rect 7414 10848 7478 10852
rect 7494 10908 7558 10912
rect 7494 10852 7498 10908
rect 7498 10852 7554 10908
rect 7554 10852 7558 10908
rect 7494 10848 7558 10852
rect 13556 10908 13620 10912
rect 13556 10852 13560 10908
rect 13560 10852 13616 10908
rect 13616 10852 13620 10908
rect 13556 10848 13620 10852
rect 13636 10908 13700 10912
rect 13636 10852 13640 10908
rect 13640 10852 13696 10908
rect 13696 10852 13700 10908
rect 13636 10848 13700 10852
rect 13716 10908 13780 10912
rect 13716 10852 13720 10908
rect 13720 10852 13776 10908
rect 13776 10852 13780 10908
rect 13716 10848 13780 10852
rect 13796 10908 13860 10912
rect 13796 10852 13800 10908
rect 13800 10852 13856 10908
rect 13856 10852 13860 10908
rect 13796 10848 13860 10852
rect 19858 10908 19922 10912
rect 19858 10852 19862 10908
rect 19862 10852 19918 10908
rect 19918 10852 19922 10908
rect 19858 10848 19922 10852
rect 19938 10908 20002 10912
rect 19938 10852 19942 10908
rect 19942 10852 19998 10908
rect 19998 10852 20002 10908
rect 19938 10848 20002 10852
rect 20018 10908 20082 10912
rect 20018 10852 20022 10908
rect 20022 10852 20078 10908
rect 20078 10852 20082 10908
rect 20018 10848 20082 10852
rect 20098 10908 20162 10912
rect 20098 10852 20102 10908
rect 20102 10852 20158 10908
rect 20158 10852 20162 10908
rect 20098 10848 20162 10852
rect 26160 10908 26224 10912
rect 26160 10852 26164 10908
rect 26164 10852 26220 10908
rect 26220 10852 26224 10908
rect 26160 10848 26224 10852
rect 26240 10908 26304 10912
rect 26240 10852 26244 10908
rect 26244 10852 26300 10908
rect 26300 10852 26304 10908
rect 26240 10848 26304 10852
rect 26320 10908 26384 10912
rect 26320 10852 26324 10908
rect 26324 10852 26380 10908
rect 26380 10852 26384 10908
rect 26320 10848 26384 10852
rect 26400 10908 26464 10912
rect 26400 10852 26404 10908
rect 26404 10852 26460 10908
rect 26460 10852 26464 10908
rect 26400 10848 26464 10852
rect 4103 10364 4167 10368
rect 4103 10308 4107 10364
rect 4107 10308 4163 10364
rect 4163 10308 4167 10364
rect 4103 10304 4167 10308
rect 4183 10364 4247 10368
rect 4183 10308 4187 10364
rect 4187 10308 4243 10364
rect 4243 10308 4247 10364
rect 4183 10304 4247 10308
rect 4263 10364 4327 10368
rect 4263 10308 4267 10364
rect 4267 10308 4323 10364
rect 4323 10308 4327 10364
rect 4263 10304 4327 10308
rect 4343 10364 4407 10368
rect 4343 10308 4347 10364
rect 4347 10308 4403 10364
rect 4403 10308 4407 10364
rect 4343 10304 4407 10308
rect 10405 10364 10469 10368
rect 10405 10308 10409 10364
rect 10409 10308 10465 10364
rect 10465 10308 10469 10364
rect 10405 10304 10469 10308
rect 10485 10364 10549 10368
rect 10485 10308 10489 10364
rect 10489 10308 10545 10364
rect 10545 10308 10549 10364
rect 10485 10304 10549 10308
rect 10565 10364 10629 10368
rect 10565 10308 10569 10364
rect 10569 10308 10625 10364
rect 10625 10308 10629 10364
rect 10565 10304 10629 10308
rect 10645 10364 10709 10368
rect 10645 10308 10649 10364
rect 10649 10308 10705 10364
rect 10705 10308 10709 10364
rect 10645 10304 10709 10308
rect 16707 10364 16771 10368
rect 16707 10308 16711 10364
rect 16711 10308 16767 10364
rect 16767 10308 16771 10364
rect 16707 10304 16771 10308
rect 16787 10364 16851 10368
rect 16787 10308 16791 10364
rect 16791 10308 16847 10364
rect 16847 10308 16851 10364
rect 16787 10304 16851 10308
rect 16867 10364 16931 10368
rect 16867 10308 16871 10364
rect 16871 10308 16927 10364
rect 16927 10308 16931 10364
rect 16867 10304 16931 10308
rect 16947 10364 17011 10368
rect 16947 10308 16951 10364
rect 16951 10308 17007 10364
rect 17007 10308 17011 10364
rect 16947 10304 17011 10308
rect 23009 10364 23073 10368
rect 23009 10308 23013 10364
rect 23013 10308 23069 10364
rect 23069 10308 23073 10364
rect 23009 10304 23073 10308
rect 23089 10364 23153 10368
rect 23089 10308 23093 10364
rect 23093 10308 23149 10364
rect 23149 10308 23153 10364
rect 23089 10304 23153 10308
rect 23169 10364 23233 10368
rect 23169 10308 23173 10364
rect 23173 10308 23229 10364
rect 23229 10308 23233 10364
rect 23169 10304 23233 10308
rect 23249 10364 23313 10368
rect 23249 10308 23253 10364
rect 23253 10308 23309 10364
rect 23309 10308 23313 10364
rect 23249 10304 23313 10308
rect 7254 9820 7318 9824
rect 7254 9764 7258 9820
rect 7258 9764 7314 9820
rect 7314 9764 7318 9820
rect 7254 9760 7318 9764
rect 7334 9820 7398 9824
rect 7334 9764 7338 9820
rect 7338 9764 7394 9820
rect 7394 9764 7398 9820
rect 7334 9760 7398 9764
rect 7414 9820 7478 9824
rect 7414 9764 7418 9820
rect 7418 9764 7474 9820
rect 7474 9764 7478 9820
rect 7414 9760 7478 9764
rect 7494 9820 7558 9824
rect 7494 9764 7498 9820
rect 7498 9764 7554 9820
rect 7554 9764 7558 9820
rect 7494 9760 7558 9764
rect 13556 9820 13620 9824
rect 13556 9764 13560 9820
rect 13560 9764 13616 9820
rect 13616 9764 13620 9820
rect 13556 9760 13620 9764
rect 13636 9820 13700 9824
rect 13636 9764 13640 9820
rect 13640 9764 13696 9820
rect 13696 9764 13700 9820
rect 13636 9760 13700 9764
rect 13716 9820 13780 9824
rect 13716 9764 13720 9820
rect 13720 9764 13776 9820
rect 13776 9764 13780 9820
rect 13716 9760 13780 9764
rect 13796 9820 13860 9824
rect 13796 9764 13800 9820
rect 13800 9764 13856 9820
rect 13856 9764 13860 9820
rect 13796 9760 13860 9764
rect 19858 9820 19922 9824
rect 19858 9764 19862 9820
rect 19862 9764 19918 9820
rect 19918 9764 19922 9820
rect 19858 9760 19922 9764
rect 19938 9820 20002 9824
rect 19938 9764 19942 9820
rect 19942 9764 19998 9820
rect 19998 9764 20002 9820
rect 19938 9760 20002 9764
rect 20018 9820 20082 9824
rect 20018 9764 20022 9820
rect 20022 9764 20078 9820
rect 20078 9764 20082 9820
rect 20018 9760 20082 9764
rect 20098 9820 20162 9824
rect 20098 9764 20102 9820
rect 20102 9764 20158 9820
rect 20158 9764 20162 9820
rect 20098 9760 20162 9764
rect 26160 9820 26224 9824
rect 26160 9764 26164 9820
rect 26164 9764 26220 9820
rect 26220 9764 26224 9820
rect 26160 9760 26224 9764
rect 26240 9820 26304 9824
rect 26240 9764 26244 9820
rect 26244 9764 26300 9820
rect 26300 9764 26304 9820
rect 26240 9760 26304 9764
rect 26320 9820 26384 9824
rect 26320 9764 26324 9820
rect 26324 9764 26380 9820
rect 26380 9764 26384 9820
rect 26320 9760 26384 9764
rect 26400 9820 26464 9824
rect 26400 9764 26404 9820
rect 26404 9764 26460 9820
rect 26460 9764 26464 9820
rect 26400 9760 26464 9764
rect 4103 9276 4167 9280
rect 4103 9220 4107 9276
rect 4107 9220 4163 9276
rect 4163 9220 4167 9276
rect 4103 9216 4167 9220
rect 4183 9276 4247 9280
rect 4183 9220 4187 9276
rect 4187 9220 4243 9276
rect 4243 9220 4247 9276
rect 4183 9216 4247 9220
rect 4263 9276 4327 9280
rect 4263 9220 4267 9276
rect 4267 9220 4323 9276
rect 4323 9220 4327 9276
rect 4263 9216 4327 9220
rect 4343 9276 4407 9280
rect 4343 9220 4347 9276
rect 4347 9220 4403 9276
rect 4403 9220 4407 9276
rect 4343 9216 4407 9220
rect 10405 9276 10469 9280
rect 10405 9220 10409 9276
rect 10409 9220 10465 9276
rect 10465 9220 10469 9276
rect 10405 9216 10469 9220
rect 10485 9276 10549 9280
rect 10485 9220 10489 9276
rect 10489 9220 10545 9276
rect 10545 9220 10549 9276
rect 10485 9216 10549 9220
rect 10565 9276 10629 9280
rect 10565 9220 10569 9276
rect 10569 9220 10625 9276
rect 10625 9220 10629 9276
rect 10565 9216 10629 9220
rect 10645 9276 10709 9280
rect 10645 9220 10649 9276
rect 10649 9220 10705 9276
rect 10705 9220 10709 9276
rect 10645 9216 10709 9220
rect 16707 9276 16771 9280
rect 16707 9220 16711 9276
rect 16711 9220 16767 9276
rect 16767 9220 16771 9276
rect 16707 9216 16771 9220
rect 16787 9276 16851 9280
rect 16787 9220 16791 9276
rect 16791 9220 16847 9276
rect 16847 9220 16851 9276
rect 16787 9216 16851 9220
rect 16867 9276 16931 9280
rect 16867 9220 16871 9276
rect 16871 9220 16927 9276
rect 16927 9220 16931 9276
rect 16867 9216 16931 9220
rect 16947 9276 17011 9280
rect 16947 9220 16951 9276
rect 16951 9220 17007 9276
rect 17007 9220 17011 9276
rect 16947 9216 17011 9220
rect 23009 9276 23073 9280
rect 23009 9220 23013 9276
rect 23013 9220 23069 9276
rect 23069 9220 23073 9276
rect 23009 9216 23073 9220
rect 23089 9276 23153 9280
rect 23089 9220 23093 9276
rect 23093 9220 23149 9276
rect 23149 9220 23153 9276
rect 23089 9216 23153 9220
rect 23169 9276 23233 9280
rect 23169 9220 23173 9276
rect 23173 9220 23229 9276
rect 23229 9220 23233 9276
rect 23169 9216 23233 9220
rect 23249 9276 23313 9280
rect 23249 9220 23253 9276
rect 23253 9220 23309 9276
rect 23309 9220 23313 9276
rect 23249 9216 23313 9220
rect 7254 8732 7318 8736
rect 7254 8676 7258 8732
rect 7258 8676 7314 8732
rect 7314 8676 7318 8732
rect 7254 8672 7318 8676
rect 7334 8732 7398 8736
rect 7334 8676 7338 8732
rect 7338 8676 7394 8732
rect 7394 8676 7398 8732
rect 7334 8672 7398 8676
rect 7414 8732 7478 8736
rect 7414 8676 7418 8732
rect 7418 8676 7474 8732
rect 7474 8676 7478 8732
rect 7414 8672 7478 8676
rect 7494 8732 7558 8736
rect 7494 8676 7498 8732
rect 7498 8676 7554 8732
rect 7554 8676 7558 8732
rect 7494 8672 7558 8676
rect 13556 8732 13620 8736
rect 13556 8676 13560 8732
rect 13560 8676 13616 8732
rect 13616 8676 13620 8732
rect 13556 8672 13620 8676
rect 13636 8732 13700 8736
rect 13636 8676 13640 8732
rect 13640 8676 13696 8732
rect 13696 8676 13700 8732
rect 13636 8672 13700 8676
rect 13716 8732 13780 8736
rect 13716 8676 13720 8732
rect 13720 8676 13776 8732
rect 13776 8676 13780 8732
rect 13716 8672 13780 8676
rect 13796 8732 13860 8736
rect 13796 8676 13800 8732
rect 13800 8676 13856 8732
rect 13856 8676 13860 8732
rect 13796 8672 13860 8676
rect 19858 8732 19922 8736
rect 19858 8676 19862 8732
rect 19862 8676 19918 8732
rect 19918 8676 19922 8732
rect 19858 8672 19922 8676
rect 19938 8732 20002 8736
rect 19938 8676 19942 8732
rect 19942 8676 19998 8732
rect 19998 8676 20002 8732
rect 19938 8672 20002 8676
rect 20018 8732 20082 8736
rect 20018 8676 20022 8732
rect 20022 8676 20078 8732
rect 20078 8676 20082 8732
rect 20018 8672 20082 8676
rect 20098 8732 20162 8736
rect 20098 8676 20102 8732
rect 20102 8676 20158 8732
rect 20158 8676 20162 8732
rect 20098 8672 20162 8676
rect 26160 8732 26224 8736
rect 26160 8676 26164 8732
rect 26164 8676 26220 8732
rect 26220 8676 26224 8732
rect 26160 8672 26224 8676
rect 26240 8732 26304 8736
rect 26240 8676 26244 8732
rect 26244 8676 26300 8732
rect 26300 8676 26304 8732
rect 26240 8672 26304 8676
rect 26320 8732 26384 8736
rect 26320 8676 26324 8732
rect 26324 8676 26380 8732
rect 26380 8676 26384 8732
rect 26320 8672 26384 8676
rect 26400 8732 26464 8736
rect 26400 8676 26404 8732
rect 26404 8676 26460 8732
rect 26460 8676 26464 8732
rect 26400 8672 26464 8676
rect 4103 8188 4167 8192
rect 4103 8132 4107 8188
rect 4107 8132 4163 8188
rect 4163 8132 4167 8188
rect 4103 8128 4167 8132
rect 4183 8188 4247 8192
rect 4183 8132 4187 8188
rect 4187 8132 4243 8188
rect 4243 8132 4247 8188
rect 4183 8128 4247 8132
rect 4263 8188 4327 8192
rect 4263 8132 4267 8188
rect 4267 8132 4323 8188
rect 4323 8132 4327 8188
rect 4263 8128 4327 8132
rect 4343 8188 4407 8192
rect 4343 8132 4347 8188
rect 4347 8132 4403 8188
rect 4403 8132 4407 8188
rect 4343 8128 4407 8132
rect 10405 8188 10469 8192
rect 10405 8132 10409 8188
rect 10409 8132 10465 8188
rect 10465 8132 10469 8188
rect 10405 8128 10469 8132
rect 10485 8188 10549 8192
rect 10485 8132 10489 8188
rect 10489 8132 10545 8188
rect 10545 8132 10549 8188
rect 10485 8128 10549 8132
rect 10565 8188 10629 8192
rect 10565 8132 10569 8188
rect 10569 8132 10625 8188
rect 10625 8132 10629 8188
rect 10565 8128 10629 8132
rect 10645 8188 10709 8192
rect 10645 8132 10649 8188
rect 10649 8132 10705 8188
rect 10705 8132 10709 8188
rect 10645 8128 10709 8132
rect 16707 8188 16771 8192
rect 16707 8132 16711 8188
rect 16711 8132 16767 8188
rect 16767 8132 16771 8188
rect 16707 8128 16771 8132
rect 16787 8188 16851 8192
rect 16787 8132 16791 8188
rect 16791 8132 16847 8188
rect 16847 8132 16851 8188
rect 16787 8128 16851 8132
rect 16867 8188 16931 8192
rect 16867 8132 16871 8188
rect 16871 8132 16927 8188
rect 16927 8132 16931 8188
rect 16867 8128 16931 8132
rect 16947 8188 17011 8192
rect 16947 8132 16951 8188
rect 16951 8132 17007 8188
rect 17007 8132 17011 8188
rect 16947 8128 17011 8132
rect 23009 8188 23073 8192
rect 23009 8132 23013 8188
rect 23013 8132 23069 8188
rect 23069 8132 23073 8188
rect 23009 8128 23073 8132
rect 23089 8188 23153 8192
rect 23089 8132 23093 8188
rect 23093 8132 23149 8188
rect 23149 8132 23153 8188
rect 23089 8128 23153 8132
rect 23169 8188 23233 8192
rect 23169 8132 23173 8188
rect 23173 8132 23229 8188
rect 23229 8132 23233 8188
rect 23169 8128 23233 8132
rect 23249 8188 23313 8192
rect 23249 8132 23253 8188
rect 23253 8132 23309 8188
rect 23309 8132 23313 8188
rect 23249 8128 23313 8132
rect 7254 7644 7318 7648
rect 7254 7588 7258 7644
rect 7258 7588 7314 7644
rect 7314 7588 7318 7644
rect 7254 7584 7318 7588
rect 7334 7644 7398 7648
rect 7334 7588 7338 7644
rect 7338 7588 7394 7644
rect 7394 7588 7398 7644
rect 7334 7584 7398 7588
rect 7414 7644 7478 7648
rect 7414 7588 7418 7644
rect 7418 7588 7474 7644
rect 7474 7588 7478 7644
rect 7414 7584 7478 7588
rect 7494 7644 7558 7648
rect 7494 7588 7498 7644
rect 7498 7588 7554 7644
rect 7554 7588 7558 7644
rect 7494 7584 7558 7588
rect 13556 7644 13620 7648
rect 13556 7588 13560 7644
rect 13560 7588 13616 7644
rect 13616 7588 13620 7644
rect 13556 7584 13620 7588
rect 13636 7644 13700 7648
rect 13636 7588 13640 7644
rect 13640 7588 13696 7644
rect 13696 7588 13700 7644
rect 13636 7584 13700 7588
rect 13716 7644 13780 7648
rect 13716 7588 13720 7644
rect 13720 7588 13776 7644
rect 13776 7588 13780 7644
rect 13716 7584 13780 7588
rect 13796 7644 13860 7648
rect 13796 7588 13800 7644
rect 13800 7588 13856 7644
rect 13856 7588 13860 7644
rect 13796 7584 13860 7588
rect 19858 7644 19922 7648
rect 19858 7588 19862 7644
rect 19862 7588 19918 7644
rect 19918 7588 19922 7644
rect 19858 7584 19922 7588
rect 19938 7644 20002 7648
rect 19938 7588 19942 7644
rect 19942 7588 19998 7644
rect 19998 7588 20002 7644
rect 19938 7584 20002 7588
rect 20018 7644 20082 7648
rect 20018 7588 20022 7644
rect 20022 7588 20078 7644
rect 20078 7588 20082 7644
rect 20018 7584 20082 7588
rect 20098 7644 20162 7648
rect 20098 7588 20102 7644
rect 20102 7588 20158 7644
rect 20158 7588 20162 7644
rect 20098 7584 20162 7588
rect 26160 7644 26224 7648
rect 26160 7588 26164 7644
rect 26164 7588 26220 7644
rect 26220 7588 26224 7644
rect 26160 7584 26224 7588
rect 26240 7644 26304 7648
rect 26240 7588 26244 7644
rect 26244 7588 26300 7644
rect 26300 7588 26304 7644
rect 26240 7584 26304 7588
rect 26320 7644 26384 7648
rect 26320 7588 26324 7644
rect 26324 7588 26380 7644
rect 26380 7588 26384 7644
rect 26320 7584 26384 7588
rect 26400 7644 26464 7648
rect 26400 7588 26404 7644
rect 26404 7588 26460 7644
rect 26460 7588 26464 7644
rect 26400 7584 26464 7588
rect 4103 7100 4167 7104
rect 4103 7044 4107 7100
rect 4107 7044 4163 7100
rect 4163 7044 4167 7100
rect 4103 7040 4167 7044
rect 4183 7100 4247 7104
rect 4183 7044 4187 7100
rect 4187 7044 4243 7100
rect 4243 7044 4247 7100
rect 4183 7040 4247 7044
rect 4263 7100 4327 7104
rect 4263 7044 4267 7100
rect 4267 7044 4323 7100
rect 4323 7044 4327 7100
rect 4263 7040 4327 7044
rect 4343 7100 4407 7104
rect 4343 7044 4347 7100
rect 4347 7044 4403 7100
rect 4403 7044 4407 7100
rect 4343 7040 4407 7044
rect 10405 7100 10469 7104
rect 10405 7044 10409 7100
rect 10409 7044 10465 7100
rect 10465 7044 10469 7100
rect 10405 7040 10469 7044
rect 10485 7100 10549 7104
rect 10485 7044 10489 7100
rect 10489 7044 10545 7100
rect 10545 7044 10549 7100
rect 10485 7040 10549 7044
rect 10565 7100 10629 7104
rect 10565 7044 10569 7100
rect 10569 7044 10625 7100
rect 10625 7044 10629 7100
rect 10565 7040 10629 7044
rect 10645 7100 10709 7104
rect 10645 7044 10649 7100
rect 10649 7044 10705 7100
rect 10705 7044 10709 7100
rect 10645 7040 10709 7044
rect 16707 7100 16771 7104
rect 16707 7044 16711 7100
rect 16711 7044 16767 7100
rect 16767 7044 16771 7100
rect 16707 7040 16771 7044
rect 16787 7100 16851 7104
rect 16787 7044 16791 7100
rect 16791 7044 16847 7100
rect 16847 7044 16851 7100
rect 16787 7040 16851 7044
rect 16867 7100 16931 7104
rect 16867 7044 16871 7100
rect 16871 7044 16927 7100
rect 16927 7044 16931 7100
rect 16867 7040 16931 7044
rect 16947 7100 17011 7104
rect 16947 7044 16951 7100
rect 16951 7044 17007 7100
rect 17007 7044 17011 7100
rect 16947 7040 17011 7044
rect 23009 7100 23073 7104
rect 23009 7044 23013 7100
rect 23013 7044 23069 7100
rect 23069 7044 23073 7100
rect 23009 7040 23073 7044
rect 23089 7100 23153 7104
rect 23089 7044 23093 7100
rect 23093 7044 23149 7100
rect 23149 7044 23153 7100
rect 23089 7040 23153 7044
rect 23169 7100 23233 7104
rect 23169 7044 23173 7100
rect 23173 7044 23229 7100
rect 23229 7044 23233 7100
rect 23169 7040 23233 7044
rect 23249 7100 23313 7104
rect 23249 7044 23253 7100
rect 23253 7044 23309 7100
rect 23309 7044 23313 7100
rect 23249 7040 23313 7044
rect 7254 6556 7318 6560
rect 7254 6500 7258 6556
rect 7258 6500 7314 6556
rect 7314 6500 7318 6556
rect 7254 6496 7318 6500
rect 7334 6556 7398 6560
rect 7334 6500 7338 6556
rect 7338 6500 7394 6556
rect 7394 6500 7398 6556
rect 7334 6496 7398 6500
rect 7414 6556 7478 6560
rect 7414 6500 7418 6556
rect 7418 6500 7474 6556
rect 7474 6500 7478 6556
rect 7414 6496 7478 6500
rect 7494 6556 7558 6560
rect 7494 6500 7498 6556
rect 7498 6500 7554 6556
rect 7554 6500 7558 6556
rect 7494 6496 7558 6500
rect 13556 6556 13620 6560
rect 13556 6500 13560 6556
rect 13560 6500 13616 6556
rect 13616 6500 13620 6556
rect 13556 6496 13620 6500
rect 13636 6556 13700 6560
rect 13636 6500 13640 6556
rect 13640 6500 13696 6556
rect 13696 6500 13700 6556
rect 13636 6496 13700 6500
rect 13716 6556 13780 6560
rect 13716 6500 13720 6556
rect 13720 6500 13776 6556
rect 13776 6500 13780 6556
rect 13716 6496 13780 6500
rect 13796 6556 13860 6560
rect 13796 6500 13800 6556
rect 13800 6500 13856 6556
rect 13856 6500 13860 6556
rect 13796 6496 13860 6500
rect 19858 6556 19922 6560
rect 19858 6500 19862 6556
rect 19862 6500 19918 6556
rect 19918 6500 19922 6556
rect 19858 6496 19922 6500
rect 19938 6556 20002 6560
rect 19938 6500 19942 6556
rect 19942 6500 19998 6556
rect 19998 6500 20002 6556
rect 19938 6496 20002 6500
rect 20018 6556 20082 6560
rect 20018 6500 20022 6556
rect 20022 6500 20078 6556
rect 20078 6500 20082 6556
rect 20018 6496 20082 6500
rect 20098 6556 20162 6560
rect 20098 6500 20102 6556
rect 20102 6500 20158 6556
rect 20158 6500 20162 6556
rect 20098 6496 20162 6500
rect 26160 6556 26224 6560
rect 26160 6500 26164 6556
rect 26164 6500 26220 6556
rect 26220 6500 26224 6556
rect 26160 6496 26224 6500
rect 26240 6556 26304 6560
rect 26240 6500 26244 6556
rect 26244 6500 26300 6556
rect 26300 6500 26304 6556
rect 26240 6496 26304 6500
rect 26320 6556 26384 6560
rect 26320 6500 26324 6556
rect 26324 6500 26380 6556
rect 26380 6500 26384 6556
rect 26320 6496 26384 6500
rect 26400 6556 26464 6560
rect 26400 6500 26404 6556
rect 26404 6500 26460 6556
rect 26460 6500 26464 6556
rect 26400 6496 26464 6500
rect 4103 6012 4167 6016
rect 4103 5956 4107 6012
rect 4107 5956 4163 6012
rect 4163 5956 4167 6012
rect 4103 5952 4167 5956
rect 4183 6012 4247 6016
rect 4183 5956 4187 6012
rect 4187 5956 4243 6012
rect 4243 5956 4247 6012
rect 4183 5952 4247 5956
rect 4263 6012 4327 6016
rect 4263 5956 4267 6012
rect 4267 5956 4323 6012
rect 4323 5956 4327 6012
rect 4263 5952 4327 5956
rect 4343 6012 4407 6016
rect 4343 5956 4347 6012
rect 4347 5956 4403 6012
rect 4403 5956 4407 6012
rect 4343 5952 4407 5956
rect 10405 6012 10469 6016
rect 10405 5956 10409 6012
rect 10409 5956 10465 6012
rect 10465 5956 10469 6012
rect 10405 5952 10469 5956
rect 10485 6012 10549 6016
rect 10485 5956 10489 6012
rect 10489 5956 10545 6012
rect 10545 5956 10549 6012
rect 10485 5952 10549 5956
rect 10565 6012 10629 6016
rect 10565 5956 10569 6012
rect 10569 5956 10625 6012
rect 10625 5956 10629 6012
rect 10565 5952 10629 5956
rect 10645 6012 10709 6016
rect 10645 5956 10649 6012
rect 10649 5956 10705 6012
rect 10705 5956 10709 6012
rect 10645 5952 10709 5956
rect 16707 6012 16771 6016
rect 16707 5956 16711 6012
rect 16711 5956 16767 6012
rect 16767 5956 16771 6012
rect 16707 5952 16771 5956
rect 16787 6012 16851 6016
rect 16787 5956 16791 6012
rect 16791 5956 16847 6012
rect 16847 5956 16851 6012
rect 16787 5952 16851 5956
rect 16867 6012 16931 6016
rect 16867 5956 16871 6012
rect 16871 5956 16927 6012
rect 16927 5956 16931 6012
rect 16867 5952 16931 5956
rect 16947 6012 17011 6016
rect 16947 5956 16951 6012
rect 16951 5956 17007 6012
rect 17007 5956 17011 6012
rect 16947 5952 17011 5956
rect 23009 6012 23073 6016
rect 23009 5956 23013 6012
rect 23013 5956 23069 6012
rect 23069 5956 23073 6012
rect 23009 5952 23073 5956
rect 23089 6012 23153 6016
rect 23089 5956 23093 6012
rect 23093 5956 23149 6012
rect 23149 5956 23153 6012
rect 23089 5952 23153 5956
rect 23169 6012 23233 6016
rect 23169 5956 23173 6012
rect 23173 5956 23229 6012
rect 23229 5956 23233 6012
rect 23169 5952 23233 5956
rect 23249 6012 23313 6016
rect 23249 5956 23253 6012
rect 23253 5956 23309 6012
rect 23309 5956 23313 6012
rect 23249 5952 23313 5956
rect 7254 5468 7318 5472
rect 7254 5412 7258 5468
rect 7258 5412 7314 5468
rect 7314 5412 7318 5468
rect 7254 5408 7318 5412
rect 7334 5468 7398 5472
rect 7334 5412 7338 5468
rect 7338 5412 7394 5468
rect 7394 5412 7398 5468
rect 7334 5408 7398 5412
rect 7414 5468 7478 5472
rect 7414 5412 7418 5468
rect 7418 5412 7474 5468
rect 7474 5412 7478 5468
rect 7414 5408 7478 5412
rect 7494 5468 7558 5472
rect 7494 5412 7498 5468
rect 7498 5412 7554 5468
rect 7554 5412 7558 5468
rect 7494 5408 7558 5412
rect 13556 5468 13620 5472
rect 13556 5412 13560 5468
rect 13560 5412 13616 5468
rect 13616 5412 13620 5468
rect 13556 5408 13620 5412
rect 13636 5468 13700 5472
rect 13636 5412 13640 5468
rect 13640 5412 13696 5468
rect 13696 5412 13700 5468
rect 13636 5408 13700 5412
rect 13716 5468 13780 5472
rect 13716 5412 13720 5468
rect 13720 5412 13776 5468
rect 13776 5412 13780 5468
rect 13716 5408 13780 5412
rect 13796 5468 13860 5472
rect 13796 5412 13800 5468
rect 13800 5412 13856 5468
rect 13856 5412 13860 5468
rect 13796 5408 13860 5412
rect 19858 5468 19922 5472
rect 19858 5412 19862 5468
rect 19862 5412 19918 5468
rect 19918 5412 19922 5468
rect 19858 5408 19922 5412
rect 19938 5468 20002 5472
rect 19938 5412 19942 5468
rect 19942 5412 19998 5468
rect 19998 5412 20002 5468
rect 19938 5408 20002 5412
rect 20018 5468 20082 5472
rect 20018 5412 20022 5468
rect 20022 5412 20078 5468
rect 20078 5412 20082 5468
rect 20018 5408 20082 5412
rect 20098 5468 20162 5472
rect 20098 5412 20102 5468
rect 20102 5412 20158 5468
rect 20158 5412 20162 5468
rect 20098 5408 20162 5412
rect 26160 5468 26224 5472
rect 26160 5412 26164 5468
rect 26164 5412 26220 5468
rect 26220 5412 26224 5468
rect 26160 5408 26224 5412
rect 26240 5468 26304 5472
rect 26240 5412 26244 5468
rect 26244 5412 26300 5468
rect 26300 5412 26304 5468
rect 26240 5408 26304 5412
rect 26320 5468 26384 5472
rect 26320 5412 26324 5468
rect 26324 5412 26380 5468
rect 26380 5412 26384 5468
rect 26320 5408 26384 5412
rect 26400 5468 26464 5472
rect 26400 5412 26404 5468
rect 26404 5412 26460 5468
rect 26460 5412 26464 5468
rect 26400 5408 26464 5412
rect 4103 4924 4167 4928
rect 4103 4868 4107 4924
rect 4107 4868 4163 4924
rect 4163 4868 4167 4924
rect 4103 4864 4167 4868
rect 4183 4924 4247 4928
rect 4183 4868 4187 4924
rect 4187 4868 4243 4924
rect 4243 4868 4247 4924
rect 4183 4864 4247 4868
rect 4263 4924 4327 4928
rect 4263 4868 4267 4924
rect 4267 4868 4323 4924
rect 4323 4868 4327 4924
rect 4263 4864 4327 4868
rect 4343 4924 4407 4928
rect 4343 4868 4347 4924
rect 4347 4868 4403 4924
rect 4403 4868 4407 4924
rect 4343 4864 4407 4868
rect 10405 4924 10469 4928
rect 10405 4868 10409 4924
rect 10409 4868 10465 4924
rect 10465 4868 10469 4924
rect 10405 4864 10469 4868
rect 10485 4924 10549 4928
rect 10485 4868 10489 4924
rect 10489 4868 10545 4924
rect 10545 4868 10549 4924
rect 10485 4864 10549 4868
rect 10565 4924 10629 4928
rect 10565 4868 10569 4924
rect 10569 4868 10625 4924
rect 10625 4868 10629 4924
rect 10565 4864 10629 4868
rect 10645 4924 10709 4928
rect 10645 4868 10649 4924
rect 10649 4868 10705 4924
rect 10705 4868 10709 4924
rect 10645 4864 10709 4868
rect 16707 4924 16771 4928
rect 16707 4868 16711 4924
rect 16711 4868 16767 4924
rect 16767 4868 16771 4924
rect 16707 4864 16771 4868
rect 16787 4924 16851 4928
rect 16787 4868 16791 4924
rect 16791 4868 16847 4924
rect 16847 4868 16851 4924
rect 16787 4864 16851 4868
rect 16867 4924 16931 4928
rect 16867 4868 16871 4924
rect 16871 4868 16927 4924
rect 16927 4868 16931 4924
rect 16867 4864 16931 4868
rect 16947 4924 17011 4928
rect 16947 4868 16951 4924
rect 16951 4868 17007 4924
rect 17007 4868 17011 4924
rect 16947 4864 17011 4868
rect 23009 4924 23073 4928
rect 23009 4868 23013 4924
rect 23013 4868 23069 4924
rect 23069 4868 23073 4924
rect 23009 4864 23073 4868
rect 23089 4924 23153 4928
rect 23089 4868 23093 4924
rect 23093 4868 23149 4924
rect 23149 4868 23153 4924
rect 23089 4864 23153 4868
rect 23169 4924 23233 4928
rect 23169 4868 23173 4924
rect 23173 4868 23229 4924
rect 23229 4868 23233 4924
rect 23169 4864 23233 4868
rect 23249 4924 23313 4928
rect 23249 4868 23253 4924
rect 23253 4868 23309 4924
rect 23309 4868 23313 4924
rect 23249 4864 23313 4868
rect 7254 4380 7318 4384
rect 7254 4324 7258 4380
rect 7258 4324 7314 4380
rect 7314 4324 7318 4380
rect 7254 4320 7318 4324
rect 7334 4380 7398 4384
rect 7334 4324 7338 4380
rect 7338 4324 7394 4380
rect 7394 4324 7398 4380
rect 7334 4320 7398 4324
rect 7414 4380 7478 4384
rect 7414 4324 7418 4380
rect 7418 4324 7474 4380
rect 7474 4324 7478 4380
rect 7414 4320 7478 4324
rect 7494 4380 7558 4384
rect 7494 4324 7498 4380
rect 7498 4324 7554 4380
rect 7554 4324 7558 4380
rect 7494 4320 7558 4324
rect 13556 4380 13620 4384
rect 13556 4324 13560 4380
rect 13560 4324 13616 4380
rect 13616 4324 13620 4380
rect 13556 4320 13620 4324
rect 13636 4380 13700 4384
rect 13636 4324 13640 4380
rect 13640 4324 13696 4380
rect 13696 4324 13700 4380
rect 13636 4320 13700 4324
rect 13716 4380 13780 4384
rect 13716 4324 13720 4380
rect 13720 4324 13776 4380
rect 13776 4324 13780 4380
rect 13716 4320 13780 4324
rect 13796 4380 13860 4384
rect 13796 4324 13800 4380
rect 13800 4324 13856 4380
rect 13856 4324 13860 4380
rect 13796 4320 13860 4324
rect 19858 4380 19922 4384
rect 19858 4324 19862 4380
rect 19862 4324 19918 4380
rect 19918 4324 19922 4380
rect 19858 4320 19922 4324
rect 19938 4380 20002 4384
rect 19938 4324 19942 4380
rect 19942 4324 19998 4380
rect 19998 4324 20002 4380
rect 19938 4320 20002 4324
rect 20018 4380 20082 4384
rect 20018 4324 20022 4380
rect 20022 4324 20078 4380
rect 20078 4324 20082 4380
rect 20018 4320 20082 4324
rect 20098 4380 20162 4384
rect 20098 4324 20102 4380
rect 20102 4324 20158 4380
rect 20158 4324 20162 4380
rect 20098 4320 20162 4324
rect 26160 4380 26224 4384
rect 26160 4324 26164 4380
rect 26164 4324 26220 4380
rect 26220 4324 26224 4380
rect 26160 4320 26224 4324
rect 26240 4380 26304 4384
rect 26240 4324 26244 4380
rect 26244 4324 26300 4380
rect 26300 4324 26304 4380
rect 26240 4320 26304 4324
rect 26320 4380 26384 4384
rect 26320 4324 26324 4380
rect 26324 4324 26380 4380
rect 26380 4324 26384 4380
rect 26320 4320 26384 4324
rect 26400 4380 26464 4384
rect 26400 4324 26404 4380
rect 26404 4324 26460 4380
rect 26460 4324 26464 4380
rect 26400 4320 26464 4324
rect 4103 3836 4167 3840
rect 4103 3780 4107 3836
rect 4107 3780 4163 3836
rect 4163 3780 4167 3836
rect 4103 3776 4167 3780
rect 4183 3836 4247 3840
rect 4183 3780 4187 3836
rect 4187 3780 4243 3836
rect 4243 3780 4247 3836
rect 4183 3776 4247 3780
rect 4263 3836 4327 3840
rect 4263 3780 4267 3836
rect 4267 3780 4323 3836
rect 4323 3780 4327 3836
rect 4263 3776 4327 3780
rect 4343 3836 4407 3840
rect 4343 3780 4347 3836
rect 4347 3780 4403 3836
rect 4403 3780 4407 3836
rect 4343 3776 4407 3780
rect 10405 3836 10469 3840
rect 10405 3780 10409 3836
rect 10409 3780 10465 3836
rect 10465 3780 10469 3836
rect 10405 3776 10469 3780
rect 10485 3836 10549 3840
rect 10485 3780 10489 3836
rect 10489 3780 10545 3836
rect 10545 3780 10549 3836
rect 10485 3776 10549 3780
rect 10565 3836 10629 3840
rect 10565 3780 10569 3836
rect 10569 3780 10625 3836
rect 10625 3780 10629 3836
rect 10565 3776 10629 3780
rect 10645 3836 10709 3840
rect 10645 3780 10649 3836
rect 10649 3780 10705 3836
rect 10705 3780 10709 3836
rect 10645 3776 10709 3780
rect 16707 3836 16771 3840
rect 16707 3780 16711 3836
rect 16711 3780 16767 3836
rect 16767 3780 16771 3836
rect 16707 3776 16771 3780
rect 16787 3836 16851 3840
rect 16787 3780 16791 3836
rect 16791 3780 16847 3836
rect 16847 3780 16851 3836
rect 16787 3776 16851 3780
rect 16867 3836 16931 3840
rect 16867 3780 16871 3836
rect 16871 3780 16927 3836
rect 16927 3780 16931 3836
rect 16867 3776 16931 3780
rect 16947 3836 17011 3840
rect 16947 3780 16951 3836
rect 16951 3780 17007 3836
rect 17007 3780 17011 3836
rect 16947 3776 17011 3780
rect 23009 3836 23073 3840
rect 23009 3780 23013 3836
rect 23013 3780 23069 3836
rect 23069 3780 23073 3836
rect 23009 3776 23073 3780
rect 23089 3836 23153 3840
rect 23089 3780 23093 3836
rect 23093 3780 23149 3836
rect 23149 3780 23153 3836
rect 23089 3776 23153 3780
rect 23169 3836 23233 3840
rect 23169 3780 23173 3836
rect 23173 3780 23229 3836
rect 23229 3780 23233 3836
rect 23169 3776 23233 3780
rect 23249 3836 23313 3840
rect 23249 3780 23253 3836
rect 23253 3780 23309 3836
rect 23309 3780 23313 3836
rect 23249 3776 23313 3780
rect 7254 3292 7318 3296
rect 7254 3236 7258 3292
rect 7258 3236 7314 3292
rect 7314 3236 7318 3292
rect 7254 3232 7318 3236
rect 7334 3292 7398 3296
rect 7334 3236 7338 3292
rect 7338 3236 7394 3292
rect 7394 3236 7398 3292
rect 7334 3232 7398 3236
rect 7414 3292 7478 3296
rect 7414 3236 7418 3292
rect 7418 3236 7474 3292
rect 7474 3236 7478 3292
rect 7414 3232 7478 3236
rect 7494 3292 7558 3296
rect 7494 3236 7498 3292
rect 7498 3236 7554 3292
rect 7554 3236 7558 3292
rect 7494 3232 7558 3236
rect 13556 3292 13620 3296
rect 13556 3236 13560 3292
rect 13560 3236 13616 3292
rect 13616 3236 13620 3292
rect 13556 3232 13620 3236
rect 13636 3292 13700 3296
rect 13636 3236 13640 3292
rect 13640 3236 13696 3292
rect 13696 3236 13700 3292
rect 13636 3232 13700 3236
rect 13716 3292 13780 3296
rect 13716 3236 13720 3292
rect 13720 3236 13776 3292
rect 13776 3236 13780 3292
rect 13716 3232 13780 3236
rect 13796 3292 13860 3296
rect 13796 3236 13800 3292
rect 13800 3236 13856 3292
rect 13856 3236 13860 3292
rect 13796 3232 13860 3236
rect 19858 3292 19922 3296
rect 19858 3236 19862 3292
rect 19862 3236 19918 3292
rect 19918 3236 19922 3292
rect 19858 3232 19922 3236
rect 19938 3292 20002 3296
rect 19938 3236 19942 3292
rect 19942 3236 19998 3292
rect 19998 3236 20002 3292
rect 19938 3232 20002 3236
rect 20018 3292 20082 3296
rect 20018 3236 20022 3292
rect 20022 3236 20078 3292
rect 20078 3236 20082 3292
rect 20018 3232 20082 3236
rect 20098 3292 20162 3296
rect 20098 3236 20102 3292
rect 20102 3236 20158 3292
rect 20158 3236 20162 3292
rect 20098 3232 20162 3236
rect 26160 3292 26224 3296
rect 26160 3236 26164 3292
rect 26164 3236 26220 3292
rect 26220 3236 26224 3292
rect 26160 3232 26224 3236
rect 26240 3292 26304 3296
rect 26240 3236 26244 3292
rect 26244 3236 26300 3292
rect 26300 3236 26304 3292
rect 26240 3232 26304 3236
rect 26320 3292 26384 3296
rect 26320 3236 26324 3292
rect 26324 3236 26380 3292
rect 26380 3236 26384 3292
rect 26320 3232 26384 3236
rect 26400 3292 26464 3296
rect 26400 3236 26404 3292
rect 26404 3236 26460 3292
rect 26460 3236 26464 3292
rect 26400 3232 26464 3236
rect 4103 2748 4167 2752
rect 4103 2692 4107 2748
rect 4107 2692 4163 2748
rect 4163 2692 4167 2748
rect 4103 2688 4167 2692
rect 4183 2748 4247 2752
rect 4183 2692 4187 2748
rect 4187 2692 4243 2748
rect 4243 2692 4247 2748
rect 4183 2688 4247 2692
rect 4263 2748 4327 2752
rect 4263 2692 4267 2748
rect 4267 2692 4323 2748
rect 4323 2692 4327 2748
rect 4263 2688 4327 2692
rect 4343 2748 4407 2752
rect 4343 2692 4347 2748
rect 4347 2692 4403 2748
rect 4403 2692 4407 2748
rect 4343 2688 4407 2692
rect 10405 2748 10469 2752
rect 10405 2692 10409 2748
rect 10409 2692 10465 2748
rect 10465 2692 10469 2748
rect 10405 2688 10469 2692
rect 10485 2748 10549 2752
rect 10485 2692 10489 2748
rect 10489 2692 10545 2748
rect 10545 2692 10549 2748
rect 10485 2688 10549 2692
rect 10565 2748 10629 2752
rect 10565 2692 10569 2748
rect 10569 2692 10625 2748
rect 10625 2692 10629 2748
rect 10565 2688 10629 2692
rect 10645 2748 10709 2752
rect 10645 2692 10649 2748
rect 10649 2692 10705 2748
rect 10705 2692 10709 2748
rect 10645 2688 10709 2692
rect 16707 2748 16771 2752
rect 16707 2692 16711 2748
rect 16711 2692 16767 2748
rect 16767 2692 16771 2748
rect 16707 2688 16771 2692
rect 16787 2748 16851 2752
rect 16787 2692 16791 2748
rect 16791 2692 16847 2748
rect 16847 2692 16851 2748
rect 16787 2688 16851 2692
rect 16867 2748 16931 2752
rect 16867 2692 16871 2748
rect 16871 2692 16927 2748
rect 16927 2692 16931 2748
rect 16867 2688 16931 2692
rect 16947 2748 17011 2752
rect 16947 2692 16951 2748
rect 16951 2692 17007 2748
rect 17007 2692 17011 2748
rect 16947 2688 17011 2692
rect 23009 2748 23073 2752
rect 23009 2692 23013 2748
rect 23013 2692 23069 2748
rect 23069 2692 23073 2748
rect 23009 2688 23073 2692
rect 23089 2748 23153 2752
rect 23089 2692 23093 2748
rect 23093 2692 23149 2748
rect 23149 2692 23153 2748
rect 23089 2688 23153 2692
rect 23169 2748 23233 2752
rect 23169 2692 23173 2748
rect 23173 2692 23229 2748
rect 23229 2692 23233 2748
rect 23169 2688 23233 2692
rect 23249 2748 23313 2752
rect 23249 2692 23253 2748
rect 23253 2692 23309 2748
rect 23309 2692 23313 2748
rect 23249 2688 23313 2692
rect 7254 2204 7318 2208
rect 7254 2148 7258 2204
rect 7258 2148 7314 2204
rect 7314 2148 7318 2204
rect 7254 2144 7318 2148
rect 7334 2204 7398 2208
rect 7334 2148 7338 2204
rect 7338 2148 7394 2204
rect 7394 2148 7398 2204
rect 7334 2144 7398 2148
rect 7414 2204 7478 2208
rect 7414 2148 7418 2204
rect 7418 2148 7474 2204
rect 7474 2148 7478 2204
rect 7414 2144 7478 2148
rect 7494 2204 7558 2208
rect 7494 2148 7498 2204
rect 7498 2148 7554 2204
rect 7554 2148 7558 2204
rect 7494 2144 7558 2148
rect 13556 2204 13620 2208
rect 13556 2148 13560 2204
rect 13560 2148 13616 2204
rect 13616 2148 13620 2204
rect 13556 2144 13620 2148
rect 13636 2204 13700 2208
rect 13636 2148 13640 2204
rect 13640 2148 13696 2204
rect 13696 2148 13700 2204
rect 13636 2144 13700 2148
rect 13716 2204 13780 2208
rect 13716 2148 13720 2204
rect 13720 2148 13776 2204
rect 13776 2148 13780 2204
rect 13716 2144 13780 2148
rect 13796 2204 13860 2208
rect 13796 2148 13800 2204
rect 13800 2148 13856 2204
rect 13856 2148 13860 2204
rect 13796 2144 13860 2148
rect 19858 2204 19922 2208
rect 19858 2148 19862 2204
rect 19862 2148 19918 2204
rect 19918 2148 19922 2204
rect 19858 2144 19922 2148
rect 19938 2204 20002 2208
rect 19938 2148 19942 2204
rect 19942 2148 19998 2204
rect 19998 2148 20002 2204
rect 19938 2144 20002 2148
rect 20018 2204 20082 2208
rect 20018 2148 20022 2204
rect 20022 2148 20078 2204
rect 20078 2148 20082 2204
rect 20018 2144 20082 2148
rect 20098 2204 20162 2208
rect 20098 2148 20102 2204
rect 20102 2148 20158 2204
rect 20158 2148 20162 2204
rect 20098 2144 20162 2148
rect 26160 2204 26224 2208
rect 26160 2148 26164 2204
rect 26164 2148 26220 2204
rect 26220 2148 26224 2204
rect 26160 2144 26224 2148
rect 26240 2204 26304 2208
rect 26240 2148 26244 2204
rect 26244 2148 26300 2204
rect 26300 2148 26304 2204
rect 26240 2144 26304 2148
rect 26320 2204 26384 2208
rect 26320 2148 26324 2204
rect 26324 2148 26380 2204
rect 26380 2148 26384 2204
rect 26320 2144 26384 2148
rect 26400 2204 26464 2208
rect 26400 2148 26404 2204
rect 26404 2148 26460 2204
rect 26460 2148 26464 2204
rect 26400 2144 26464 2148
<< metal4 >>
rect 4095 26688 4415 27248
rect 4095 26624 4103 26688
rect 4167 26624 4183 26688
rect 4247 26624 4263 26688
rect 4327 26624 4343 26688
rect 4407 26624 4415 26688
rect 4095 25600 4415 26624
rect 4095 25536 4103 25600
rect 4167 25536 4183 25600
rect 4247 25536 4263 25600
rect 4327 25536 4343 25600
rect 4407 25536 4415 25600
rect 4095 24512 4415 25536
rect 7246 27232 7566 27248
rect 7246 27168 7254 27232
rect 7318 27168 7334 27232
rect 7398 27168 7414 27232
rect 7478 27168 7494 27232
rect 7558 27168 7566 27232
rect 7246 26144 7566 27168
rect 7246 26080 7254 26144
rect 7318 26080 7334 26144
rect 7398 26080 7414 26144
rect 7478 26080 7494 26144
rect 7558 26080 7566 26144
rect 7246 25056 7566 26080
rect 7246 24992 7254 25056
rect 7318 24992 7334 25056
rect 7398 24992 7414 25056
rect 7478 24992 7494 25056
rect 7558 24992 7566 25056
rect 6499 24716 6565 24717
rect 6499 24652 6500 24716
rect 6564 24652 6565 24716
rect 6499 24651 6565 24652
rect 4095 24448 4103 24512
rect 4167 24448 4183 24512
rect 4247 24448 4263 24512
rect 4327 24448 4343 24512
rect 4407 24448 4415 24512
rect 4095 23424 4415 24448
rect 4095 23360 4103 23424
rect 4167 23360 4183 23424
rect 4247 23360 4263 23424
rect 4327 23360 4343 23424
rect 4407 23360 4415 23424
rect 4095 22336 4415 23360
rect 4095 22272 4103 22336
rect 4167 22272 4183 22336
rect 4247 22272 4263 22336
rect 4327 22272 4343 22336
rect 4407 22272 4415 22336
rect 4095 21248 4415 22272
rect 4095 21184 4103 21248
rect 4167 21184 4183 21248
rect 4247 21184 4263 21248
rect 4327 21184 4343 21248
rect 4407 21184 4415 21248
rect 4095 20160 4415 21184
rect 4095 20096 4103 20160
rect 4167 20096 4183 20160
rect 4247 20096 4263 20160
rect 4327 20096 4343 20160
rect 4407 20096 4415 20160
rect 4095 19072 4415 20096
rect 4095 19008 4103 19072
rect 4167 19008 4183 19072
rect 4247 19008 4263 19072
rect 4327 19008 4343 19072
rect 4407 19008 4415 19072
rect 4095 17984 4415 19008
rect 4095 17920 4103 17984
rect 4167 17920 4183 17984
rect 4247 17920 4263 17984
rect 4327 17920 4343 17984
rect 4407 17920 4415 17984
rect 4095 16896 4415 17920
rect 4095 16832 4103 16896
rect 4167 16832 4183 16896
rect 4247 16832 4263 16896
rect 4327 16832 4343 16896
rect 4407 16832 4415 16896
rect 4095 15808 4415 16832
rect 4095 15744 4103 15808
rect 4167 15744 4183 15808
rect 4247 15744 4263 15808
rect 4327 15744 4343 15808
rect 4407 15744 4415 15808
rect 4095 14720 4415 15744
rect 6502 14925 6562 24651
rect 7246 23968 7566 24992
rect 7246 23904 7254 23968
rect 7318 23904 7334 23968
rect 7398 23904 7414 23968
rect 7478 23904 7494 23968
rect 7558 23904 7566 23968
rect 7246 22880 7566 23904
rect 7246 22816 7254 22880
rect 7318 22816 7334 22880
rect 7398 22816 7414 22880
rect 7478 22816 7494 22880
rect 7558 22816 7566 22880
rect 7246 21792 7566 22816
rect 7246 21728 7254 21792
rect 7318 21728 7334 21792
rect 7398 21728 7414 21792
rect 7478 21728 7494 21792
rect 7558 21728 7566 21792
rect 7246 20704 7566 21728
rect 7246 20640 7254 20704
rect 7318 20640 7334 20704
rect 7398 20640 7414 20704
rect 7478 20640 7494 20704
rect 7558 20640 7566 20704
rect 7246 19616 7566 20640
rect 7246 19552 7254 19616
rect 7318 19552 7334 19616
rect 7398 19552 7414 19616
rect 7478 19552 7494 19616
rect 7558 19552 7566 19616
rect 7246 18528 7566 19552
rect 7246 18464 7254 18528
rect 7318 18464 7334 18528
rect 7398 18464 7414 18528
rect 7478 18464 7494 18528
rect 7558 18464 7566 18528
rect 7246 17440 7566 18464
rect 7246 17376 7254 17440
rect 7318 17376 7334 17440
rect 7398 17376 7414 17440
rect 7478 17376 7494 17440
rect 7558 17376 7566 17440
rect 7246 16352 7566 17376
rect 7246 16288 7254 16352
rect 7318 16288 7334 16352
rect 7398 16288 7414 16352
rect 7478 16288 7494 16352
rect 7558 16288 7566 16352
rect 7246 15264 7566 16288
rect 7246 15200 7254 15264
rect 7318 15200 7334 15264
rect 7398 15200 7414 15264
rect 7478 15200 7494 15264
rect 7558 15200 7566 15264
rect 6499 14924 6565 14925
rect 6499 14860 6500 14924
rect 6564 14860 6565 14924
rect 6499 14859 6565 14860
rect 4095 14656 4103 14720
rect 4167 14656 4183 14720
rect 4247 14656 4263 14720
rect 4327 14656 4343 14720
rect 4407 14656 4415 14720
rect 4095 13632 4415 14656
rect 4095 13568 4103 13632
rect 4167 13568 4183 13632
rect 4247 13568 4263 13632
rect 4327 13568 4343 13632
rect 4407 13568 4415 13632
rect 4095 12544 4415 13568
rect 4095 12480 4103 12544
rect 4167 12480 4183 12544
rect 4247 12480 4263 12544
rect 4327 12480 4343 12544
rect 4407 12480 4415 12544
rect 4095 11456 4415 12480
rect 4095 11392 4103 11456
rect 4167 11392 4183 11456
rect 4247 11392 4263 11456
rect 4327 11392 4343 11456
rect 4407 11392 4415 11456
rect 4095 10368 4415 11392
rect 4095 10304 4103 10368
rect 4167 10304 4183 10368
rect 4247 10304 4263 10368
rect 4327 10304 4343 10368
rect 4407 10304 4415 10368
rect 4095 9280 4415 10304
rect 4095 9216 4103 9280
rect 4167 9216 4183 9280
rect 4247 9216 4263 9280
rect 4327 9216 4343 9280
rect 4407 9216 4415 9280
rect 4095 8192 4415 9216
rect 4095 8128 4103 8192
rect 4167 8128 4183 8192
rect 4247 8128 4263 8192
rect 4327 8128 4343 8192
rect 4407 8128 4415 8192
rect 4095 7104 4415 8128
rect 4095 7040 4103 7104
rect 4167 7040 4183 7104
rect 4247 7040 4263 7104
rect 4327 7040 4343 7104
rect 4407 7040 4415 7104
rect 4095 6016 4415 7040
rect 4095 5952 4103 6016
rect 4167 5952 4183 6016
rect 4247 5952 4263 6016
rect 4327 5952 4343 6016
rect 4407 5952 4415 6016
rect 4095 4928 4415 5952
rect 4095 4864 4103 4928
rect 4167 4864 4183 4928
rect 4247 4864 4263 4928
rect 4327 4864 4343 4928
rect 4407 4864 4415 4928
rect 4095 3840 4415 4864
rect 4095 3776 4103 3840
rect 4167 3776 4183 3840
rect 4247 3776 4263 3840
rect 4327 3776 4343 3840
rect 4407 3776 4415 3840
rect 4095 2752 4415 3776
rect 4095 2688 4103 2752
rect 4167 2688 4183 2752
rect 4247 2688 4263 2752
rect 4327 2688 4343 2752
rect 4407 2688 4415 2752
rect 4095 2128 4415 2688
rect 7246 14176 7566 15200
rect 7246 14112 7254 14176
rect 7318 14112 7334 14176
rect 7398 14112 7414 14176
rect 7478 14112 7494 14176
rect 7558 14112 7566 14176
rect 7246 13088 7566 14112
rect 7246 13024 7254 13088
rect 7318 13024 7334 13088
rect 7398 13024 7414 13088
rect 7478 13024 7494 13088
rect 7558 13024 7566 13088
rect 7246 12000 7566 13024
rect 7246 11936 7254 12000
rect 7318 11936 7334 12000
rect 7398 11936 7414 12000
rect 7478 11936 7494 12000
rect 7558 11936 7566 12000
rect 7246 10912 7566 11936
rect 7246 10848 7254 10912
rect 7318 10848 7334 10912
rect 7398 10848 7414 10912
rect 7478 10848 7494 10912
rect 7558 10848 7566 10912
rect 7246 9824 7566 10848
rect 7246 9760 7254 9824
rect 7318 9760 7334 9824
rect 7398 9760 7414 9824
rect 7478 9760 7494 9824
rect 7558 9760 7566 9824
rect 7246 8736 7566 9760
rect 7246 8672 7254 8736
rect 7318 8672 7334 8736
rect 7398 8672 7414 8736
rect 7478 8672 7494 8736
rect 7558 8672 7566 8736
rect 7246 7648 7566 8672
rect 7246 7584 7254 7648
rect 7318 7584 7334 7648
rect 7398 7584 7414 7648
rect 7478 7584 7494 7648
rect 7558 7584 7566 7648
rect 7246 6560 7566 7584
rect 7246 6496 7254 6560
rect 7318 6496 7334 6560
rect 7398 6496 7414 6560
rect 7478 6496 7494 6560
rect 7558 6496 7566 6560
rect 7246 5472 7566 6496
rect 7246 5408 7254 5472
rect 7318 5408 7334 5472
rect 7398 5408 7414 5472
rect 7478 5408 7494 5472
rect 7558 5408 7566 5472
rect 7246 4384 7566 5408
rect 7246 4320 7254 4384
rect 7318 4320 7334 4384
rect 7398 4320 7414 4384
rect 7478 4320 7494 4384
rect 7558 4320 7566 4384
rect 7246 3296 7566 4320
rect 7246 3232 7254 3296
rect 7318 3232 7334 3296
rect 7398 3232 7414 3296
rect 7478 3232 7494 3296
rect 7558 3232 7566 3296
rect 7246 2208 7566 3232
rect 7246 2144 7254 2208
rect 7318 2144 7334 2208
rect 7398 2144 7414 2208
rect 7478 2144 7494 2208
rect 7558 2144 7566 2208
rect 7246 2128 7566 2144
rect 10397 26688 10717 27248
rect 10397 26624 10405 26688
rect 10469 26624 10485 26688
rect 10549 26624 10565 26688
rect 10629 26624 10645 26688
rect 10709 26624 10717 26688
rect 10397 25600 10717 26624
rect 10397 25536 10405 25600
rect 10469 25536 10485 25600
rect 10549 25536 10565 25600
rect 10629 25536 10645 25600
rect 10709 25536 10717 25600
rect 10397 24512 10717 25536
rect 10397 24448 10405 24512
rect 10469 24448 10485 24512
rect 10549 24448 10565 24512
rect 10629 24448 10645 24512
rect 10709 24448 10717 24512
rect 10397 23424 10717 24448
rect 10397 23360 10405 23424
rect 10469 23360 10485 23424
rect 10549 23360 10565 23424
rect 10629 23360 10645 23424
rect 10709 23360 10717 23424
rect 10397 22336 10717 23360
rect 10397 22272 10405 22336
rect 10469 22272 10485 22336
rect 10549 22272 10565 22336
rect 10629 22272 10645 22336
rect 10709 22272 10717 22336
rect 10397 21248 10717 22272
rect 10397 21184 10405 21248
rect 10469 21184 10485 21248
rect 10549 21184 10565 21248
rect 10629 21184 10645 21248
rect 10709 21184 10717 21248
rect 10397 20160 10717 21184
rect 10397 20096 10405 20160
rect 10469 20096 10485 20160
rect 10549 20096 10565 20160
rect 10629 20096 10645 20160
rect 10709 20096 10717 20160
rect 10397 19072 10717 20096
rect 10397 19008 10405 19072
rect 10469 19008 10485 19072
rect 10549 19008 10565 19072
rect 10629 19008 10645 19072
rect 10709 19008 10717 19072
rect 10397 17984 10717 19008
rect 10397 17920 10405 17984
rect 10469 17920 10485 17984
rect 10549 17920 10565 17984
rect 10629 17920 10645 17984
rect 10709 17920 10717 17984
rect 10397 16896 10717 17920
rect 10397 16832 10405 16896
rect 10469 16832 10485 16896
rect 10549 16832 10565 16896
rect 10629 16832 10645 16896
rect 10709 16832 10717 16896
rect 10397 15808 10717 16832
rect 10397 15744 10405 15808
rect 10469 15744 10485 15808
rect 10549 15744 10565 15808
rect 10629 15744 10645 15808
rect 10709 15744 10717 15808
rect 10397 14720 10717 15744
rect 10397 14656 10405 14720
rect 10469 14656 10485 14720
rect 10549 14656 10565 14720
rect 10629 14656 10645 14720
rect 10709 14656 10717 14720
rect 10397 13632 10717 14656
rect 10397 13568 10405 13632
rect 10469 13568 10485 13632
rect 10549 13568 10565 13632
rect 10629 13568 10645 13632
rect 10709 13568 10717 13632
rect 10397 12544 10717 13568
rect 10397 12480 10405 12544
rect 10469 12480 10485 12544
rect 10549 12480 10565 12544
rect 10629 12480 10645 12544
rect 10709 12480 10717 12544
rect 10397 11456 10717 12480
rect 10397 11392 10405 11456
rect 10469 11392 10485 11456
rect 10549 11392 10565 11456
rect 10629 11392 10645 11456
rect 10709 11392 10717 11456
rect 10397 10368 10717 11392
rect 10397 10304 10405 10368
rect 10469 10304 10485 10368
rect 10549 10304 10565 10368
rect 10629 10304 10645 10368
rect 10709 10304 10717 10368
rect 10397 9280 10717 10304
rect 10397 9216 10405 9280
rect 10469 9216 10485 9280
rect 10549 9216 10565 9280
rect 10629 9216 10645 9280
rect 10709 9216 10717 9280
rect 10397 8192 10717 9216
rect 10397 8128 10405 8192
rect 10469 8128 10485 8192
rect 10549 8128 10565 8192
rect 10629 8128 10645 8192
rect 10709 8128 10717 8192
rect 10397 7104 10717 8128
rect 10397 7040 10405 7104
rect 10469 7040 10485 7104
rect 10549 7040 10565 7104
rect 10629 7040 10645 7104
rect 10709 7040 10717 7104
rect 10397 6016 10717 7040
rect 10397 5952 10405 6016
rect 10469 5952 10485 6016
rect 10549 5952 10565 6016
rect 10629 5952 10645 6016
rect 10709 5952 10717 6016
rect 10397 4928 10717 5952
rect 10397 4864 10405 4928
rect 10469 4864 10485 4928
rect 10549 4864 10565 4928
rect 10629 4864 10645 4928
rect 10709 4864 10717 4928
rect 10397 3840 10717 4864
rect 10397 3776 10405 3840
rect 10469 3776 10485 3840
rect 10549 3776 10565 3840
rect 10629 3776 10645 3840
rect 10709 3776 10717 3840
rect 10397 2752 10717 3776
rect 10397 2688 10405 2752
rect 10469 2688 10485 2752
rect 10549 2688 10565 2752
rect 10629 2688 10645 2752
rect 10709 2688 10717 2752
rect 10397 2128 10717 2688
rect 13548 27232 13868 27248
rect 13548 27168 13556 27232
rect 13620 27168 13636 27232
rect 13700 27168 13716 27232
rect 13780 27168 13796 27232
rect 13860 27168 13868 27232
rect 13548 26144 13868 27168
rect 13548 26080 13556 26144
rect 13620 26080 13636 26144
rect 13700 26080 13716 26144
rect 13780 26080 13796 26144
rect 13860 26080 13868 26144
rect 13548 25056 13868 26080
rect 13548 24992 13556 25056
rect 13620 24992 13636 25056
rect 13700 24992 13716 25056
rect 13780 24992 13796 25056
rect 13860 24992 13868 25056
rect 13548 23968 13868 24992
rect 13548 23904 13556 23968
rect 13620 23904 13636 23968
rect 13700 23904 13716 23968
rect 13780 23904 13796 23968
rect 13860 23904 13868 23968
rect 13548 22880 13868 23904
rect 13548 22816 13556 22880
rect 13620 22816 13636 22880
rect 13700 22816 13716 22880
rect 13780 22816 13796 22880
rect 13860 22816 13868 22880
rect 13548 21792 13868 22816
rect 13548 21728 13556 21792
rect 13620 21728 13636 21792
rect 13700 21728 13716 21792
rect 13780 21728 13796 21792
rect 13860 21728 13868 21792
rect 13548 20704 13868 21728
rect 13548 20640 13556 20704
rect 13620 20640 13636 20704
rect 13700 20640 13716 20704
rect 13780 20640 13796 20704
rect 13860 20640 13868 20704
rect 13548 19616 13868 20640
rect 13548 19552 13556 19616
rect 13620 19552 13636 19616
rect 13700 19552 13716 19616
rect 13780 19552 13796 19616
rect 13860 19552 13868 19616
rect 13548 18528 13868 19552
rect 13548 18464 13556 18528
rect 13620 18464 13636 18528
rect 13700 18464 13716 18528
rect 13780 18464 13796 18528
rect 13860 18464 13868 18528
rect 13548 17440 13868 18464
rect 13548 17376 13556 17440
rect 13620 17376 13636 17440
rect 13700 17376 13716 17440
rect 13780 17376 13796 17440
rect 13860 17376 13868 17440
rect 13548 16352 13868 17376
rect 13548 16288 13556 16352
rect 13620 16288 13636 16352
rect 13700 16288 13716 16352
rect 13780 16288 13796 16352
rect 13860 16288 13868 16352
rect 13548 15264 13868 16288
rect 13548 15200 13556 15264
rect 13620 15200 13636 15264
rect 13700 15200 13716 15264
rect 13780 15200 13796 15264
rect 13860 15200 13868 15264
rect 13548 14176 13868 15200
rect 13548 14112 13556 14176
rect 13620 14112 13636 14176
rect 13700 14112 13716 14176
rect 13780 14112 13796 14176
rect 13860 14112 13868 14176
rect 13548 13088 13868 14112
rect 13548 13024 13556 13088
rect 13620 13024 13636 13088
rect 13700 13024 13716 13088
rect 13780 13024 13796 13088
rect 13860 13024 13868 13088
rect 13548 12000 13868 13024
rect 13548 11936 13556 12000
rect 13620 11936 13636 12000
rect 13700 11936 13716 12000
rect 13780 11936 13796 12000
rect 13860 11936 13868 12000
rect 13548 10912 13868 11936
rect 13548 10848 13556 10912
rect 13620 10848 13636 10912
rect 13700 10848 13716 10912
rect 13780 10848 13796 10912
rect 13860 10848 13868 10912
rect 13548 9824 13868 10848
rect 13548 9760 13556 9824
rect 13620 9760 13636 9824
rect 13700 9760 13716 9824
rect 13780 9760 13796 9824
rect 13860 9760 13868 9824
rect 13548 8736 13868 9760
rect 13548 8672 13556 8736
rect 13620 8672 13636 8736
rect 13700 8672 13716 8736
rect 13780 8672 13796 8736
rect 13860 8672 13868 8736
rect 13548 7648 13868 8672
rect 13548 7584 13556 7648
rect 13620 7584 13636 7648
rect 13700 7584 13716 7648
rect 13780 7584 13796 7648
rect 13860 7584 13868 7648
rect 13548 6560 13868 7584
rect 13548 6496 13556 6560
rect 13620 6496 13636 6560
rect 13700 6496 13716 6560
rect 13780 6496 13796 6560
rect 13860 6496 13868 6560
rect 13548 5472 13868 6496
rect 13548 5408 13556 5472
rect 13620 5408 13636 5472
rect 13700 5408 13716 5472
rect 13780 5408 13796 5472
rect 13860 5408 13868 5472
rect 13548 4384 13868 5408
rect 13548 4320 13556 4384
rect 13620 4320 13636 4384
rect 13700 4320 13716 4384
rect 13780 4320 13796 4384
rect 13860 4320 13868 4384
rect 13548 3296 13868 4320
rect 13548 3232 13556 3296
rect 13620 3232 13636 3296
rect 13700 3232 13716 3296
rect 13780 3232 13796 3296
rect 13860 3232 13868 3296
rect 13548 2208 13868 3232
rect 13548 2144 13556 2208
rect 13620 2144 13636 2208
rect 13700 2144 13716 2208
rect 13780 2144 13796 2208
rect 13860 2144 13868 2208
rect 13548 2128 13868 2144
rect 16699 26688 17019 27248
rect 16699 26624 16707 26688
rect 16771 26624 16787 26688
rect 16851 26624 16867 26688
rect 16931 26624 16947 26688
rect 17011 26624 17019 26688
rect 16699 25600 17019 26624
rect 16699 25536 16707 25600
rect 16771 25536 16787 25600
rect 16851 25536 16867 25600
rect 16931 25536 16947 25600
rect 17011 25536 17019 25600
rect 16699 24512 17019 25536
rect 16699 24448 16707 24512
rect 16771 24448 16787 24512
rect 16851 24448 16867 24512
rect 16931 24448 16947 24512
rect 17011 24448 17019 24512
rect 16699 23424 17019 24448
rect 16699 23360 16707 23424
rect 16771 23360 16787 23424
rect 16851 23360 16867 23424
rect 16931 23360 16947 23424
rect 17011 23360 17019 23424
rect 16699 22336 17019 23360
rect 16699 22272 16707 22336
rect 16771 22272 16787 22336
rect 16851 22272 16867 22336
rect 16931 22272 16947 22336
rect 17011 22272 17019 22336
rect 16699 21248 17019 22272
rect 16699 21184 16707 21248
rect 16771 21184 16787 21248
rect 16851 21184 16867 21248
rect 16931 21184 16947 21248
rect 17011 21184 17019 21248
rect 16699 20160 17019 21184
rect 16699 20096 16707 20160
rect 16771 20096 16787 20160
rect 16851 20096 16867 20160
rect 16931 20096 16947 20160
rect 17011 20096 17019 20160
rect 16699 19072 17019 20096
rect 16699 19008 16707 19072
rect 16771 19008 16787 19072
rect 16851 19008 16867 19072
rect 16931 19008 16947 19072
rect 17011 19008 17019 19072
rect 16699 17984 17019 19008
rect 16699 17920 16707 17984
rect 16771 17920 16787 17984
rect 16851 17920 16867 17984
rect 16931 17920 16947 17984
rect 17011 17920 17019 17984
rect 16699 16896 17019 17920
rect 16699 16832 16707 16896
rect 16771 16832 16787 16896
rect 16851 16832 16867 16896
rect 16931 16832 16947 16896
rect 17011 16832 17019 16896
rect 16699 15808 17019 16832
rect 16699 15744 16707 15808
rect 16771 15744 16787 15808
rect 16851 15744 16867 15808
rect 16931 15744 16947 15808
rect 17011 15744 17019 15808
rect 16699 14720 17019 15744
rect 16699 14656 16707 14720
rect 16771 14656 16787 14720
rect 16851 14656 16867 14720
rect 16931 14656 16947 14720
rect 17011 14656 17019 14720
rect 16699 13632 17019 14656
rect 16699 13568 16707 13632
rect 16771 13568 16787 13632
rect 16851 13568 16867 13632
rect 16931 13568 16947 13632
rect 17011 13568 17019 13632
rect 16699 12544 17019 13568
rect 16699 12480 16707 12544
rect 16771 12480 16787 12544
rect 16851 12480 16867 12544
rect 16931 12480 16947 12544
rect 17011 12480 17019 12544
rect 16699 11456 17019 12480
rect 16699 11392 16707 11456
rect 16771 11392 16787 11456
rect 16851 11392 16867 11456
rect 16931 11392 16947 11456
rect 17011 11392 17019 11456
rect 16699 10368 17019 11392
rect 16699 10304 16707 10368
rect 16771 10304 16787 10368
rect 16851 10304 16867 10368
rect 16931 10304 16947 10368
rect 17011 10304 17019 10368
rect 16699 9280 17019 10304
rect 16699 9216 16707 9280
rect 16771 9216 16787 9280
rect 16851 9216 16867 9280
rect 16931 9216 16947 9280
rect 17011 9216 17019 9280
rect 16699 8192 17019 9216
rect 16699 8128 16707 8192
rect 16771 8128 16787 8192
rect 16851 8128 16867 8192
rect 16931 8128 16947 8192
rect 17011 8128 17019 8192
rect 16699 7104 17019 8128
rect 16699 7040 16707 7104
rect 16771 7040 16787 7104
rect 16851 7040 16867 7104
rect 16931 7040 16947 7104
rect 17011 7040 17019 7104
rect 16699 6016 17019 7040
rect 16699 5952 16707 6016
rect 16771 5952 16787 6016
rect 16851 5952 16867 6016
rect 16931 5952 16947 6016
rect 17011 5952 17019 6016
rect 16699 4928 17019 5952
rect 16699 4864 16707 4928
rect 16771 4864 16787 4928
rect 16851 4864 16867 4928
rect 16931 4864 16947 4928
rect 17011 4864 17019 4928
rect 16699 3840 17019 4864
rect 16699 3776 16707 3840
rect 16771 3776 16787 3840
rect 16851 3776 16867 3840
rect 16931 3776 16947 3840
rect 17011 3776 17019 3840
rect 16699 2752 17019 3776
rect 16699 2688 16707 2752
rect 16771 2688 16787 2752
rect 16851 2688 16867 2752
rect 16931 2688 16947 2752
rect 17011 2688 17019 2752
rect 16699 2128 17019 2688
rect 19850 27232 20170 27248
rect 19850 27168 19858 27232
rect 19922 27168 19938 27232
rect 20002 27168 20018 27232
rect 20082 27168 20098 27232
rect 20162 27168 20170 27232
rect 19850 26144 20170 27168
rect 19850 26080 19858 26144
rect 19922 26080 19938 26144
rect 20002 26080 20018 26144
rect 20082 26080 20098 26144
rect 20162 26080 20170 26144
rect 19850 25056 20170 26080
rect 19850 24992 19858 25056
rect 19922 24992 19938 25056
rect 20002 24992 20018 25056
rect 20082 24992 20098 25056
rect 20162 24992 20170 25056
rect 19850 23968 20170 24992
rect 19850 23904 19858 23968
rect 19922 23904 19938 23968
rect 20002 23904 20018 23968
rect 20082 23904 20098 23968
rect 20162 23904 20170 23968
rect 19850 22880 20170 23904
rect 19850 22816 19858 22880
rect 19922 22816 19938 22880
rect 20002 22816 20018 22880
rect 20082 22816 20098 22880
rect 20162 22816 20170 22880
rect 19850 21792 20170 22816
rect 19850 21728 19858 21792
rect 19922 21728 19938 21792
rect 20002 21728 20018 21792
rect 20082 21728 20098 21792
rect 20162 21728 20170 21792
rect 19850 20704 20170 21728
rect 19850 20640 19858 20704
rect 19922 20640 19938 20704
rect 20002 20640 20018 20704
rect 20082 20640 20098 20704
rect 20162 20640 20170 20704
rect 19850 19616 20170 20640
rect 19850 19552 19858 19616
rect 19922 19552 19938 19616
rect 20002 19552 20018 19616
rect 20082 19552 20098 19616
rect 20162 19552 20170 19616
rect 19850 18528 20170 19552
rect 19850 18464 19858 18528
rect 19922 18464 19938 18528
rect 20002 18464 20018 18528
rect 20082 18464 20098 18528
rect 20162 18464 20170 18528
rect 19850 17440 20170 18464
rect 19850 17376 19858 17440
rect 19922 17376 19938 17440
rect 20002 17376 20018 17440
rect 20082 17376 20098 17440
rect 20162 17376 20170 17440
rect 19850 16352 20170 17376
rect 19850 16288 19858 16352
rect 19922 16288 19938 16352
rect 20002 16288 20018 16352
rect 20082 16288 20098 16352
rect 20162 16288 20170 16352
rect 19850 15264 20170 16288
rect 19850 15200 19858 15264
rect 19922 15200 19938 15264
rect 20002 15200 20018 15264
rect 20082 15200 20098 15264
rect 20162 15200 20170 15264
rect 19850 14176 20170 15200
rect 19850 14112 19858 14176
rect 19922 14112 19938 14176
rect 20002 14112 20018 14176
rect 20082 14112 20098 14176
rect 20162 14112 20170 14176
rect 19850 13088 20170 14112
rect 19850 13024 19858 13088
rect 19922 13024 19938 13088
rect 20002 13024 20018 13088
rect 20082 13024 20098 13088
rect 20162 13024 20170 13088
rect 19850 12000 20170 13024
rect 19850 11936 19858 12000
rect 19922 11936 19938 12000
rect 20002 11936 20018 12000
rect 20082 11936 20098 12000
rect 20162 11936 20170 12000
rect 19850 10912 20170 11936
rect 19850 10848 19858 10912
rect 19922 10848 19938 10912
rect 20002 10848 20018 10912
rect 20082 10848 20098 10912
rect 20162 10848 20170 10912
rect 19850 9824 20170 10848
rect 19850 9760 19858 9824
rect 19922 9760 19938 9824
rect 20002 9760 20018 9824
rect 20082 9760 20098 9824
rect 20162 9760 20170 9824
rect 19850 8736 20170 9760
rect 19850 8672 19858 8736
rect 19922 8672 19938 8736
rect 20002 8672 20018 8736
rect 20082 8672 20098 8736
rect 20162 8672 20170 8736
rect 19850 7648 20170 8672
rect 19850 7584 19858 7648
rect 19922 7584 19938 7648
rect 20002 7584 20018 7648
rect 20082 7584 20098 7648
rect 20162 7584 20170 7648
rect 19850 6560 20170 7584
rect 19850 6496 19858 6560
rect 19922 6496 19938 6560
rect 20002 6496 20018 6560
rect 20082 6496 20098 6560
rect 20162 6496 20170 6560
rect 19850 5472 20170 6496
rect 19850 5408 19858 5472
rect 19922 5408 19938 5472
rect 20002 5408 20018 5472
rect 20082 5408 20098 5472
rect 20162 5408 20170 5472
rect 19850 4384 20170 5408
rect 19850 4320 19858 4384
rect 19922 4320 19938 4384
rect 20002 4320 20018 4384
rect 20082 4320 20098 4384
rect 20162 4320 20170 4384
rect 19850 3296 20170 4320
rect 19850 3232 19858 3296
rect 19922 3232 19938 3296
rect 20002 3232 20018 3296
rect 20082 3232 20098 3296
rect 20162 3232 20170 3296
rect 19850 2208 20170 3232
rect 19850 2144 19858 2208
rect 19922 2144 19938 2208
rect 20002 2144 20018 2208
rect 20082 2144 20098 2208
rect 20162 2144 20170 2208
rect 19850 2128 20170 2144
rect 23001 26688 23321 27248
rect 23001 26624 23009 26688
rect 23073 26624 23089 26688
rect 23153 26624 23169 26688
rect 23233 26624 23249 26688
rect 23313 26624 23321 26688
rect 23001 25600 23321 26624
rect 23001 25536 23009 25600
rect 23073 25536 23089 25600
rect 23153 25536 23169 25600
rect 23233 25536 23249 25600
rect 23313 25536 23321 25600
rect 23001 24512 23321 25536
rect 23001 24448 23009 24512
rect 23073 24448 23089 24512
rect 23153 24448 23169 24512
rect 23233 24448 23249 24512
rect 23313 24448 23321 24512
rect 23001 23424 23321 24448
rect 23001 23360 23009 23424
rect 23073 23360 23089 23424
rect 23153 23360 23169 23424
rect 23233 23360 23249 23424
rect 23313 23360 23321 23424
rect 23001 22336 23321 23360
rect 23001 22272 23009 22336
rect 23073 22272 23089 22336
rect 23153 22272 23169 22336
rect 23233 22272 23249 22336
rect 23313 22272 23321 22336
rect 23001 21248 23321 22272
rect 23001 21184 23009 21248
rect 23073 21184 23089 21248
rect 23153 21184 23169 21248
rect 23233 21184 23249 21248
rect 23313 21184 23321 21248
rect 23001 20160 23321 21184
rect 23001 20096 23009 20160
rect 23073 20096 23089 20160
rect 23153 20096 23169 20160
rect 23233 20096 23249 20160
rect 23313 20096 23321 20160
rect 23001 19072 23321 20096
rect 23001 19008 23009 19072
rect 23073 19008 23089 19072
rect 23153 19008 23169 19072
rect 23233 19008 23249 19072
rect 23313 19008 23321 19072
rect 23001 17984 23321 19008
rect 23001 17920 23009 17984
rect 23073 17920 23089 17984
rect 23153 17920 23169 17984
rect 23233 17920 23249 17984
rect 23313 17920 23321 17984
rect 23001 16896 23321 17920
rect 23001 16832 23009 16896
rect 23073 16832 23089 16896
rect 23153 16832 23169 16896
rect 23233 16832 23249 16896
rect 23313 16832 23321 16896
rect 23001 15808 23321 16832
rect 23001 15744 23009 15808
rect 23073 15744 23089 15808
rect 23153 15744 23169 15808
rect 23233 15744 23249 15808
rect 23313 15744 23321 15808
rect 23001 14720 23321 15744
rect 23001 14656 23009 14720
rect 23073 14656 23089 14720
rect 23153 14656 23169 14720
rect 23233 14656 23249 14720
rect 23313 14656 23321 14720
rect 23001 13632 23321 14656
rect 23001 13568 23009 13632
rect 23073 13568 23089 13632
rect 23153 13568 23169 13632
rect 23233 13568 23249 13632
rect 23313 13568 23321 13632
rect 23001 12544 23321 13568
rect 23001 12480 23009 12544
rect 23073 12480 23089 12544
rect 23153 12480 23169 12544
rect 23233 12480 23249 12544
rect 23313 12480 23321 12544
rect 23001 11456 23321 12480
rect 23001 11392 23009 11456
rect 23073 11392 23089 11456
rect 23153 11392 23169 11456
rect 23233 11392 23249 11456
rect 23313 11392 23321 11456
rect 23001 10368 23321 11392
rect 23001 10304 23009 10368
rect 23073 10304 23089 10368
rect 23153 10304 23169 10368
rect 23233 10304 23249 10368
rect 23313 10304 23321 10368
rect 23001 9280 23321 10304
rect 23001 9216 23009 9280
rect 23073 9216 23089 9280
rect 23153 9216 23169 9280
rect 23233 9216 23249 9280
rect 23313 9216 23321 9280
rect 23001 8192 23321 9216
rect 23001 8128 23009 8192
rect 23073 8128 23089 8192
rect 23153 8128 23169 8192
rect 23233 8128 23249 8192
rect 23313 8128 23321 8192
rect 23001 7104 23321 8128
rect 23001 7040 23009 7104
rect 23073 7040 23089 7104
rect 23153 7040 23169 7104
rect 23233 7040 23249 7104
rect 23313 7040 23321 7104
rect 23001 6016 23321 7040
rect 23001 5952 23009 6016
rect 23073 5952 23089 6016
rect 23153 5952 23169 6016
rect 23233 5952 23249 6016
rect 23313 5952 23321 6016
rect 23001 4928 23321 5952
rect 23001 4864 23009 4928
rect 23073 4864 23089 4928
rect 23153 4864 23169 4928
rect 23233 4864 23249 4928
rect 23313 4864 23321 4928
rect 23001 3840 23321 4864
rect 23001 3776 23009 3840
rect 23073 3776 23089 3840
rect 23153 3776 23169 3840
rect 23233 3776 23249 3840
rect 23313 3776 23321 3840
rect 23001 2752 23321 3776
rect 23001 2688 23009 2752
rect 23073 2688 23089 2752
rect 23153 2688 23169 2752
rect 23233 2688 23249 2752
rect 23313 2688 23321 2752
rect 23001 2128 23321 2688
rect 26152 27232 26472 27248
rect 26152 27168 26160 27232
rect 26224 27168 26240 27232
rect 26304 27168 26320 27232
rect 26384 27168 26400 27232
rect 26464 27168 26472 27232
rect 26152 26144 26472 27168
rect 26152 26080 26160 26144
rect 26224 26080 26240 26144
rect 26304 26080 26320 26144
rect 26384 26080 26400 26144
rect 26464 26080 26472 26144
rect 26152 25056 26472 26080
rect 26152 24992 26160 25056
rect 26224 24992 26240 25056
rect 26304 24992 26320 25056
rect 26384 24992 26400 25056
rect 26464 24992 26472 25056
rect 26152 23968 26472 24992
rect 26152 23904 26160 23968
rect 26224 23904 26240 23968
rect 26304 23904 26320 23968
rect 26384 23904 26400 23968
rect 26464 23904 26472 23968
rect 26152 22880 26472 23904
rect 26152 22816 26160 22880
rect 26224 22816 26240 22880
rect 26304 22816 26320 22880
rect 26384 22816 26400 22880
rect 26464 22816 26472 22880
rect 26152 21792 26472 22816
rect 26152 21728 26160 21792
rect 26224 21728 26240 21792
rect 26304 21728 26320 21792
rect 26384 21728 26400 21792
rect 26464 21728 26472 21792
rect 26152 20704 26472 21728
rect 26152 20640 26160 20704
rect 26224 20640 26240 20704
rect 26304 20640 26320 20704
rect 26384 20640 26400 20704
rect 26464 20640 26472 20704
rect 26152 19616 26472 20640
rect 26152 19552 26160 19616
rect 26224 19552 26240 19616
rect 26304 19552 26320 19616
rect 26384 19552 26400 19616
rect 26464 19552 26472 19616
rect 26152 18528 26472 19552
rect 26152 18464 26160 18528
rect 26224 18464 26240 18528
rect 26304 18464 26320 18528
rect 26384 18464 26400 18528
rect 26464 18464 26472 18528
rect 26152 17440 26472 18464
rect 26152 17376 26160 17440
rect 26224 17376 26240 17440
rect 26304 17376 26320 17440
rect 26384 17376 26400 17440
rect 26464 17376 26472 17440
rect 26152 16352 26472 17376
rect 26152 16288 26160 16352
rect 26224 16288 26240 16352
rect 26304 16288 26320 16352
rect 26384 16288 26400 16352
rect 26464 16288 26472 16352
rect 26152 15264 26472 16288
rect 26152 15200 26160 15264
rect 26224 15200 26240 15264
rect 26304 15200 26320 15264
rect 26384 15200 26400 15264
rect 26464 15200 26472 15264
rect 26152 14176 26472 15200
rect 26152 14112 26160 14176
rect 26224 14112 26240 14176
rect 26304 14112 26320 14176
rect 26384 14112 26400 14176
rect 26464 14112 26472 14176
rect 26152 13088 26472 14112
rect 26152 13024 26160 13088
rect 26224 13024 26240 13088
rect 26304 13024 26320 13088
rect 26384 13024 26400 13088
rect 26464 13024 26472 13088
rect 26152 12000 26472 13024
rect 26152 11936 26160 12000
rect 26224 11936 26240 12000
rect 26304 11936 26320 12000
rect 26384 11936 26400 12000
rect 26464 11936 26472 12000
rect 26152 10912 26472 11936
rect 26152 10848 26160 10912
rect 26224 10848 26240 10912
rect 26304 10848 26320 10912
rect 26384 10848 26400 10912
rect 26464 10848 26472 10912
rect 26152 9824 26472 10848
rect 26152 9760 26160 9824
rect 26224 9760 26240 9824
rect 26304 9760 26320 9824
rect 26384 9760 26400 9824
rect 26464 9760 26472 9824
rect 26152 8736 26472 9760
rect 26152 8672 26160 8736
rect 26224 8672 26240 8736
rect 26304 8672 26320 8736
rect 26384 8672 26400 8736
rect 26464 8672 26472 8736
rect 26152 7648 26472 8672
rect 26152 7584 26160 7648
rect 26224 7584 26240 7648
rect 26304 7584 26320 7648
rect 26384 7584 26400 7648
rect 26464 7584 26472 7648
rect 26152 6560 26472 7584
rect 26152 6496 26160 6560
rect 26224 6496 26240 6560
rect 26304 6496 26320 6560
rect 26384 6496 26400 6560
rect 26464 6496 26472 6560
rect 26152 5472 26472 6496
rect 26152 5408 26160 5472
rect 26224 5408 26240 5472
rect 26304 5408 26320 5472
rect 26384 5408 26400 5472
rect 26464 5408 26472 5472
rect 26152 4384 26472 5408
rect 26152 4320 26160 4384
rect 26224 4320 26240 4384
rect 26304 4320 26320 4384
rect 26384 4320 26400 4384
rect 26464 4320 26472 4384
rect 26152 3296 26472 4320
rect 26152 3232 26160 3296
rect 26224 3232 26240 3296
rect 26304 3232 26320 3296
rect 26384 3232 26400 3296
rect 26464 3232 26472 3296
rect 26152 2208 26472 3232
rect 26152 2144 26160 2208
rect 26224 2144 26240 2208
rect 26304 2144 26320 2208
rect 26384 2144 26400 2208
rect 26464 2144 26472 2208
rect 26152 2128 26472 2144
use sky130_fd_sc_hd__or2b_1  _0469_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25392 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0470_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25392 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0471_
timestamp 1688980957
transform -1 0 23092 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0472_
timestamp 1688980957
transform -1 0 21712 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0473_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21712 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0474_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24564 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0475_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25024 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0476_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25024 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0477_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23920 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0478_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0479_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20976 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0480_
timestamp 1688980957
transform 1 0 20608 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0481_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24288 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0482_
timestamp 1688980957
transform 1 0 19780 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0483_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0484_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0486_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0487_
timestamp 1688980957
transform 1 0 7176 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0488_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _0489_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20976 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0490_
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1688980957
transform -1 0 21712 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0492_
timestamp 1688980957
transform 1 0 21068 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0493_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0494_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21988 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0495_
timestamp 1688980957
transform 1 0 21804 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0496_
timestamp 1688980957
transform -1 0 22356 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0497_
timestamp 1688980957
transform 1 0 20700 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0498_
timestamp 1688980957
transform 1 0 20148 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0499_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19780 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0500_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25760 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0501_
timestamp 1688980957
transform 1 0 19320 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0502_
timestamp 1688980957
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1688980957
transform 1 0 23828 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0504_
timestamp 1688980957
transform -1 0 24932 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0505_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0506_
timestamp 1688980957
transform 1 0 20700 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0507_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23092 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0508_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1688980957
transform 1 0 14904 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0510_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0511_
timestamp 1688980957
transform -1 0 13984 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0512_
timestamp 1688980957
transform -1 0 13984 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0513_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15364 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0514_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15364 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0515_
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0516_
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0517_
timestamp 1688980957
transform 1 0 14444 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _0518_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14628 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0519_
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0520_
timestamp 1688980957
transform -1 0 25300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0521_
timestamp 1688980957
transform 1 0 16192 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _0522_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16192 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0523_
timestamp 1688980957
transform 1 0 13156 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0524_
timestamp 1688980957
transform 1 0 13156 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0525_
timestamp 1688980957
transform 1 0 14628 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_2  _0526_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14628 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _0527_
timestamp 1688980957
transform -1 0 15180 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0528_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15732 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0529_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22448 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0530_
timestamp 1688980957
transform -1 0 22908 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0531_
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _0532_
timestamp 1688980957
transform -1 0 22908 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0533_
timestamp 1688980957
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _0534_
timestamp 1688980957
transform -1 0 23644 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0535_
timestamp 1688980957
transform -1 0 21344 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0536_
timestamp 1688980957
transform -1 0 4140 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1688980957
transform 1 0 5520 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0538_
timestamp 1688980957
transform 1 0 4140 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0539_
timestamp 1688980957
transform 1 0 2392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0540_
timestamp 1688980957
transform -1 0 4784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0541_
timestamp 1688980957
transform 1 0 5060 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0542_
timestamp 1688980957
transform 1 0 2024 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0543_
timestamp 1688980957
transform -1 0 4968 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0544_
timestamp 1688980957
transform -1 0 3680 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0545_
timestamp 1688980957
transform -1 0 3036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _0546_
timestamp 1688980957
transform -1 0 4508 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0547_
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0548_
timestamp 1688980957
transform -1 0 25300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0549_
timestamp 1688980957
transform 1 0 2852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0550_
timestamp 1688980957
transform 1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _0551_
timestamp 1688980957
transform -1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0552_
timestamp 1688980957
transform 1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0553_
timestamp 1688980957
transform -1 0 4876 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_2  _0554_
timestamp 1688980957
transform 1 0 2760 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _0555_
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0556_
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1688980957
transform -1 0 20976 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0558_
timestamp 1688980957
transform -1 0 21620 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0559_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23000 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0560_
timestamp 1688980957
transform 1 0 23460 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0561_
timestamp 1688980957
transform -1 0 20792 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0562_
timestamp 1688980957
transform 1 0 20240 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_8  _0563_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__a22o_1  _0564_
timestamp 1688980957
transform 1 0 16008 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0565_
timestamp 1688980957
transform 1 0 3956 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0566_
timestamp 1688980957
transform -1 0 5612 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0567_
timestamp 1688980957
transform 1 0 6072 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0568_
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0569_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _0570_
timestamp 1688980957
transform 1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0571_
timestamp 1688980957
transform -1 0 6900 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0572_
timestamp 1688980957
transform 1 0 7176 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0573_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7636 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0574_
timestamp 1688980957
transform 1 0 4416 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o2111ai_1  _0575_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5704 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0576_
timestamp 1688980957
transform 1 0 7636 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0577_
timestamp 1688980957
transform 1 0 6348 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_4  _0578_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _0579_
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0580_
timestamp 1688980957
transform 1 0 5796 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0581_
timestamp 1688980957
transform -1 0 6992 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0582_
timestamp 1688980957
transform -1 0 14720 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0583_
timestamp 1688980957
transform -1 0 6716 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1688980957
transform 1 0 6440 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0585_
timestamp 1688980957
transform -1 0 6992 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0586_
timestamp 1688980957
transform 1 0 6900 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0587_
timestamp 1688980957
transform 1 0 4140 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _0588_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5796 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0589_
timestamp 1688980957
transform 1 0 5704 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0590_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0591_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5704 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0592_
timestamp 1688980957
transform -1 0 5704 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0593_
timestamp 1688980957
transform -1 0 4508 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0594_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4876 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0595_
timestamp 1688980957
transform -1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0596_
timestamp 1688980957
transform 1 0 4968 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0597_
timestamp 1688980957
transform 1 0 5704 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0598_
timestamp 1688980957
transform 1 0 5520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0599_
timestamp 1688980957
transform 1 0 4508 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0600_
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0601_
timestamp 1688980957
transform 1 0 7544 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0602_
timestamp 1688980957
transform -1 0 7544 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0603_
timestamp 1688980957
transform 1 0 6348 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0604_
timestamp 1688980957
transform -1 0 6256 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0605_
timestamp 1688980957
transform 1 0 6348 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0606_
timestamp 1688980957
transform 1 0 6716 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _0607_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8832 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _0608_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7912 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0609_
timestamp 1688980957
transform -1 0 6624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0610_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18492 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _0611_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17572 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0612_
timestamp 1688980957
transform 1 0 17572 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0613_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15824 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0614_
timestamp 1688980957
transform -1 0 17664 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0615_
timestamp 1688980957
transform -1 0 18124 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0616_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16928 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _0617_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16652 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _0618_
timestamp 1688980957
transform -1 0 17112 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0619_
timestamp 1688980957
transform 1 0 15456 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0620_
timestamp 1688980957
transform -1 0 16100 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_4  _0621_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1688980957
transform -1 0 16192 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0623_
timestamp 1688980957
transform 1 0 16836 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0624_
timestamp 1688980957
transform -1 0 17112 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0625_
timestamp 1688980957
transform -1 0 13616 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0626_
timestamp 1688980957
transform -1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0627_
timestamp 1688980957
transform -1 0 13156 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0628_
timestamp 1688980957
transform -1 0 12604 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0629_
timestamp 1688980957
transform -1 0 16744 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0630_
timestamp 1688980957
transform -1 0 16468 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0631_
timestamp 1688980957
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0632_
timestamp 1688980957
transform -1 0 14720 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0633_
timestamp 1688980957
transform -1 0 13156 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_4  _0634_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__a21oi_4  _0635_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0636_
timestamp 1688980957
transform -1 0 10120 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0637_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13248 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0638_
timestamp 1688980957
transform -1 0 9660 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1688980957
transform -1 0 9752 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0640_
timestamp 1688980957
transform -1 0 9660 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _0641_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8832 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0642_
timestamp 1688980957
transform -1 0 9384 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0643_
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_2  _0644_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8096 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _0645_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8832 0 1 6528
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_1  _0646_
timestamp 1688980957
transform 1 0 7544 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0647_
timestamp 1688980957
transform -1 0 13524 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0648_
timestamp 1688980957
transform 1 0 12604 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__and3b_1  _0649_
timestamp 1688980957
transform -1 0 10120 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0650_
timestamp 1688980957
transform -1 0 7636 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0651_
timestamp 1688980957
transform 1 0 4968 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0652_
timestamp 1688980957
transform 1 0 5336 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _0653_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8280 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0654_
timestamp 1688980957
transform -1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0655_
timestamp 1688980957
transform -1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0656_
timestamp 1688980957
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0657_
timestamp 1688980957
transform -1 0 13248 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _0658_
timestamp 1688980957
transform 1 0 12052 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0659_
timestamp 1688980957
transform 1 0 6900 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0660_
timestamp 1688980957
transform -1 0 7636 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _0661_
timestamp 1688980957
transform 1 0 4692 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0662_
timestamp 1688980957
transform 1 0 5060 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_4  _0663_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15640 0 -1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0664_
timestamp 1688980957
transform 1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0665_
timestamp 1688980957
transform -1 0 6808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0666_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_4  _0667_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7544 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__o21a_2  _0668_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6992 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0669_
timestamp 1688980957
transform -1 0 8648 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0670_
timestamp 1688980957
transform -1 0 6900 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0671_
timestamp 1688980957
transform -1 0 6256 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0672_
timestamp 1688980957
transform -1 0 8004 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0673_
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0674_
timestamp 1688980957
transform 1 0 6900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0675_
timestamp 1688980957
transform 1 0 7728 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _0676_
timestamp 1688980957
transform -1 0 7728 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0677_
timestamp 1688980957
transform -1 0 8832 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0678_
timestamp 1688980957
transform -1 0 7268 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0679_
timestamp 1688980957
transform 1 0 2208 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0680_
timestamp 1688980957
transform 1 0 24932 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_2  _0681_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21620 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0682_
timestamp 1688980957
transform 1 0 21804 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0683_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22448 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_4  _0684_
timestamp 1688980957
transform 1 0 21068 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__a21oi_4  _0685_
timestamp 1688980957
transform 1 0 4784 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1688980957
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0687_
timestamp 1688980957
transform 1 0 4508 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0688_
timestamp 1688980957
transform 1 0 3680 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0689_
timestamp 1688980957
transform 1 0 3312 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0690_
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0691_
timestamp 1688980957
transform 1 0 2300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0692_
timestamp 1688980957
transform 1 0 2668 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0693_
timestamp 1688980957
transform 1 0 2116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0694_
timestamp 1688980957
transform 1 0 2576 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0695_
timestamp 1688980957
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0696_
timestamp 1688980957
transform 1 0 2668 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1688980957
transform 1 0 2208 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0698_
timestamp 1688980957
transform 1 0 3680 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0699_
timestamp 1688980957
transform 1 0 2116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0700_
timestamp 1688980957
transform 1 0 2852 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0701_
timestamp 1688980957
transform 1 0 2392 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0702_
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0703_
timestamp 1688980957
transform 1 0 3128 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _0704_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_4  _0705_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19044 0 -1 16320
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _0706_
timestamp 1688980957
transform 1 0 16928 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0707_
timestamp 1688980957
transform -1 0 17020 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0708_
timestamp 1688980957
transform 1 0 17296 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0709_
timestamp 1688980957
transform -1 0 17112 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0710_
timestamp 1688980957
transform 1 0 14260 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0711_
timestamp 1688980957
transform -1 0 13984 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0712_
timestamp 1688980957
transform 1 0 14720 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0713_
timestamp 1688980957
transform -1 0 13984 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0714_
timestamp 1688980957
transform 1 0 9292 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0715_
timestamp 1688980957
transform -1 0 8832 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0716_
timestamp 1688980957
transform 1 0 9384 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0717_
timestamp 1688980957
transform 1 0 9108 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0718_
timestamp 1688980957
transform 1 0 9200 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0719_
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0720_
timestamp 1688980957
transform 1 0 9200 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0721_
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0722_
timestamp 1688980957
transform 1 0 12880 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0723_
timestamp 1688980957
transform 1 0 12604 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _0724_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20148 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _0725_
timestamp 1688980957
transform -1 0 19228 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0726_
timestamp 1688980957
transform -1 0 18124 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0727_
timestamp 1688980957
transform 1 0 18768 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0728_
timestamp 1688980957
transform -1 0 18584 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0729_
timestamp 1688980957
transform -1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0730_
timestamp 1688980957
transform 1 0 16836 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0731_
timestamp 1688980957
transform -1 0 14720 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0732_
timestamp 1688980957
transform -1 0 17572 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0733_
timestamp 1688980957
transform 1 0 17388 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0734_
timestamp 1688980957
transform 1 0 11408 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0735_
timestamp 1688980957
transform -1 0 11408 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0736_
timestamp 1688980957
transform 1 0 11592 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0737_
timestamp 1688980957
transform -1 0 11132 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0738_
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0739_
timestamp 1688980957
transform 1 0 10948 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0740_
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0741_
timestamp 1688980957
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0742_
timestamp 1688980957
transform -1 0 13984 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0743_
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0744_
timestamp 1688980957
transform -1 0 19044 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0745_
timestamp 1688980957
transform -1 0 18676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0746_
timestamp 1688980957
transform 1 0 17940 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0747_
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0749_
timestamp 1688980957
transform 1 0 17388 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0750_
timestamp 1688980957
transform 1 0 15180 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0751_
timestamp 1688980957
transform 1 0 14720 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 1688980957
transform 1 0 16560 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0753_
timestamp 1688980957
transform -1 0 16560 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0754_
timestamp 1688980957
transform 1 0 10580 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0755_
timestamp 1688980957
transform -1 0 10580 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 1688980957
transform 1 0 12972 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0757_
timestamp 1688980957
transform -1 0 11408 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0758_
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0759_
timestamp 1688980957
transform 1 0 10580 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 1688980957
transform 1 0 10580 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0761_
timestamp 1688980957
transform 1 0 10120 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0762_
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0763_
timestamp 1688980957
transform -1 0 13156 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0764_
timestamp 1688980957
transform -1 0 21252 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0765_
timestamp 1688980957
transform -1 0 19320 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_2  _0766_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19872 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0767_
timestamp 1688980957
transform 1 0 19044 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  _0768_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19964 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0769_
timestamp 1688980957
transform -1 0 20240 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0770_
timestamp 1688980957
transform -1 0 19780 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0771_
timestamp 1688980957
transform 1 0 16836 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0772_
timestamp 1688980957
transform 1 0 19780 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _0773_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12420 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0774_
timestamp 1688980957
transform 1 0 18492 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0775_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0776_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17848 0 1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _0777_
timestamp 1688980957
transform 1 0 17480 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0778_
timestamp 1688980957
transform 1 0 17020 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0779_
timestamp 1688980957
transform 1 0 16468 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0780_
timestamp 1688980957
transform 1 0 17020 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0781_
timestamp 1688980957
transform 1 0 17572 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0782_
timestamp 1688980957
transform 1 0 17296 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0783_
timestamp 1688980957
transform 1 0 14996 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0784_
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0786_
timestamp 1688980957
transform 1 0 16192 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0787_
timestamp 1688980957
transform 1 0 15824 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0788_
timestamp 1688980957
transform 1 0 18584 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0790_
timestamp 1688980957
transform 1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0791_
timestamp 1688980957
transform 1 0 10396 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0792_
timestamp 1688980957
transform 1 0 12236 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1688980957
transform -1 0 11408 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0794_
timestamp 1688980957
transform 1 0 11316 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0795_
timestamp 1688980957
transform 1 0 10396 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0796_
timestamp 1688980957
transform 1 0 11868 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0797_
timestamp 1688980957
transform 1 0 11960 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0798_
timestamp 1688980957
transform 1 0 11684 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0799_
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0800_
timestamp 1688980957
transform 1 0 13248 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0802_
timestamp 1688980957
transform 1 0 9476 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0803_
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0804_
timestamp 1688980957
transform 1 0 11408 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1688980957
transform 1 0 10120 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0806_
timestamp 1688980957
transform 1 0 9844 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0807_
timestamp 1688980957
transform 1 0 14812 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0808_
timestamp 1688980957
transform 1 0 15548 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp 1688980957
transform 1 0 14076 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0810_
timestamp 1688980957
transform -1 0 14352 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0811_
timestamp 1688980957
transform -1 0 16560 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0812_
timestamp 1688980957
transform -1 0 16100 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0813_
timestamp 1688980957
transform -1 0 13984 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp 1688980957
transform 1 0 12144 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0815_
timestamp 1688980957
transform 1 0 11868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0816_
timestamp 1688980957
transform 1 0 7268 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0817_
timestamp 1688980957
transform 1 0 10304 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0818_
timestamp 1688980957
transform -1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0819_
timestamp 1688980957
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1688980957
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0821_
timestamp 1688980957
transform -1 0 9200 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0822_
timestamp 1688980957
transform -1 0 11960 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0823_
timestamp 1688980957
transform 1 0 11224 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1688980957
transform 1 0 13156 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0825_
timestamp 1688980957
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0826_
timestamp 1688980957
transform 1 0 10856 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0827_
timestamp 1688980957
transform -1 0 10580 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0828_
timestamp 1688980957
transform -1 0 10304 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0829_
timestamp 1688980957
transform 1 0 9200 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _0830_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8832 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0831_
timestamp 1688980957
transform 1 0 8832 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0832_
timestamp 1688980957
transform -1 0 9200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _0833_
timestamp 1688980957
transform 1 0 14168 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _0834_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14536 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0835_
timestamp 1688980957
transform 1 0 14904 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0836_
timestamp 1688980957
transform -1 0 13432 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0837_
timestamp 1688980957
transform -1 0 11868 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0838_
timestamp 1688980957
transform -1 0 8372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0839_
timestamp 1688980957
transform -1 0 7636 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_2  _0840_
timestamp 1688980957
transform -1 0 7636 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1688980957
transform -1 0 10396 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0842_
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0843_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0844_
timestamp 1688980957
transform -1 0 7452 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0845_
timestamp 1688980957
transform -1 0 8832 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0846_
timestamp 1688980957
transform 1 0 9844 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0847_
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0848_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11132 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0849_
timestamp 1688980957
transform 1 0 10672 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0850_
timestamp 1688980957
transform -1 0 7268 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0851_
timestamp 1688980957
transform 1 0 10488 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0852_
timestamp 1688980957
transform 1 0 9568 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0853_
timestamp 1688980957
transform 1 0 9844 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0854_
timestamp 1688980957
transform 1 0 10856 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0855_
timestamp 1688980957
transform 1 0 9292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0856_
timestamp 1688980957
transform -1 0 8924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0857_
timestamp 1688980957
transform -1 0 8464 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0858_
timestamp 1688980957
transform -1 0 6624 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0859_
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0860_
timestamp 1688980957
transform 1 0 2668 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0861_
timestamp 1688980957
transform -1 0 4784 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0862_
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0863_
timestamp 1688980957
transform 1 0 7912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0864_
timestamp 1688980957
transform -1 0 7360 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0865_
timestamp 1688980957
transform -1 0 6808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0866_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6256 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0867_
timestamp 1688980957
transform 1 0 5612 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0868_
timestamp 1688980957
transform -1 0 7636 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1688980957
transform 1 0 7544 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0870_
timestamp 1688980957
transform -1 0 7452 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0871_
timestamp 1688980957
transform -1 0 8188 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0872_
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _0873_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6256 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0874_
timestamp 1688980957
transform -1 0 7176 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0875_
timestamp 1688980957
transform -1 0 6808 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0876_
timestamp 1688980957
transform -1 0 6348 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0877_
timestamp 1688980957
transform 1 0 5612 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0878_
timestamp 1688980957
transform -1 0 4140 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0879_
timestamp 1688980957
transform 1 0 5888 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0880_
timestamp 1688980957
transform -1 0 5612 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0881_
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0882_
timestamp 1688980957
transform -1 0 5980 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0883_
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0884_
timestamp 1688980957
transform 1 0 5428 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0885_
timestamp 1688980957
transform 1 0 2392 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0886_
timestamp 1688980957
transform -1 0 17296 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0887_
timestamp 1688980957
transform -1 0 17204 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0888_
timestamp 1688980957
transform -1 0 19136 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0889_
timestamp 1688980957
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0890_
timestamp 1688980957
transform -1 0 18308 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0891_
timestamp 1688980957
transform -1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0892_
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0893_
timestamp 1688980957
transform -1 0 16560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0894_
timestamp 1688980957
transform -1 0 12512 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0895_
timestamp 1688980957
transform 1 0 11960 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0896_
timestamp 1688980957
transform 1 0 13248 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0897_
timestamp 1688980957
transform 1 0 12512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0898_
timestamp 1688980957
transform -1 0 12328 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0899_
timestamp 1688980957
transform 1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0900_
timestamp 1688980957
transform -1 0 11408 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0902_
timestamp 1688980957
transform 1 0 14812 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0903_
timestamp 1688980957
transform -1 0 15180 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0904_
timestamp 1688980957
transform -1 0 19136 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0905_
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0906_
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0907_
timestamp 1688980957
transform 1 0 18584 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0908_
timestamp 1688980957
transform 1 0 15548 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0909_
timestamp 1688980957
transform -1 0 14444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0910_
timestamp 1688980957
transform 1 0 15364 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0911_
timestamp 1688980957
transform 1 0 14996 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0912_
timestamp 1688980957
transform -1 0 10488 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0913_
timestamp 1688980957
transform 1 0 10120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0914_
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0915_
timestamp 1688980957
transform 1 0 8280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0916_
timestamp 1688980957
transform 1 0 7452 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0917_
timestamp 1688980957
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0918_
timestamp 1688980957
transform 1 0 10120 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0919_
timestamp 1688980957
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0920_
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0921_
timestamp 1688980957
transform 1 0 13248 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0922_
timestamp 1688980957
transform -1 0 18216 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0923_
timestamp 1688980957
transform -1 0 17848 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0924_
timestamp 1688980957
transform 1 0 15916 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0925_
timestamp 1688980957
transform 1 0 15548 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0926_
timestamp 1688980957
transform 1 0 15640 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0927_
timestamp 1688980957
transform -1 0 14996 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0928_
timestamp 1688980957
transform 1 0 15916 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0929_
timestamp 1688980957
transform -1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0930_
timestamp 1688980957
transform 1 0 14260 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0931_
timestamp 1688980957
transform -1 0 13984 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0932_
timestamp 1688980957
transform 1 0 9200 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0933_
timestamp 1688980957
transform 1 0 8832 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0934_
timestamp 1688980957
transform 1 0 9292 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0935_
timestamp 1688980957
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0936_
timestamp 1688980957
transform 1 0 9108 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0937_
timestamp 1688980957
transform 1 0 9108 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0938_
timestamp 1688980957
transform 1 0 8740 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0939_
timestamp 1688980957
transform -1 0 8832 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0940_
timestamp 1688980957
transform 1 0 12696 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0941_
timestamp 1688980957
transform -1 0 12144 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0942_
timestamp 1688980957
transform -1 0 20884 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0943_
timestamp 1688980957
transform -1 0 21528 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0944_
timestamp 1688980957
transform 1 0 22816 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0945_
timestamp 1688980957
transform -1 0 21712 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0946_
timestamp 1688980957
transform -1 0 23368 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0947_
timestamp 1688980957
transform -1 0 23460 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0948_
timestamp 1688980957
transform 1 0 19964 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0949_
timestamp 1688980957
transform -1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0950_
timestamp 1688980957
transform -1 0 21712 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0951_
timestamp 1688980957
transform 1 0 23460 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0952_
timestamp 1688980957
transform 1 0 22448 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0953_
timestamp 1688980957
transform -1 0 22264 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0954_
timestamp 1688980957
transform 1 0 20792 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0955_
timestamp 1688980957
transform -1 0 19136 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _0956_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25300 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0957_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19872 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0958_
timestamp 1688980957
transform -1 0 22908 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0959_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22172 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0960_
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0961_
timestamp 1688980957
transform 1 0 20148 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0962_
timestamp 1688980957
transform 1 0 18400 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _0963_
timestamp 1688980957
transform 1 0 22356 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0964_
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0965_
timestamp 1688980957
transform 1 0 19872 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0966_
timestamp 1688980957
transform 1 0 19412 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0967_
timestamp 1688980957
transform -1 0 23736 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0968_
timestamp 1688980957
transform 1 0 20424 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0969_
timestamp 1688980957
transform 1 0 21804 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0970_
timestamp 1688980957
transform 1 0 20424 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0971_
timestamp 1688980957
transform 1 0 14444 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0972_
timestamp 1688980957
transform 1 0 18492 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0973_
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0974_
timestamp 1688980957
transform 1 0 4416 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0975_
timestamp 1688980957
transform 1 0 4968 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0976_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2668 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0977_
timestamp 1688980957
transform -1 0 8280 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0978_
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0979_
timestamp 1688980957
transform 1 0 5612 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0980_
timestamp 1688980957
transform -1 0 23644 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0981_
timestamp 1688980957
transform -1 0 23644 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0982_
timestamp 1688980957
transform -1 0 24196 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0983_
timestamp 1688980957
transform -1 0 23644 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0984_
timestamp 1688980957
transform 1 0 21896 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0985_
timestamp 1688980957
transform 1 0 19688 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0986_
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0987_
timestamp 1688980957
transform 1 0 7728 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0988_
timestamp 1688980957
transform 1 0 5152 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0989_
timestamp 1688980957
transform 1 0 13064 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0990_
timestamp 1688980957
transform 1 0 6992 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0991_
timestamp 1688980957
transform 1 0 6256 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0992_
timestamp 1688980957
transform 1 0 5520 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0993_
timestamp 1688980957
transform 1 0 6532 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0994_
timestamp 1688980957
transform 1 0 6992 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0995_
timestamp 1688980957
transform -1 0 5704 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0996_
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0997_
timestamp 1688980957
transform 1 0 4048 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0998_
timestamp 1688980957
transform 1 0 2760 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0999_
timestamp 1688980957
transform 1 0 1564 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1000_
timestamp 1688980957
transform 1 0 1564 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1001_
timestamp 1688980957
transform 1 0 1564 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1002_
timestamp 1688980957
transform 1 0 1564 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1003_
timestamp 1688980957
transform 1 0 1564 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1004_
timestamp 1688980957
transform 1 0 1564 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1005_
timestamp 1688980957
transform 1 0 2760 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1006_
timestamp 1688980957
transform -1 0 25760 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1007_
timestamp 1688980957
transform 1 0 23460 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1008_
timestamp 1688980957
transform 1 0 23184 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1009_
timestamp 1688980957
transform 1 0 22448 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1010_
timestamp 1688980957
transform -1 0 25852 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1011_
timestamp 1688980957
transform 1 0 20516 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1012_
timestamp 1688980957
transform -1 0 24288 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1013_
timestamp 1688980957
transform 1 0 20424 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1014_
timestamp 1688980957
transform -1 0 25852 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1015_
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1016_
timestamp 1688980957
transform -1 0 25484 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1017_
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1018_
timestamp 1688980957
transform -1 0 22172 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1019_
timestamp 1688980957
transform -1 0 20148 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1020_
timestamp 1688980957
transform -1 0 20056 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1021_
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1022_
timestamp 1688980957
transform 1 0 17112 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1023_
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1024_
timestamp 1688980957
transform 1 0 13984 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1025_
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1026_
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1027_
timestamp 1688980957
transform 1 0 8280 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1028_
timestamp 1688980957
transform 1 0 8464 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1029_
timestamp 1688980957
transform 1 0 12144 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1030_
timestamp 1688980957
transform 1 0 16928 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1031_
timestamp 1688980957
transform -1 0 19872 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1032_
timestamp 1688980957
transform 1 0 14996 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1033_
timestamp 1688980957
transform 1 0 16468 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1034_
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1035_
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1036_
timestamp 1688980957
transform 1 0 10672 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1037_
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1038_
timestamp 1688980957
transform 1 0 13156 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1039_
timestamp 1688980957
transform 1 0 16100 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1040_
timestamp 1688980957
transform 1 0 17112 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1041_
timestamp 1688980957
transform 1 0 14536 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1042_
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1043_
timestamp 1688980957
transform 1 0 10764 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1044_
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1045_
timestamp 1688980957
transform 1 0 10212 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1046_
timestamp 1688980957
transform 1 0 9568 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1047_
timestamp 1688980957
transform 1 0 12972 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1048_
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1049_
timestamp 1688980957
transform 1 0 16928 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1050_
timestamp 1688980957
transform 1 0 16008 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1051_
timestamp 1688980957
transform 1 0 15640 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1052_
timestamp 1688980957
transform 1 0 10948 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1053_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1054_
timestamp 1688980957
transform -1 0 9568 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1055_
timestamp 1688980957
transform 1 0 9568 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1056_
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1057_
timestamp 1688980957
transform 1 0 11592 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1058_
timestamp 1688980957
transform 1 0 8004 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1059_
timestamp 1688980957
transform 1 0 10488 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1060_
timestamp 1688980957
transform 1 0 11592 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1061_
timestamp 1688980957
transform 1 0 1748 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1062_
timestamp 1688980957
transform -1 0 4876 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1063_
timestamp 1688980957
transform -1 0 3588 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1064_
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1065_
timestamp 1688980957
transform 1 0 22264 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1066_
timestamp 1688980957
transform 1 0 23644 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1067_
timestamp 1688980957
transform 1 0 23828 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1068_
timestamp 1688980957
transform -1 0 22540 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1069_
timestamp 1688980957
transform 1 0 17020 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1070_
timestamp 1688980957
transform 1 0 18584 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1071_
timestamp 1688980957
transform -1 0 18952 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1072_
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1073_
timestamp 1688980957
transform 1 0 10856 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1074_
timestamp 1688980957
transform 1 0 12052 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1075_
timestamp 1688980957
transform 1 0 10212 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1076_
timestamp 1688980957
transform 1 0 10580 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1077_
timestamp 1688980957
transform -1 0 16008 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1078_
timestamp 1688980957
transform -1 0 19320 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1079_
timestamp 1688980957
transform 1 0 18308 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1080_
timestamp 1688980957
transform 1 0 14444 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1081_
timestamp 1688980957
transform 1 0 14352 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1082_
timestamp 1688980957
transform -1 0 10212 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1083_
timestamp 1688980957
transform 1 0 7636 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1084_
timestamp 1688980957
transform 1 0 5612 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1085_
timestamp 1688980957
transform 1 0 9016 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1086_
timestamp 1688980957
transform 1 0 12696 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1087_
timestamp 1688980957
transform 1 0 14720 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1088_
timestamp 1688980957
transform 1 0 14720 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1089_
timestamp 1688980957
transform 1 0 13340 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1090_
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1091_
timestamp 1688980957
transform 1 0 8372 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1092_
timestamp 1688980957
transform 1 0 8372 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1093_
timestamp 1688980957
transform 1 0 8188 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1094_
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1095_
timestamp 1688980957
transform 1 0 11868 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1096_
timestamp 1688980957
transform -1 0 20332 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1097_
timestamp 1688980957
transform -1 0 21988 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1098_
timestamp 1688980957
transform 1 0 21068 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1099_
timestamp 1688980957
transform 1 0 21712 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1100_
timestamp 1688980957
transform -1 0 24288 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1101_
timestamp 1688980957
transform 1 0 19044 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1102_
timestamp 1688980957
transform -1 0 21620 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1103_
timestamp 1688980957
transform 1 0 22264 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1104_
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15364 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1688980957
transform -1 0 5612 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1688980957
transform -1 0 10856 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1688980957
transform 1 0 10396 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1688980957
transform -1 0 9936 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1688980957
transform 1 0 12512 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1688980957
transform 1 0 12512 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1688980957
transform -1 0 18216 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1688980957
transform 1 0 17296 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1688980957
transform 1 0 22908 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1688980957
transform 1 0 17572 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1688980957
transform -1 0 20240 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1688980957
transform -1 0 22908 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1688980957
transform -1 0 22816 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout29
timestamp 1688980957
transform -1 0 3312 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout30
timestamp 1688980957
transform 1 0 10304 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout31
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout32
timestamp 1688980957
transform 1 0 20240 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout33
timestamp 1688980957
transform 1 0 17848 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout34
timestamp 1688980957
transform 1 0 14352 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout35
timestamp 1688980957
transform -1 0 21160 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout36 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6808 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_37
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49
timestamp 1688980957
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1688980957
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_69 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_79
timestamp 1688980957
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_163
timestamp 1688980957
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1688980957
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_197 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_205
timestamp 1688980957
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_259
timestamp 1688980957
transform 1 0 24932 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_267
timestamp 1688980957
transform 1 0 25668 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_62
timestamp 1688980957
transform 1 0 6808 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_74
timestamp 1688980957
transform 1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_99
timestamp 1688980957
transform 1 0 10212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_122
timestamp 1688980957
transform 1 0 12328 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_127
timestamp 1688980957
transform 1 0 12788 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_139
timestamp 1688980957
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_143
timestamp 1688980957
transform 1 0 14260 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_164
timestamp 1688980957
transform 1 0 16192 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_173
timestamp 1688980957
transform 1 0 17020 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_194
timestamp 1688980957
transform 1 0 18952 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_206
timestamp 1688980957
transform 1 0 20056 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_218
timestamp 1688980957
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_269
timestamp 1688980957
transform 1 0 25852 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_81
timestamp 1688980957
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_94
timestamp 1688980957
transform 1 0 9752 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_98
timestamp 1688980957
transform 1 0 10120 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_188
timestamp 1688980957
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_201
timestamp 1688980957
transform 1 0 19596 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_222
timestamp 1688980957
transform 1 0 21528 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_101
timestamp 1688980957
transform 1 0 10396 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_141
timestamp 1688980957
transform 1 0 14076 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_154
timestamp 1688980957
transform 1 0 15272 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_164
timestamp 1688980957
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_187
timestamp 1688980957
transform 1 0 18308 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_199
timestamp 1688980957
transform 1 0 19412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_211
timestamp 1688980957
transform 1 0 20516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_245
timestamp 1688980957
transform 1 0 23644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_257
timestamp 1688980957
transform 1 0 24748 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_269
timestamp 1688980957
transform 1 0 25852 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_9
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_21
timestamp 1688980957
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_49
timestamp 1688980957
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_56
timestamp 1688980957
transform 1 0 6256 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_62
timestamp 1688980957
transform 1 0 6808 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_66
timestamp 1688980957
transform 1 0 7176 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_78
timestamp 1688980957
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_102
timestamp 1688980957
transform 1 0 10488 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_123
timestamp 1688980957
transform 1 0 12420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp 1688980957
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_166
timestamp 1688980957
transform 1 0 16376 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_174
timestamp 1688980957
transform 1 0 17112 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_186
timestamp 1688980957
transform 1 0 18216 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_192
timestamp 1688980957
transform 1 0 18768 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_71
timestamp 1688980957
transform 1 0 7636 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_75
timestamp 1688980957
transform 1 0 8004 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_79
timestamp 1688980957
transform 1 0 8372 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_83
timestamp 1688980957
transform 1 0 8740 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_90
timestamp 1688980957
transform 1 0 9384 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_94
timestamp 1688980957
transform 1 0 9752 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_106
timestamp 1688980957
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_135
timestamp 1688980957
transform 1 0 13524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_147
timestamp 1688980957
transform 1 0 14628 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_159
timestamp 1688980957
transform 1 0 15732 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_164
timestamp 1688980957
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_178
timestamp 1688980957
transform 1 0 17480 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_189
timestamp 1688980957
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_211
timestamp 1688980957
transform 1 0 20516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_233
timestamp 1688980957
transform 1 0 22540 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_244
timestamp 1688980957
transform 1 0 23552 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_256
timestamp 1688980957
transform 1 0 24656 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_268
timestamp 1688980957
transform 1 0 25760 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_37
timestamp 1688980957
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_62
timestamp 1688980957
transform 1 0 6808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_71
timestamp 1688980957
transform 1 0 7636 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_90
timestamp 1688980957
transform 1 0 9384 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_107
timestamp 1688980957
transform 1 0 10948 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_111
timestamp 1688980957
transform 1 0 11316 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_117
timestamp 1688980957
transform 1 0 11868 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_125
timestamp 1688980957
transform 1 0 12604 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_134
timestamp 1688980957
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_163
timestamp 1688980957
transform 1 0 16100 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_175
timestamp 1688980957
transform 1 0 17204 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_206
timestamp 1688980957
transform 1 0 20056 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_239
timestamp 1688980957
transform 1 0 23092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_23
timestamp 1688980957
transform 1 0 3220 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_35
timestamp 1688980957
transform 1 0 4324 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_64
timestamp 1688980957
transform 1 0 6992 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_83
timestamp 1688980957
transform 1 0 8740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_106
timestamp 1688980957
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_124
timestamp 1688980957
transform 1 0 12512 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_130
timestamp 1688980957
transform 1 0 13064 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_139
timestamp 1688980957
transform 1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_158
timestamp 1688980957
transform 1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 1688980957
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_185
timestamp 1688980957
transform 1 0 18124 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_208
timestamp 1688980957
transform 1 0 20240 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_220
timestamp 1688980957
transform 1 0 21344 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_265
timestamp 1688980957
transform 1 0 25484 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_11
timestamp 1688980957
transform 1 0 2116 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_18
timestamp 1688980957
transform 1 0 2760 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_49
timestamp 1688980957
transform 1 0 5612 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_58
timestamp 1688980957
transform 1 0 6440 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_96
timestamp 1688980957
transform 1 0 9936 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_104
timestamp 1688980957
transform 1 0 10672 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_126
timestamp 1688980957
transform 1 0 12696 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_131
timestamp 1688980957
transform 1 0 13156 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_174
timestamp 1688980957
transform 1 0 17112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_180
timestamp 1688980957
transform 1 0 17664 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_188
timestamp 1688980957
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_193
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_217
timestamp 1688980957
transform 1 0 21068 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_239
timestamp 1688980957
transform 1 0 23092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_258
timestamp 1688980957
transform 1 0 24840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_269
timestamp 1688980957
transform 1 0 25852 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_85
timestamp 1688980957
transform 1 0 8924 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_92
timestamp 1688980957
transform 1 0 9568 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_104
timestamp 1688980957
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_121
timestamp 1688980957
transform 1 0 12236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_140
timestamp 1688980957
transform 1 0 13984 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_155
timestamp 1688980957
transform 1 0 15364 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_163
timestamp 1688980957
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_177
timestamp 1688980957
transform 1 0 17388 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_198
timestamp 1688980957
transform 1 0 19320 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_210
timestamp 1688980957
transform 1 0 20424 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_219
timestamp 1688980957
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_265
timestamp 1688980957
transform 1 0 25484 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_22
timestamp 1688980957
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_32
timestamp 1688980957
transform 1 0 4048 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_78
timestamp 1688980957
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_105
timestamp 1688980957
transform 1 0 10764 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_132
timestamp 1688980957
transform 1 0 13248 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_148
timestamp 1688980957
transform 1 0 14720 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_170
timestamp 1688980957
transform 1 0 16744 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_200
timestamp 1688980957
transform 1 0 19504 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_6
timestamp 1688980957
transform 1 0 1656 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_44
timestamp 1688980957
transform 1 0 5152 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_82
timestamp 1688980957
transform 1 0 8648 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_94
timestamp 1688980957
transform 1 0 9752 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_107
timestamp 1688980957
transform 1 0 10948 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_134
timestamp 1688980957
transform 1 0 13432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_209
timestamp 1688980957
transform 1 0 20332 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_219
timestamp 1688980957
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_233
timestamp 1688980957
transform 1 0 22540 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_267
timestamp 1688980957
transform 1 0 25668 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1688980957
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_42
timestamp 1688980957
transform 1 0 4968 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_51
timestamp 1688980957
transform 1 0 5796 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_59
timestamp 1688980957
transform 1 0 6532 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_63
timestamp 1688980957
transform 1 0 6900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_79
timestamp 1688980957
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_100
timestamp 1688980957
transform 1 0 10304 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_108
timestamp 1688980957
transform 1 0 11040 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_119
timestamp 1688980957
transform 1 0 12052 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_131
timestamp 1688980957
transform 1 0 13156 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_135
timestamp 1688980957
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_162
timestamp 1688980957
transform 1 0 16008 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_166
timestamp 1688980957
transform 1 0 16376 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_205
timestamp 1688980957
transform 1 0 19964 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_227
timestamp 1688980957
transform 1 0 21988 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_250
timestamp 1688980957
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_9
timestamp 1688980957
transform 1 0 1932 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_14
timestamp 1688980957
transform 1 0 2392 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_40
timestamp 1688980957
transform 1 0 4784 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_52
timestamp 1688980957
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_62
timestamp 1688980957
transform 1 0 6808 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_74
timestamp 1688980957
transform 1 0 7912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_78
timestamp 1688980957
transform 1 0 8280 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_88
timestamp 1688980957
transform 1 0 9200 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_92
timestamp 1688980957
transform 1 0 9568 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_97
timestamp 1688980957
transform 1 0 10028 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_158
timestamp 1688980957
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1688980957
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_189
timestamp 1688980957
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 1688980957
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_233
timestamp 1688980957
transform 1 0 22540 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_241
timestamp 1688980957
transform 1 0 23276 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_263
timestamp 1688980957
transform 1 0 25300 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_270
timestamp 1688980957
transform 1 0 25944 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_11
timestamp 1688980957
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_20
timestamp 1688980957
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_42
timestamp 1688980957
transform 1 0 4968 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_66
timestamp 1688980957
transform 1 0 7176 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_106
timestamp 1688980957
transform 1 0 10856 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_118
timestamp 1688980957
transform 1 0 11960 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_130
timestamp 1688980957
transform 1 0 13064 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1688980957
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_157
timestamp 1688980957
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_178
timestamp 1688980957
transform 1 0 17480 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_190
timestamp 1688980957
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_203
timestamp 1688980957
transform 1 0 19780 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_224
timestamp 1688980957
transform 1 0 21712 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_230
timestamp 1688980957
transform 1 0 22264 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_270
timestamp 1688980957
transform 1 0 25944 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_33
timestamp 1688980957
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_45
timestamp 1688980957
transform 1 0 5244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1688980957
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_71
timestamp 1688980957
transform 1 0 7636 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_88
timestamp 1688980957
transform 1 0 9200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1688980957
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_166
timestamp 1688980957
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_187
timestamp 1688980957
transform 1 0 18308 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_222
timestamp 1688980957
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_228
timestamp 1688980957
transform 1 0 22080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_252
timestamp 1688980957
transform 1 0 24288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_270
timestamp 1688980957
transform 1 0 25944 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_19
timestamp 1688980957
transform 1 0 2852 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_63
timestamp 1688980957
transform 1 0 6900 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_71
timestamp 1688980957
transform 1 0 7636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_80
timestamp 1688980957
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_93
timestamp 1688980957
transform 1 0 9660 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_113
timestamp 1688980957
transform 1 0 11500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_137
timestamp 1688980957
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_149
timestamp 1688980957
transform 1 0 14812 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_161
timestamp 1688980957
transform 1 0 15916 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_184
timestamp 1688980957
transform 1 0 18032 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_248
timestamp 1688980957
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_268
timestamp 1688980957
transform 1 0 25760 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_20
timestamp 1688980957
transform 1 0 2944 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_62
timestamp 1688980957
transform 1 0 6808 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_74
timestamp 1688980957
transform 1 0 7912 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_86
timestamp 1688980957
transform 1 0 9016 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_94
timestamp 1688980957
transform 1 0 9752 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_134
timestamp 1688980957
transform 1 0 13432 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_140
timestamp 1688980957
transform 1 0 13984 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_147
timestamp 1688980957
transform 1 0 14628 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_162
timestamp 1688980957
transform 1 0 16008 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_187
timestamp 1688980957
transform 1 0 18308 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_222
timestamp 1688980957
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_231
timestamp 1688980957
transform 1 0 22356 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_239
timestamp 1688980957
transform 1 0 23092 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_263
timestamp 1688980957
transform 1 0 25300 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_6
timestamp 1688980957
transform 1 0 1656 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_49
timestamp 1688980957
transform 1 0 5612 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_67
timestamp 1688980957
transform 1 0 7268 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_79
timestamp 1688980957
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_93
timestamp 1688980957
transform 1 0 9660 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_101
timestamp 1688980957
transform 1 0 10396 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_160
timestamp 1688980957
transform 1 0 15824 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_172
timestamp 1688980957
transform 1 0 16928 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_188
timestamp 1688980957
transform 1 0 18400 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_209
timestamp 1688980957
transform 1 0 20332 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_230
timestamp 1688980957
transform 1 0 22264 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_242
timestamp 1688980957
transform 1 0 23368 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1688980957
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_265
timestamp 1688980957
transform 1 0 25484 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_23
timestamp 1688980957
transform 1 0 3220 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_31
timestamp 1688980957
transform 1 0 3956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_66
timestamp 1688980957
transform 1 0 7176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_96
timestamp 1688980957
transform 1 0 9936 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_129
timestamp 1688980957
transform 1 0 12972 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_200
timestamp 1688980957
transform 1 0 19504 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_208
timestamp 1688980957
transform 1 0 20240 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_220
timestamp 1688980957
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_231
timestamp 1688980957
transform 1 0 22356 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_240
timestamp 1688980957
transform 1 0 23184 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_263
timestamp 1688980957
transform 1 0 25300 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_23
timestamp 1688980957
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_50
timestamp 1688980957
transform 1 0 5704 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_57
timestamp 1688980957
transform 1 0 6348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_91
timestamp 1688980957
transform 1 0 9476 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_103
timestamp 1688980957
transform 1 0 10580 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_115
timestamp 1688980957
transform 1 0 11684 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_126
timestamp 1688980957
transform 1 0 12696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_130
timestamp 1688980957
transform 1 0 13064 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_134
timestamp 1688980957
transform 1 0 13432 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_158
timestamp 1688980957
transform 1 0 15640 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_191
timestamp 1688980957
transform 1 0 18676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_221
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_266
timestamp 1688980957
transform 1 0 25576 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_60
timestamp 1688980957
transform 1 0 6624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_122
timestamp 1688980957
transform 1 0 12328 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_134
timestamp 1688980957
transform 1 0 13432 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_140
timestamp 1688980957
transform 1 0 13984 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_153
timestamp 1688980957
transform 1 0 15180 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_161
timestamp 1688980957
transform 1 0 15916 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_178
timestamp 1688980957
transform 1 0 17480 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_207
timestamp 1688980957
transform 1 0 20148 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_215
timestamp 1688980957
transform 1 0 20884 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_243
timestamp 1688980957
transform 1 0 23460 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_268
timestamp 1688980957
transform 1 0 25760 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_64
timestamp 1688980957
transform 1 0 6992 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_72
timestamp 1688980957
transform 1 0 7728 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_80
timestamp 1688980957
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_94
timestamp 1688980957
transform 1 0 9752 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_127
timestamp 1688980957
transform 1 0 12788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_161
timestamp 1688980957
transform 1 0 15916 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_173
timestamp 1688980957
transform 1 0 17020 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_185
timestamp 1688980957
transform 1 0 18124 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1688980957
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_208
timestamp 1688980957
transform 1 0 20240 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 1688980957
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_268
timestamp 1688980957
transform 1 0 25760 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_37
timestamp 1688980957
transform 1 0 4508 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_49
timestamp 1688980957
transform 1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_61
timestamp 1688980957
transform 1 0 6716 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_71
timestamp 1688980957
transform 1 0 7636 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_85
timestamp 1688980957
transform 1 0 8924 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_97
timestamp 1688980957
transform 1 0 10028 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_133
timestamp 1688980957
transform 1 0 13340 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_155
timestamp 1688980957
transform 1 0 15364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1688980957
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_206
timestamp 1688980957
transform 1 0 20056 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_214
timestamp 1688980957
transform 1 0 20792 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_269
timestamp 1688980957
transform 1 0 25852 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_38
timestamp 1688980957
transform 1 0 4600 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_114
timestamp 1688980957
transform 1 0 11592 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_127
timestamp 1688980957
transform 1 0 12788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_144
timestamp 1688980957
transform 1 0 14352 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_156
timestamp 1688980957
transform 1 0 15456 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_168
timestamp 1688980957
transform 1 0 16560 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_246
timestamp 1688980957
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_261
timestamp 1688980957
transform 1 0 25116 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_269
timestamp 1688980957
transform 1 0 25852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_9
timestamp 1688980957
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_25
timestamp 1688980957
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_37
timestamp 1688980957
transform 1 0 4508 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_50
timestamp 1688980957
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_78
timestamp 1688980957
transform 1 0 8280 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_107
timestamp 1688980957
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_137
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_145
timestamp 1688980957
transform 1 0 14444 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_166
timestamp 1688980957
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_177
timestamp 1688980957
transform 1 0 17388 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_211
timestamp 1688980957
transform 1 0 20516 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_248
timestamp 1688980957
transform 1 0 23920 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_269
timestamp 1688980957
transform 1 0 25852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_9
timestamp 1688980957
transform 1 0 1932 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_14
timestamp 1688980957
transform 1 0 2392 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1688980957
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_77
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1688980957
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 1688980957
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1688980957
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_265
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_28
timestamp 1688980957
transform 1 0 3680 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_32
timestamp 1688980957
transform 1 0 4048 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_66
timestamp 1688980957
transform 1 0 7176 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_78
timestamp 1688980957
transform 1 0 8280 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_87
timestamp 1688980957
transform 1 0 9108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_98
timestamp 1688980957
transform 1 0 10120 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_133
timestamp 1688980957
transform 1 0 13340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_141
timestamp 1688980957
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_152
timestamp 1688980957
transform 1 0 15088 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_162
timestamp 1688980957
transform 1 0 16008 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_177
timestamp 1688980957
transform 1 0 17388 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_197
timestamp 1688980957
transform 1 0 19228 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_208
timestamp 1688980957
transform 1 0 20240 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_237
timestamp 1688980957
transform 1 0 22908 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1688980957
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_261
timestamp 1688980957
transform 1 0 25116 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_267
timestamp 1688980957
transform 1 0 25668 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_63
timestamp 1688980957
transform 1 0 6900 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_79
timestamp 1688980957
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_107
timestamp 1688980957
transform 1 0 10948 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_121
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_133
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_170
timestamp 1688980957
transform 1 0 16744 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_193
timestamp 1688980957
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_221
timestamp 1688980957
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_250
timestamp 1688980957
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_265
timestamp 1688980957
transform 1 0 25484 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_11
timestamp 1688980957
transform 1 0 2116 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_34
timestamp 1688980957
transform 1 0 4232 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_49
timestamp 1688980957
transform 1 0 5612 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1688980957
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_64
timestamp 1688980957
transform 1 0 6992 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_108
timestamp 1688980957
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_129
timestamp 1688980957
transform 1 0 12972 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_153
timestamp 1688980957
transform 1 0 15180 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_162
timestamp 1688980957
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_180
timestamp 1688980957
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_212
timestamp 1688980957
transform 1 0 20608 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_246
timestamp 1688980957
transform 1 0 23736 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_258
timestamp 1688980957
transform 1 0 24840 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_270
timestamp 1688980957
transform 1 0 25944 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_54
timestamp 1688980957
transform 1 0 6072 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_66
timestamp 1688980957
transform 1 0 7176 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_78
timestamp 1688980957
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_98
timestamp 1688980957
transform 1 0 10120 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_108
timestamp 1688980957
transform 1 0 11040 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_116
timestamp 1688980957
transform 1 0 11776 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_125
timestamp 1688980957
transform 1 0 12604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_137
timestamp 1688980957
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_147
timestamp 1688980957
transform 1 0 14628 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1688980957
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_206
timestamp 1688980957
transform 1 0 20056 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_230
timestamp 1688980957
transform 1 0 22264 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_256
timestamp 1688980957
transform 1 0 24656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_268
timestamp 1688980957
transform 1 0 25760 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_37
timestamp 1688980957
transform 1 0 4508 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_60
timestamp 1688980957
transform 1 0 6624 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_64
timestamp 1688980957
transform 1 0 6992 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_73
timestamp 1688980957
transform 1 0 7820 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_107
timestamp 1688980957
transform 1 0 10948 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_133
timestamp 1688980957
transform 1 0 13340 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_145
timestamp 1688980957
transform 1 0 14444 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_194
timestamp 1688980957
transform 1 0 18952 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_261
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_269
timestamp 1688980957
transform 1 0 25852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_33
timestamp 1688980957
transform 1 0 4140 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_76
timestamp 1688980957
transform 1 0 8096 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_80
timestamp 1688980957
transform 1 0 8464 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_105
timestamp 1688980957
transform 1 0 10764 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 1688980957
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_149
timestamp 1688980957
transform 1 0 14812 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_161
timestamp 1688980957
transform 1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_173
timestamp 1688980957
transform 1 0 17020 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_185
timestamp 1688980957
transform 1 0 18124 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_209
timestamp 1688980957
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_216
timestamp 1688980957
transform 1 0 20976 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_224
timestamp 1688980957
transform 1 0 21712 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_250
timestamp 1688980957
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_265
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_17
timestamp 1688980957
transform 1 0 2668 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_28
timestamp 1688980957
transform 1 0 3680 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_40
timestamp 1688980957
transform 1 0 4784 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_48
timestamp 1688980957
transform 1 0 5520 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_65
timestamp 1688980957
transform 1 0 7084 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_77
timestamp 1688980957
transform 1 0 8188 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_85
timestamp 1688980957
transform 1 0 8924 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_99
timestamp 1688980957
transform 1 0 10212 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_108
timestamp 1688980957
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_123
timestamp 1688980957
transform 1 0 12420 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_129
timestamp 1688980957
transform 1 0 12972 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_150
timestamp 1688980957
transform 1 0 14904 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_158
timestamp 1688980957
transform 1 0 15640 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_198
timestamp 1688980957
transform 1 0 19320 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_210
timestamp 1688980957
transform 1 0 20424 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_218
timestamp 1688980957
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_252
timestamp 1688980957
transform 1 0 24288 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_263
timestamp 1688980957
transform 1 0 25300 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_21
timestamp 1688980957
transform 1 0 3036 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_25
timestamp 1688980957
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_38
timestamp 1688980957
transform 1 0 4600 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_46
timestamp 1688980957
transform 1 0 5336 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_56
timestamp 1688980957
transform 1 0 6256 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_74
timestamp 1688980957
transform 1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_82
timestamp 1688980957
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_96
timestamp 1688980957
transform 1 0 9936 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_108
timestamp 1688980957
transform 1 0 11040 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_120
timestamp 1688980957
transform 1 0 12144 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_135
timestamp 1688980957
transform 1 0 13524 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_161
timestamp 1688980957
transform 1 0 15916 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1688980957
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_217
timestamp 1688980957
transform 1 0 21068 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_244
timestamp 1688980957
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_265
timestamp 1688980957
transform 1 0 25484 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_9
timestamp 1688980957
transform 1 0 1932 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_17
timestamp 1688980957
transform 1 0 2668 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_41
timestamp 1688980957
transform 1 0 4876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_53
timestamp 1688980957
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_76
timestamp 1688980957
transform 1 0 8096 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_106
timestamp 1688980957
transform 1 0 10856 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_122
timestamp 1688980957
transform 1 0 12328 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_189
timestamp 1688980957
transform 1 0 18492 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_197
timestamp 1688980957
transform 1 0 19228 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_219
timestamp 1688980957
transform 1 0 21252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1688980957
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_234
timestamp 1688980957
transform 1 0 22632 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_248
timestamp 1688980957
transform 1 0 23920 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_260
timestamp 1688980957
transform 1 0 25024 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_266
timestamp 1688980957
transform 1 0 25576 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_47
timestamp 1688980957
transform 1 0 5428 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_68
timestamp 1688980957
transform 1 0 7360 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_80
timestamp 1688980957
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_135
timestamp 1688980957
transform 1 0 13524 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_180
timestamp 1688980957
transform 1 0 17664 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 1688980957
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_214
timestamp 1688980957
transform 1 0 20792 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_241
timestamp 1688980957
transform 1 0 23276 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_249
timestamp 1688980957
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_265
timestamp 1688980957
transform 1 0 25484 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_38
timestamp 1688980957
transform 1 0 4600 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_53
timestamp 1688980957
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_68
timestamp 1688980957
transform 1 0 7360 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_76
timestamp 1688980957
transform 1 0 8096 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_105
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_110
timestamp 1688980957
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_130
timestamp 1688980957
transform 1 0 13064 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_142
timestamp 1688980957
transform 1 0 14168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_152
timestamp 1688980957
transform 1 0 15088 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_164
timestamp 1688980957
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_193
timestamp 1688980957
transform 1 0 18860 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_250
timestamp 1688980957
transform 1 0 24104 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_262
timestamp 1688980957
transform 1 0 25208 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_270
timestamp 1688980957
transform 1 0 25944 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_55
timestamp 1688980957
transform 1 0 6164 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_96
timestamp 1688980957
transform 1 0 9936 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_119
timestamp 1688980957
transform 1 0 12052 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_131
timestamp 1688980957
transform 1 0 13156 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_153
timestamp 1688980957
transform 1 0 15180 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_161
timestamp 1688980957
transform 1 0 15916 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_169
timestamp 1688980957
transform 1 0 16652 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_175
timestamp 1688980957
transform 1 0 17204 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_185
timestamp 1688980957
transform 1 0 18124 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_189
timestamp 1688980957
transform 1 0 18492 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_231
timestamp 1688980957
transform 1 0 22356 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_242
timestamp 1688980957
transform 1 0 23368 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_265
timestamp 1688980957
transform 1 0 25484 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_35
timestamp 1688980957
transform 1 0 4324 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_90
timestamp 1688980957
transform 1 0 9384 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_102
timestamp 1688980957
transform 1 0 10488 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_106
timestamp 1688980957
transform 1 0 10856 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_117
timestamp 1688980957
transform 1 0 11868 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_126
timestamp 1688980957
transform 1 0 12696 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_151
timestamp 1688980957
transform 1 0 14996 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1688980957
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_252
timestamp 1688980957
transform 1 0 24288 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_264
timestamp 1688980957
transform 1 0 25392 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_270
timestamp 1688980957
transform 1 0 25944 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_52
timestamp 1688980957
transform 1 0 5888 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_64
timestamp 1688980957
transform 1 0 6992 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_78
timestamp 1688980957
transform 1 0 8280 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_101
timestamp 1688980957
transform 1 0 10396 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_162
timestamp 1688980957
transform 1 0 16008 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_205
timestamp 1688980957
transform 1 0 19964 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_246
timestamp 1688980957
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_35
timestamp 1688980957
transform 1 0 4324 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_71
timestamp 1688980957
transform 1 0 7636 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_122
timestamp 1688980957
transform 1 0 12328 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_128
timestamp 1688980957
transform 1 0 12880 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_165
timestamp 1688980957
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_192
timestamp 1688980957
transform 1 0 18768 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_251
timestamp 1688980957
transform 1 0 24196 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_263
timestamp 1688980957
transform 1 0 25300 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_6
timestamp 1688980957
transform 1 0 1656 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_18
timestamp 1688980957
transform 1 0 2760 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_26
timestamp 1688980957
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_74
timestamp 1688980957
transform 1 0 7912 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_80
timestamp 1688980957
transform 1 0 8464 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_137
timestamp 1688980957
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_171
timestamp 1688980957
transform 1 0 16836 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 1688980957
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_261
timestamp 1688980957
transform 1 0 25116 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_47
timestamp 1688980957
transform 1 0 5428 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_78
timestamp 1688980957
transform 1 0 8280 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_209
timestamp 1688980957
transform 1 0 20332 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_222
timestamp 1688980957
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_246
timestamp 1688980957
transform 1 0 23736 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_258
timestamp 1688980957
transform 1 0 24840 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_270
timestamp 1688980957
transform 1 0 25944 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_113
timestamp 1688980957
transform 1 0 11500 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_137
timestamp 1688980957
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_156
timestamp 1688980957
transform 1 0 15456 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_160
timestamp 1688980957
transform 1 0 15824 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_194
timestamp 1688980957
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_240
timestamp 1688980957
transform 1 0 23184 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_9
timestamp 1688980957
transform 1 0 1932 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_21
timestamp 1688980957
transform 1 0 3036 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_35
timestamp 1688980957
transform 1 0 4324 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_47
timestamp 1688980957
transform 1 0 5428 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_65
timestamp 1688980957
transform 1 0 7084 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_85
timestamp 1688980957
transform 1 0 8924 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_104
timestamp 1688980957
transform 1 0 10672 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_118
timestamp 1688980957
transform 1 0 11960 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_135
timestamp 1688980957
transform 1 0 13524 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_139
timestamp 1688980957
transform 1 0 13892 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_141
timestamp 1688980957
transform 1 0 14076 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_153
timestamp 1688980957
transform 1 0 15180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_163
timestamp 1688980957
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_173
timestamp 1688980957
transform 1 0 17020 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_185
timestamp 1688980957
transform 1 0 18124 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_193
timestamp 1688980957
transform 1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_197
timestamp 1688980957
transform 1 0 19228 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_202
timestamp 1688980957
transform 1 0 19688 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_208
timestamp 1688980957
transform 1 0 20240 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_218
timestamp 1688980957
transform 1 0 21160 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_237
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_244
timestamp 1688980957
transform 1 0 23552 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_253
timestamp 1688980957
transform 1 0 24380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_265
timestamp 1688980957
transform 1 0 25484 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 23184 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 25116 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 17480 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 25116 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 4232 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 7452 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 23092 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 21804 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform -1 0 22540 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform -1 0 21528 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 11960 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 25852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 22816 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 22264 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform -1 0 5980 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 25116 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 25024 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform -1 0 6256 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 23184 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform 1 0 23368 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform -1 0 22540 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform -1 0 20332 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform -1 0 24012 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform 1 0 23092 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform -1 0 3680 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform -1 0 21528 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 21620 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform -1 0 23644 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 24472 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform -1 0 25944 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform -1 0 25116 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform -1 0 24380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform -1 0 21712 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform 1 0 4876 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform -1 0 19228 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform -1 0 8096 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform -1 0 23092 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 7820 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform -1 0 17020 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform -1 0 12880 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform -1 0 20608 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform -1 0 7636 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform -1 0 13340 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform -1 0 19964 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform -1 0 8924 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform -1 0 13064 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform -1 0 18492 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform -1 0 8280 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform -1 0 12604 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform -1 0 18952 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform -1 0 17480 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform -1 0 16560 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform -1 0 12696 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform -1 0 14812 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform -1 0 16192 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform 1 0 18584 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform -1 0 10396 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform -1 0 18400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform -1 0 13340 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform -1 0 10764 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform -1 0 10948 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform -1 0 15548 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform -1 0 17388 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform -1 0 13248 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform -1 0 19044 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform -1 0 11040 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform 1 0 15180 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform -1 0 19044 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform -1 0 17388 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform 1 0 19136 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform -1 0 11500 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform -1 0 14720 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform -1 0 16008 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform -1 0 14812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform -1 0 10948 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform -1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform -1 0 16284 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform -1 0 22448 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform -1 0 19780 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform -1 0 10948 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform -1 0 13340 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform -1 0 18492 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform -1 0 23644 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform 1 0 4876 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform -1 0 10856 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform 1 0 22632 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform -1 0 17388 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform 1 0 20516 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform 1 0 22448 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform -1 0 20056 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform -1 0 23920 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform -1 0 9108 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform -1 0 24288 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform -1 0 18032 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform -1 0 20792 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform -1 0 19504 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 7176 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform -1 0 11960 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26036 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 23276 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 25760 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 19688 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 25760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap28
timestamp 1688980957
transform 1 0 12788 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 1688980957
transform -1 0 1932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 1688980957
transform -1 0 4324 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1688980957
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1688980957
transform -1 0 4508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1688980957
transform 1 0 7820 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1688980957
transform -1 0 12236 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25668 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1688980957
transform 1 0 25668 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1688980957
transform -1 0 1932 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1688980957
transform 1 0 15548 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1688980957
transform -1 0 16100 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1688980957
transform -1 0 1932 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform -1 0 1932 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1688980957
transform 1 0 25668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 26312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 26312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 26312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 26312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 26312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 26312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 26312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 26312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 26312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 26312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 26312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 26312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 26312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 26312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 26312 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 26312 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 26312 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 26312 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 26312 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 26312 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 26312 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 26312 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 26312 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 26312 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 26312 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 26312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 26312 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 26312 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 26312 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 26312 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 26312 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 26312 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 26312 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 26312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 26312 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 26312 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 26312 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 26312 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 26312 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 26312 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 26312 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 26312 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 26312 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 26312 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 26312 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 26312 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 3680 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 8832 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 13984 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 19136 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 24288 0 -1 27200
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 blue
port 0 nsew signal tristate
flabel metal2 s 27066 28809 27122 29609 0 FreeSans 224 90 0 0 clk
port 1 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 nrst
port 2 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 pb[0]
port 3 nsew signal input
flabel metal2 s 7102 28809 7158 29609 0 FreeSans 224 90 0 0 pb[1]
port 4 nsew signal input
flabel metal2 s 11610 28809 11666 29609 0 FreeSans 224 90 0 0 pb[2]
port 5 nsew signal input
flabel metal3 s 26665 8168 27465 8288 0 FreeSans 480 0 0 0 pb[3]
port 6 nsew signal input
flabel metal2 s 23202 28809 23258 29609 0 FreeSans 224 90 0 0 pb[4]
port 7 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 pb[5]
port 8 nsew signal input
flabel metal3 s 26665 17008 27465 17128 0 FreeSans 480 0 0 0 pb[6]
port 9 nsew signal input
flabel metal2 s 19338 28809 19394 29609 0 FreeSans 224 90 0 0 pb[7]
port 10 nsew signal input
flabel metal3 s 26665 8 27465 128 0 FreeSans 480 0 0 0 pb[8]
port 11 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 pb[9]
port 12 nsew signal input
flabel metal2 s 3238 28809 3294 29609 0 FreeSans 224 90 0 0 red
port 13 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 ss[0]
port 14 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 ss[10]
port 15 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 ss[11]
port 16 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 ss[12]
port 17 nsew signal tristate
flabel metal3 s 26665 4088 27465 4208 0 FreeSans 480 0 0 0 ss[13]
port 18 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 ss[1]
port 19 nsew signal tristate
flabel metal3 s 26665 21088 27465 21208 0 FreeSans 480 0 0 0 ss[2]
port 20 nsew signal tristate
flabel metal3 s 26665 25168 27465 25288 0 FreeSans 480 0 0 0 ss[3]
port 21 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 ss[4]
port 22 nsew signal tristate
flabel metal2 s 15474 28809 15530 29609 0 FreeSans 224 90 0 0 ss[5]
port 23 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 ss[6]
port 24 nsew signal tristate
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 ss[7]
port 25 nsew signal tristate
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 ss[8]
port 26 nsew signal tristate
flabel metal3 s 26665 12928 27465 13048 0 FreeSans 480 0 0 0 ss[9]
port 27 nsew signal tristate
flabel metal4 s 4095 2128 4415 27248 0 FreeSans 1920 90 0 0 vccd1
port 28 nsew power bidirectional
flabel metal4 s 10397 2128 10717 27248 0 FreeSans 1920 90 0 0 vccd1
port 28 nsew power bidirectional
flabel metal4 s 16699 2128 17019 27248 0 FreeSans 1920 90 0 0 vccd1
port 28 nsew power bidirectional
flabel metal4 s 23001 2128 23321 27248 0 FreeSans 1920 90 0 0 vccd1
port 28 nsew power bidirectional
flabel metal4 s 7246 2128 7566 27248 0 FreeSans 1920 90 0 0 vssd1
port 29 nsew ground bidirectional
flabel metal4 s 13548 2128 13868 27248 0 FreeSans 1920 90 0 0 vssd1
port 29 nsew ground bidirectional
flabel metal4 s 19850 2128 20170 27248 0 FreeSans 1920 90 0 0 vssd1
port 29 nsew ground bidirectional
flabel metal4 s 26152 2128 26472 27248 0 FreeSans 1920 90 0 0 vssd1
port 29 nsew ground bidirectional
rlabel metal1 13708 26656 13708 26656 0 vccd1
rlabel via1 13788 27200 13788 27200 0 vssd1
rlabel metal2 22126 16558 22126 16558 0 _0000_
rlabel metal1 19734 21624 19734 21624 0 _0001_
rlabel metal2 23506 16150 23506 16150 0 _0002_
rlabel metal1 21015 10234 21015 10234 0 _0003_
rlabel metal2 21574 10914 21574 10914 0 _0004_
rlabel metal1 22540 10574 22540 10574 0 _0005_
rlabel metal1 23966 19346 23966 19346 0 _0006_
rlabel metal1 20884 14858 20884 14858 0 _0007_
rlabel metal1 20470 19278 20470 19278 0 _0008_
rlabel metal1 23092 17714 23092 17714 0 _0009_
rlabel metal2 21022 18530 21022 18530 0 _0010_
rlabel metal1 25622 10234 25622 10234 0 _0011_
rlabel metal1 19458 10778 19458 10778 0 _0012_
rlabel metal2 20746 8194 20746 8194 0 _0013_
rlabel metal1 18676 11322 18676 11322 0 _0014_
rlabel metal1 16836 23290 16836 23290 0 _0015_
rlabel metal1 7866 17850 7866 17850 0 _0016_
rlabel metal1 5474 15368 5474 15368 0 _0017_
rlabel metal2 14122 21114 14122 21114 0 _0018_
rlabel metal1 7038 15130 7038 15130 0 _0019_
rlabel metal1 6578 19720 6578 19720 0 _0020_
rlabel metal1 6118 21046 6118 21046 0 _0021_
rlabel metal2 6946 23426 6946 23426 0 _0022_
rlabel metal1 7222 22746 7222 22746 0 _0023_
rlabel metal1 5520 13362 5520 13362 0 _0024_
rlabel metal1 1702 6392 1702 6392 0 _0025_
rlabel metal1 4370 22984 4370 22984 0 _0026_
rlabel metal1 3220 13974 3220 13974 0 _0027_
rlabel metal1 2109 15674 2109 15674 0 _0028_
rlabel metal1 2024 16762 2024 16762 0 _0029_
rlabel metal1 1978 15062 1978 15062 0 _0030_
rlabel metal1 2070 18394 2070 18394 0 _0031_
rlabel metal1 2024 19414 2024 19414 0 _0032_
rlabel metal1 2162 19890 2162 19890 0 _0033_
rlabel metal1 3128 21114 3128 21114 0 _0034_
rlabel metal1 17020 25942 17020 25942 0 _0035_
rlabel metal1 17342 19278 17342 19278 0 _0036_
rlabel metal1 14168 17578 14168 17578 0 _0037_
rlabel metal2 13938 21726 13938 21726 0 _0038_
rlabel metal1 9016 16490 9016 16490 0 _0039_
rlabel metal2 9246 20060 9246 20060 0 _0040_
rlabel metal1 8786 21862 8786 21862 0 _0041_
rlabel metal1 8878 25466 8878 25466 0 _0042_
rlabel metal1 12512 25942 12512 25942 0 _0043_
rlabel metal1 18354 24310 18354 24310 0 _0044_
rlabel metal1 19182 17850 19182 17850 0 _0045_
rlabel metal1 14986 16762 14986 16762 0 _0046_
rlabel metal2 17434 21420 17434 21420 0 _0047_
rlabel metal2 11822 17442 11822 17442 0 _0048_
rlabel metal1 11270 19754 11270 19754 0 _0049_
rlabel metal2 10994 22168 10994 22168 0 _0050_
rlabel metal1 10573 25466 10573 25466 0 _0051_
rlabel metal1 13478 23800 13478 23800 0 _0052_
rlabel metal1 16461 24378 16461 24378 0 _0053_
rlabel metal2 17434 18530 17434 18530 0 _0054_
rlabel metal1 14812 16150 14812 16150 0 _0055_
rlabel metal2 16514 21726 16514 21726 0 _0056_
rlabel metal1 10994 16626 10994 16626 0 _0057_
rlabel metal1 11592 19278 11592 19278 0 _0058_
rlabel metal1 10442 23154 10442 23154 0 _0059_
rlabel metal1 10028 24378 10028 24378 0 _0060_
rlabel metal1 13202 24378 13202 24378 0 _0061_
rlabel metal1 17020 9622 17020 9622 0 _0062_
rlabel metal1 17296 12410 17296 12410 0 _0063_
rlabel metal2 16330 13532 16330 13532 0 _0064_
rlabel metal1 16047 10234 16047 10234 0 _0065_
rlabel metal1 11316 14450 11316 14450 0 _0066_
rlabel metal1 11776 15062 11776 15062 0 _0067_
rlabel metal1 9292 13974 9292 13974 0 _0068_
rlabel metal2 9890 14110 9890 14110 0 _0069_
rlabel metal2 14398 14892 14398 14892 0 _0070_
rlabel metal2 11914 12206 11914 12206 0 _0071_
rlabel metal1 8648 12410 8648 12410 0 _0072_
rlabel metal1 10764 12614 10764 12614 0 _0073_
rlabel metal1 11822 11186 11822 11186 0 _0074_
rlabel metal1 2392 11866 2392 11866 0 _0075_
rlabel metal1 4554 11832 4554 11832 0 _0076_
rlabel metal1 3680 10710 3680 10710 0 _0077_
rlabel metal1 2070 9010 2070 9010 0 _0078_
rlabel metal1 17296 7786 17296 7786 0 _0079_
rlabel metal1 18952 4794 18952 4794 0 _0080_
rlabel metal1 18492 3094 18492 3094 0 _0081_
rlabel metal1 16560 3162 16560 3162 0 _0082_
rlabel metal1 11539 6970 11539 6970 0 _0083_
rlabel metal2 12374 3298 12374 3298 0 _0084_
rlabel metal1 11171 3706 11171 3706 0 _0085_
rlabel metal1 11362 4250 11362 4250 0 _0086_
rlabel metal1 15502 9010 15502 9010 0 _0087_
rlabel metal1 18998 7480 18998 7480 0 _0088_
rlabel metal2 18630 6426 18630 6426 0 _0089_
rlabel metal1 14766 3400 14766 3400 0 _0090_
rlabel metal1 14858 3094 14858 3094 0 _0091_
rlabel metal1 9890 3128 9890 3128 0 _0092_
rlabel metal1 8142 3706 8142 3706 0 _0093_
rlabel metal1 6256 3162 6256 3162 0 _0094_
rlabel metal1 9384 6358 9384 6358 0 _0095_
rlabel metal1 13156 9146 13156 9146 0 _0096_
rlabel metal1 15318 25806 15318 25806 0 _0097_
rlabel metal1 15042 18938 15042 18938 0 _0098_
rlabel metal2 13662 18020 13662 18020 0 _0099_
rlabel metal1 14398 20808 14398 20808 0 _0100_
rlabel metal1 8779 15878 8779 15878 0 _0101_
rlabel metal1 8648 19414 8648 19414 0 _0102_
rlabel metal1 8510 22712 8510 22712 0 _0103_
rlabel metal1 8832 25126 8832 25126 0 _0104_
rlabel via1 12183 25466 12183 25466 0 _0105_
rlabel metal1 21436 25330 21436 25330 0 _0106_
rlabel metal1 21840 21114 21840 21114 0 _0107_
rlabel metal1 23966 23800 23966 23800 0 _0108_
rlabel metal1 19366 22712 19366 22712 0 _0109_
rlabel metal2 21298 24548 21298 24548 0 _0110_
rlabel metal1 22402 22542 22402 22542 0 _0111_
rlabel metal1 19320 23018 19320 23018 0 _0112_
rlabel metal2 25898 9860 25898 9860 0 _0113_
rlabel via1 22116 6766 22116 6766 0 _0114_
rlabel metal1 22218 6630 22218 6630 0 _0115_
rlabel metal2 21344 14450 21344 14450 0 _0116_
rlabel metal1 24932 13498 24932 13498 0 _0117_
rlabel metal1 24978 13226 24978 13226 0 _0118_
rlabel metal2 24426 13668 24426 13668 0 _0119_
rlabel metal1 21206 15028 21206 15028 0 _0120_
rlabel metal1 20746 16524 20746 16524 0 _0121_
rlabel metal1 21252 20230 21252 20230 0 _0122_
rlabel metal1 20148 12818 20148 12818 0 _0123_
rlabel metal1 20608 12614 20608 12614 0 _0124_
rlabel metal1 21206 18326 21206 18326 0 _0125_
rlabel metal1 6532 24378 6532 24378 0 _0126_
rlabel metal2 21942 24735 21942 24735 0 _0127_
rlabel metal1 22678 23052 22678 23052 0 _0128_
rlabel metal1 23046 6902 23046 6902 0 _0129_
rlabel metal1 21666 11730 21666 11730 0 _0130_
rlabel metal1 22908 15674 22908 15674 0 _0131_
rlabel metal1 22172 10234 22172 10234 0 _0132_
rlabel metal1 18078 14790 18078 14790 0 _0133_
rlabel metal1 19090 11084 19090 11084 0 _0134_
rlabel metal1 21252 8534 21252 8534 0 _0135_
rlabel metal1 24334 19686 24334 19686 0 _0136_
rlabel metal1 23552 19754 23552 19754 0 _0137_
rlabel metal1 21390 19822 21390 19822 0 _0138_
rlabel metal2 15594 11917 15594 11917 0 _0139_
rlabel metal1 13892 12818 13892 12818 0 _0140_
rlabel metal1 15088 11526 15088 11526 0 _0141_
rlabel metal1 14720 11594 14720 11594 0 _0142_
rlabel metal1 14674 12172 14674 12172 0 _0143_
rlabel metal1 14812 11730 14812 11730 0 _0144_
rlabel metal1 14720 12070 14720 12070 0 _0145_
rlabel metal1 16008 12886 16008 12886 0 _0146_
rlabel metal1 14766 12954 14766 12954 0 _0147_
rlabel metal2 15594 13056 15594 13056 0 _0148_
rlabel metal1 15962 12784 15962 12784 0 _0149_
rlabel metal2 13202 13124 13202 13124 0 _0150_
rlabel metal1 15134 12886 15134 12886 0 _0151_
rlabel metal1 15778 11764 15778 11764 0 _0152_
rlabel metal1 21804 13974 21804 13974 0 _0153_
rlabel metal1 22172 13906 22172 13906 0 _0154_
rlabel metal2 21666 14076 21666 14076 0 _0155_
rlabel metal1 22034 14484 22034 14484 0 _0156_
rlabel metal2 3726 8874 3726 8874 0 _0157_
rlabel metal1 3864 8942 3864 8942 0 _0158_
rlabel metal1 2438 8432 2438 8432 0 _0159_
rlabel metal1 2300 8262 2300 8262 0 _0160_
rlabel metal1 4232 8942 4232 8942 0 _0161_
rlabel metal1 2346 8364 2346 8364 0 _0162_
rlabel metal1 3910 8500 3910 8500 0 _0163_
rlabel metal1 2944 9350 2944 9350 0 _0164_
rlabel metal1 4508 9962 4508 9962 0 _0165_
rlabel metal1 16330 9928 16330 9928 0 _0166_
rlabel metal2 2438 8262 2438 8262 0 _0167_
rlabel metal2 4922 8738 4922 8738 0 _0168_
rlabel metal1 3358 8398 3358 8398 0 _0169_
rlabel metal1 3772 7854 3772 7854 0 _0170_
rlabel metal1 21114 16218 21114 16218 0 _0171_
rlabel metal1 23552 15470 23552 15470 0 _0172_
rlabel metal1 20562 21998 20562 21998 0 _0173_
rlabel metal1 21068 16626 21068 16626 0 _0174_
rlabel metal1 5382 17204 5382 17204 0 _0175_
rlabel metal2 5566 17612 5566 17612 0 _0176_
rlabel metal1 6854 17136 6854 17136 0 _0177_
rlabel metal1 5980 16626 5980 16626 0 _0178_
rlabel metal1 6900 17034 6900 17034 0 _0179_
rlabel metal1 6762 17306 6762 17306 0 _0180_
rlabel metal1 7958 17680 7958 17680 0 _0181_
rlabel metal1 7728 17646 7728 17646 0 _0182_
rlabel metal1 5060 16762 5060 16762 0 _0183_
rlabel metal1 6164 16490 6164 16490 0 _0184_
rlabel metal1 7682 16184 7682 16184 0 _0185_
rlabel metal1 6394 14960 6394 14960 0 _0186_
rlabel metal2 6026 17153 6026 17153 0 _0187_
rlabel metal1 6348 17850 6348 17850 0 _0188_
rlabel metal2 14490 20587 14490 20587 0 _0189_
rlabel metal1 7130 14892 7130 14892 0 _0190_
rlabel metal1 5796 13294 5796 13294 0 _0191_
rlabel metal1 7084 14586 7084 14586 0 _0192_
rlabel metal1 5014 17306 5014 17306 0 _0193_
rlabel metal1 5934 17850 5934 17850 0 _0194_
rlabel metal1 5796 19482 5796 19482 0 _0195_
rlabel metal1 5336 19346 5336 19346 0 _0196_
rlabel metal1 5704 18938 5704 18938 0 _0197_
rlabel metal2 5382 20196 5382 20196 0 _0198_
rlabel metal1 5888 20366 5888 20366 0 _0199_
rlabel metal1 5566 20298 5566 20298 0 _0200_
rlabel metal1 7038 20570 7038 20570 0 _0201_
rlabel metal1 5244 20026 5244 20026 0 _0202_
rlabel metal2 5750 20060 5750 20060 0 _0203_
rlabel metal2 4922 20264 4922 20264 0 _0204_
rlabel metal2 6762 20842 6762 20842 0 _0205_
rlabel metal1 6670 20808 6670 20808 0 _0206_
rlabel metal1 6578 20978 6578 20978 0 _0207_
rlabel metal1 6394 21114 6394 21114 0 _0208_
rlabel metal1 6072 13294 6072 13294 0 _0209_
rlabel metal2 8326 14144 8326 14144 0 _0210_
rlabel metal1 6256 13974 6256 13974 0 _0211_
rlabel metal1 18078 5236 18078 5236 0 _0212_
rlabel metal1 17802 5168 17802 5168 0 _0213_
rlabel metal1 16054 5644 16054 5644 0 _0214_
rlabel metal1 13754 6800 13754 6800 0 _0215_
rlabel metal1 17434 6324 17434 6324 0 _0216_
rlabel metal1 17158 6256 17158 6256 0 _0217_
rlabel metal1 16928 6766 16928 6766 0 _0218_
rlabel metal2 15686 7616 15686 7616 0 _0219_
rlabel metal1 16652 6834 16652 6834 0 _0220_
rlabel metal1 14996 7514 14996 7514 0 _0221_
rlabel metal1 14122 6698 14122 6698 0 _0222_
rlabel metal1 13938 7378 13938 7378 0 _0223_
rlabel metal1 14582 5134 14582 5134 0 _0224_
rlabel metal1 17020 4658 17020 4658 0 _0225_
rlabel metal1 13938 6290 13938 6290 0 _0226_
rlabel metal1 12972 6766 12972 6766 0 _0227_
rlabel metal1 13892 6426 13892 6426 0 _0228_
rlabel metal1 12926 6970 12926 6970 0 _0229_
rlabel metal2 12098 8160 12098 8160 0 _0230_
rlabel metal2 16054 8126 16054 8126 0 _0231_
rlabel metal1 12926 8398 12926 8398 0 _0232_
rlabel metal1 13892 6970 13892 6970 0 _0233_
rlabel metal1 13478 8534 13478 8534 0 _0234_
rlabel metal2 12374 8636 12374 8636 0 _0235_
rlabel metal1 13156 7446 13156 7446 0 _0236_
rlabel metal1 9154 5236 9154 5236 0 _0237_
rlabel metal2 9614 6154 9614 6154 0 _0238_
rlabel metal1 12604 7922 12604 7922 0 _0239_
rlabel via1 8326 6767 8326 6767 0 _0240_
rlabel metal1 9476 5202 9476 5202 0 _0241_
rlabel metal2 9154 5338 9154 5338 0 _0242_
rlabel metal1 9192 5542 9192 5542 0 _0243_
rlabel metal1 8694 6086 8694 6086 0 _0244_
rlabel metal1 8142 6188 8142 6188 0 _0245_
rlabel metal1 8556 6426 8556 6426 0 _0246_
rlabel metal1 6946 7446 6946 7446 0 _0247_
rlabel metal1 6026 5678 6026 5678 0 _0248_
rlabel metal2 13386 4794 13386 4794 0 _0249_
rlabel metal1 6026 4663 6026 4663 0 _0250_
rlabel metal1 7590 4114 7590 4114 0 _0251_
rlabel metal1 6210 4624 6210 4624 0 _0252_
rlabel metal2 5566 5542 5566 5542 0 _0253_
rlabel metal1 6394 6766 6394 6766 0 _0254_
rlabel metal2 7774 8228 7774 8228 0 _0255_
rlabel metal2 6118 4998 6118 4998 0 _0256_
rlabel metal1 5842 5236 5842 5236 0 _0257_
rlabel metal1 5980 6290 5980 6290 0 _0258_
rlabel metal1 12788 4998 12788 4998 0 _0259_
rlabel metal1 6624 5678 6624 5678 0 _0260_
rlabel metal2 7038 4998 7038 4998 0 _0261_
rlabel metal1 6762 5746 6762 5746 0 _0262_
rlabel metal2 5290 6052 5290 6052 0 _0263_
rlabel metal1 6118 7888 6118 7888 0 _0264_
rlabel metal1 14819 8534 14819 8534 0 _0265_
rlabel metal1 6578 6256 6578 6256 0 _0266_
rlabel metal1 6854 5882 6854 5882 0 _0267_
rlabel metal1 6624 7310 6624 7310 0 _0268_
rlabel metal2 7130 8466 7130 8466 0 _0269_
rlabel metal1 7130 7378 7130 7378 0 _0270_
rlabel metal1 8004 8602 8004 8602 0 _0271_
rlabel metal1 6670 9146 6670 9146 0 _0272_
rlabel metal1 8326 12954 8326 12954 0 _0273_
rlabel metal2 9476 12750 9476 12750 0 _0274_
rlabel metal2 6992 12580 6992 12580 0 _0275_
rlabel metal2 8694 9316 8694 9316 0 _0276_
rlabel metal2 8510 9350 8510 9350 0 _0277_
rlabel metal1 8740 9690 8740 9690 0 _0278_
rlabel metal1 2438 6732 2438 6732 0 _0279_
rlabel metal1 22126 17816 22126 17816 0 _0280_
rlabel metal2 22218 17680 22218 17680 0 _0281_
rlabel metal1 22356 23290 22356 23290 0 _0282_
rlabel metal2 21942 22746 21942 22746 0 _0283_
rlabel via2 21574 21947 21574 21947 0 _0284_
rlabel metal1 4876 20978 4876 20978 0 _0285_
rlabel metal1 5658 23766 5658 23766 0 _0286_
rlabel metal1 3634 14382 3634 14382 0 _0287_
rlabel metal2 2530 15878 2530 15878 0 _0288_
rlabel metal1 2530 16422 2530 16422 0 _0289_
rlabel metal1 2254 16048 2254 16048 0 _0290_
rlabel metal1 2576 18258 2576 18258 0 _0291_
rlabel metal1 2346 20400 2346 20400 0 _0292_
rlabel metal1 2898 20366 2898 20366 0 _0293_
rlabel metal1 3588 20910 3588 20910 0 _0294_
rlabel metal1 18630 16456 18630 16456 0 _0295_
rlabel metal1 15088 17102 15088 17102 0 _0296_
rlabel metal1 17066 25466 17066 25466 0 _0297_
rlabel metal1 16882 19380 16882 19380 0 _0298_
rlabel metal1 14168 17306 14168 17306 0 _0299_
rlabel metal1 13938 21998 13938 21998 0 _0300_
rlabel metal1 8694 16558 8694 16558 0 _0301_
rlabel metal1 9384 20434 9384 20434 0 _0302_
rlabel metal1 9200 21862 9200 21862 0 _0303_
rlabel metal1 9200 25262 9200 25262 0 _0304_
rlabel metal1 12880 26350 12880 26350 0 _0305_
rlabel metal1 19182 15674 19182 15674 0 _0306_
rlabel metal1 17020 20366 17020 20366 0 _0307_
rlabel metal1 18400 23290 18400 23290 0 _0308_
rlabel metal1 18584 17646 18584 17646 0 _0309_
rlabel metal1 14674 16558 14674 16558 0 _0310_
rlabel metal2 17526 21284 17526 21284 0 _0311_
rlabel metal1 11316 17646 11316 17646 0 _0312_
rlabel metal1 10902 19924 10902 19924 0 _0313_
rlabel metal1 11362 21658 11362 21658 0 _0314_
rlabel metal1 11454 24922 11454 24922 0 _0315_
rlabel metal1 14122 24174 14122 24174 0 _0316_
rlabel metal1 18492 16762 18492 16762 0 _0317_
rlabel metal1 19826 18836 19826 18836 0 _0318_
rlabel metal1 17756 24378 17756 24378 0 _0319_
rlabel metal1 17894 18258 17894 18258 0 _0320_
rlabel via1 14950 16541 14950 16541 0 _0321_
rlabel metal1 16606 21896 16606 21896 0 _0322_
rlabel metal1 10488 17170 10488 17170 0 _0323_
rlabel metal1 12742 19720 12742 19720 0 _0324_
rlabel metal2 11546 23222 11546 23222 0 _0325_
rlabel metal1 10488 24174 10488 24174 0 _0326_
rlabel metal1 13202 24174 13202 24174 0 _0327_
rlabel metal1 20792 8602 20792 8602 0 _0328_
rlabel metal1 19550 10574 19550 10574 0 _0329_
rlabel metal1 20148 16150 20148 16150 0 _0330_
rlabel metal1 19964 16082 19964 16082 0 _0331_
rlabel metal1 20148 16014 20148 16014 0 _0332_
rlabel metal1 19688 16490 19688 16490 0 _0333_
rlabel metal2 19366 17850 19366 17850 0 _0334_
rlabel metal1 18308 15606 18308 15606 0 _0335_
rlabel metal1 15042 26248 15042 26248 0 _0336_
rlabel metal1 18906 20400 18906 20400 0 _0337_
rlabel metal1 19274 23664 19274 23664 0 _0338_
rlabel metal2 19642 17204 19642 17204 0 _0339_
rlabel metal1 17342 13804 17342 13804 0 _0340_
rlabel metal2 17526 10948 17526 10948 0 _0341_
rlabel metal2 17066 18122 17066 18122 0 _0342_
rlabel metal2 18032 15028 18032 15028 0 _0343_
rlabel metal1 17572 12206 17572 12206 0 _0344_
rlabel metal1 16652 16082 16652 16082 0 _0345_
rlabel metal1 17250 14042 17250 14042 0 _0346_
rlabel metal1 16422 13974 16422 13974 0 _0347_
rlabel metal1 18400 20434 18400 20434 0 _0348_
rlabel metal1 19136 20230 19136 20230 0 _0349_
rlabel metal1 16514 10642 16514 10642 0 _0350_
rlabel metal1 11638 18258 11638 18258 0 _0351_
rlabel metal2 12834 16490 12834 16490 0 _0352_
rlabel metal1 11408 15130 11408 15130 0 _0353_
rlabel metal1 11454 18734 11454 18734 0 _0354_
rlabel metal1 12512 15402 12512 15402 0 _0355_
rlabel metal1 11960 15470 11960 15470 0 _0356_
rlabel metal1 12857 21522 12857 21522 0 _0357_
rlabel metal2 13938 17646 13938 17646 0 _0358_
rlabel metal1 11086 14042 11086 14042 0 _0359_
rlabel metal2 11454 25466 11454 25466 0 _0360_
rlabel metal1 11914 24378 11914 24378 0 _0361_
rlabel metal1 10074 14314 10074 14314 0 _0362_
rlabel metal1 15548 24786 15548 24786 0 _0363_
rlabel metal1 15226 14042 15226 14042 0 _0364_
rlabel metal1 14168 14042 14168 14042 0 _0365_
rlabel metal1 16008 8466 16008 8466 0 _0366_
rlabel metal1 9154 9452 9154 9452 0 _0367_
rlabel metal1 13064 12410 13064 12410 0 _0368_
rlabel metal2 12098 12886 12098 12886 0 _0369_
rlabel metal1 8004 13158 8004 13158 0 _0370_
rlabel via1 11165 9554 11165 9554 0 _0371_
rlabel metal1 10166 9996 10166 9996 0 _0372_
rlabel metal1 11178 9384 11178 9384 0 _0373_
rlabel metal1 10810 9996 10810 9996 0 _0374_
rlabel metal1 9108 10642 9108 10642 0 _0375_
rlabel metal1 11684 7514 11684 7514 0 _0376_
rlabel metal1 10074 8874 10074 8874 0 _0377_
rlabel metal2 13294 8126 13294 8126 0 _0378_
rlabel metal1 11086 7888 11086 7888 0 _0379_
rlabel metal1 10258 8908 10258 8908 0 _0380_
rlabel metal1 9936 9690 9936 9690 0 _0381_
rlabel metal1 9798 9146 9798 9146 0 _0382_
rlabel metal1 8786 9996 8786 9996 0 _0383_
rlabel metal1 9246 11152 9246 11152 0 _0384_
rlabel metal2 8878 10166 8878 10166 0 _0385_
rlabel metal1 9522 11050 9522 11050 0 _0386_
rlabel metal1 14950 6086 14950 6086 0 _0387_
rlabel metal2 15318 6732 15318 6732 0 _0388_
rlabel metal1 14352 5746 14352 5746 0 _0389_
rlabel metal1 11822 5610 11822 5610 0 _0390_
rlabel metal1 7590 5780 7590 5780 0 _0391_
rlabel metal2 8142 5440 8142 5440 0 _0392_
rlabel metal1 7452 6698 7452 6698 0 _0393_
rlabel metal1 7452 10982 7452 10982 0 _0394_
rlabel metal1 9936 11526 9936 11526 0 _0395_
rlabel metal1 9062 11322 9062 11322 0 _0396_
rlabel metal1 10902 12886 10902 12886 0 _0397_
rlabel metal1 9706 9588 9706 9588 0 _0398_
rlabel metal2 9890 10387 9890 10387 0 _0399_
rlabel metal1 9982 9588 9982 9588 0 _0400_
rlabel metal1 11040 10778 11040 10778 0 _0401_
rlabel metal1 9154 13498 9154 13498 0 _0402_
rlabel metal1 10442 10234 10442 10234 0 _0403_
rlabel metal1 9752 10778 9752 10778 0 _0404_
rlabel metal1 11224 11118 11224 11118 0 _0405_
rlabel metal1 8878 7412 8878 7412 0 _0406_
rlabel metal2 7958 8772 7958 8772 0 _0407_
rlabel metal1 7452 11322 7452 11322 0 _0408_
rlabel metal1 5152 12070 5152 12070 0 _0409_
rlabel metal1 2898 11798 2898 11798 0 _0410_
rlabel metal1 5244 12614 5244 12614 0 _0411_
rlabel metal1 6992 9962 6992 9962 0 _0412_
rlabel via1 7122 10778 7122 10778 0 _0413_
rlabel metal1 6808 10438 6808 10438 0 _0414_
rlabel metal1 6716 11254 6716 11254 0 _0415_
rlabel metal1 6118 11322 6118 11322 0 _0416_
rlabel metal1 6854 10608 6854 10608 0 _0417_
rlabel metal1 7774 8534 7774 8534 0 _0418_
rlabel metal1 7912 8466 7912 8466 0 _0419_
rlabel metal1 6578 10676 6578 10676 0 _0420_
rlabel metal1 6164 10778 6164 10778 0 _0421_
rlabel metal1 6118 9350 6118 9350 0 _0422_
rlabel metal1 6256 10098 6256 10098 0 _0423_
rlabel metal1 6118 9418 6118 9418 0 _0424_
rlabel metal2 6302 12789 6302 12789 0 _0425_
rlabel metal1 4324 10642 4324 10642 0 _0426_
rlabel metal2 5934 7378 5934 7378 0 _0427_
rlabel metal1 5520 10030 5520 10030 0 _0428_
rlabel metal1 6440 10234 6440 10234 0 _0429_
rlabel metal1 5796 10234 5796 10234 0 _0430_
rlabel metal2 6440 12308 6440 12308 0 _0431_
rlabel metal1 2622 10132 2622 10132 0 _0432_
rlabel metal1 17112 8466 17112 8466 0 _0433_
rlabel metal2 19090 5066 19090 5066 0 _0434_
rlabel metal1 18216 3502 18216 3502 0 _0435_
rlabel metal1 16376 3026 16376 3026 0 _0436_
rlabel metal2 12466 6902 12466 6902 0 _0437_
rlabel metal1 13018 3026 13018 3026 0 _0438_
rlabel metal1 12144 3162 12144 3162 0 _0439_
rlabel metal1 11546 4114 11546 4114 0 _0440_
rlabel metal1 14904 9690 14904 9690 0 _0441_
rlabel metal1 19412 7854 19412 7854 0 _0442_
rlabel metal1 19044 5882 19044 5882 0 _0443_
rlabel metal1 14214 3604 14214 3604 0 _0444_
rlabel metal1 15318 4114 15318 4114 0 _0445_
rlabel metal1 10396 4114 10396 4114 0 _0446_
rlabel metal1 8740 3502 8740 3502 0 _0447_
rlabel metal1 7222 3026 7222 3026 0 _0448_
rlabel metal2 10166 6324 10166 6324 0 _0449_
rlabel metal1 13754 8942 13754 8942 0 _0450_
rlabel metal1 17756 14790 17756 14790 0 _0451_
rlabel metal2 14858 19482 14858 19482 0 _0452_
rlabel metal1 15870 26350 15870 26350 0 _0453_
rlabel metal1 14766 18768 14766 18768 0 _0454_
rlabel metal1 13386 17646 13386 17646 0 _0455_
rlabel metal1 13892 20910 13892 20910 0 _0456_
rlabel metal1 9154 15674 9154 15674 0 _0457_
rlabel metal1 9062 18938 9062 18938 0 _0458_
rlabel metal1 9246 21114 9246 21114 0 _0459_
rlabel metal1 8694 24922 8694 24922 0 _0460_
rlabel metal2 12466 26350 12466 26350 0 _0461_
rlabel metal2 20838 25126 20838 25126 0 _0462_
rlabel metal2 21482 20570 21482 20570 0 _0463_
rlabel metal1 23138 23290 23138 23290 0 _0464_
rlabel metal1 19872 23834 19872 23834 0 _0465_
rlabel metal1 22494 24276 22494 24276 0 _0466_
rlabel metal1 22356 22202 22356 22202 0 _0467_
rlabel metal1 18906 23188 18906 23188 0 _0468_
rlabel metal3 820 4148 820 4148 0 blue
rlabel metal1 15318 15096 15318 15096 0 clk
rlabel metal1 15824 14790 15824 14790 0 clknet_0_clk
rlabel metal2 1426 4930 1426 4930 0 clknet_4_0_0_clk
rlabel metal1 23874 8500 23874 8500 0 clknet_4_10_0_clk
rlabel metal1 20286 13838 20286 13838 0 clknet_4_11_0_clk
rlabel metal1 16882 19278 16882 19278 0 clknet_4_12_0_clk
rlabel metal1 19320 22066 19320 22066 0 clknet_4_13_0_clk
rlabel metal2 20470 15232 20470 15232 0 clknet_4_14_0_clk
rlabel metal1 24150 24650 24150 24650 0 clknet_4_15_0_clk
rlabel metal2 1610 15266 1610 15266 0 clknet_4_1_0_clk
rlabel metal1 12581 9554 12581 9554 0 clknet_4_2_0_clk
rlabel metal2 14122 15198 14122 15198 0 clknet_4_3_0_clk
rlabel metal2 2714 22066 2714 22066 0 clknet_4_4_0_clk
rlabel metal2 4462 23936 4462 23936 0 clknet_4_5_0_clk
rlabel metal1 14582 17714 14582 17714 0 clknet_4_6_0_clk
rlabel metal2 14490 25602 14490 25602 0 clknet_4_7_0_clk
rlabel metal1 14444 3502 14444 3502 0 clknet_4_8_0_clk
rlabel metal1 17388 12614 17388 12614 0 clknet_4_9_0_clk
rlabel metal1 6578 25160 6578 25160 0 net1
rlabel metal1 25484 2618 25484 2618 0 net10
rlabel metal1 9982 18734 9982 18734 0 net100
rlabel metal1 13708 24174 13708 24174 0 net101
rlabel metal1 16146 17170 16146 17170 0 net102
rlabel metal2 12466 20944 12466 20944 0 net103
rlabel metal1 17158 20400 17158 20400 0 net104
rlabel metal1 10120 20434 10120 20434 0 net105
rlabel metal1 15732 23834 15732 23834 0 net106
rlabel metal1 18078 19686 18078 19686 0 net107
rlabel metal1 16468 17646 16468 17646 0 net108
rlabel metal2 19642 18938 19642 18938 0 net109
rlabel metal1 1656 12410 1656 12410 0 net11
rlabel metal1 9844 25262 9844 25262 0 net110
rlabel metal2 14030 26486 14030 26486 0 net111
rlabel metal1 15042 17306 15042 17306 0 net112
rlabel metal1 13754 19754 13754 19754 0 net113
rlabel metal2 3634 10778 3634 10778 0 net114
rlabel metal1 10028 17306 10028 17306 0 net115
rlabel metal1 9476 24922 9476 24922 0 net116
rlabel metal1 15134 22610 15134 22610 0 net117
rlabel metal1 21528 23834 21528 23834 0 net118
rlabel metal1 18722 23086 18722 23086 0 net119
rlabel metal2 3174 5338 3174 5338 0 net12
rlabel metal1 9936 15470 9936 15470 0 net120
rlabel metal1 12558 12410 12558 12410 0 net121
rlabel metal1 17756 23086 17756 23086 0 net122
rlabel metal1 22678 23800 22678 23800 0 net123
rlabel metal1 6210 11696 6210 11696 0 net124
rlabel metal1 9844 20910 9844 20910 0 net125
rlabel metal1 23368 20026 23368 20026 0 net126
rlabel metal2 17158 5644 17158 5644 0 net127
rlabel metal2 21206 24956 21206 24956 0 net128
rlabel metal1 23690 24208 23690 24208 0 net129
rlabel metal1 5060 13906 5060 13906 0 net13
rlabel metal1 18814 5746 18814 5746 0 net130
rlabel metal1 23046 21658 23046 21658 0 net131
rlabel metal1 7038 22576 7038 22576 0 net132
rlabel metal1 23276 22950 23276 22950 0 net133
rlabel metal1 17204 10778 17204 10778 0 net134
rlabel metal1 19688 5746 19688 5746 0 net135
rlabel metal1 18400 12206 18400 12206 0 net136
rlabel metal1 20470 2346 20470 2346 0 net14
rlabel metal1 2024 2414 2024 2414 0 net15
rlabel metal1 4646 2414 4646 2414 0 net16
rlabel metal1 5221 2482 5221 2482 0 net17
rlabel metal2 16790 4590 16790 4590 0 net18
rlabel metal1 13156 2414 13156 2414 0 net19
rlabel metal2 1656 12852 1656 12852 0 net2
rlabel metal1 25484 20570 25484 20570 0 net20
rlabel via2 15962 12699 15962 12699 0 net21
rlabel metal1 1886 21522 1886 21522 0 net22
rlabel metal1 15548 12886 15548 12886 0 net23
rlabel metal2 15962 2587 15962 2587 0 net24
rlabel metal1 2024 16490 2024 16490 0 net25
rlabel metal2 1794 18190 1794 18190 0 net26
rlabel metal1 25484 11866 25484 11866 0 net27
rlabel metal1 12558 18224 12558 18224 0 net28
rlabel metal1 12558 3400 12558 3400 0 net29
rlabel metal1 6578 26418 6578 26418 0 net3
rlabel metal1 12926 17245 12926 17245 0 net30
rlabel metal2 12650 25432 12650 25432 0 net31
rlabel metal2 21298 3808 21298 3808 0 net32
rlabel metal2 19182 14144 19182 14144 0 net33
rlabel metal2 15502 15266 15502 15266 0 net34
rlabel metal1 21850 15980 21850 15980 0 net35
rlabel metal2 22494 22814 22494 22814 0 net36
rlabel metal1 22678 3706 22678 3706 0 net37
rlabel metal1 22287 26350 22287 26350 0 net38
rlabel metal1 24150 24854 24150 24854 0 net39
rlabel metal1 14674 25330 14674 25330 0 net4
rlabel metal1 18676 25942 18676 25942 0 net40
rlabel metal1 25162 15334 25162 15334 0 net41
rlabel metal1 23966 7480 23966 7480 0 net42
rlabel metal1 3266 22542 3266 22542 0 net43
rlabel metal1 8004 25942 8004 25942 0 net44
rlabel metal1 23874 8602 23874 8602 0 net45
rlabel metal1 20332 20978 20332 20978 0 net46
rlabel metal2 21666 8636 21666 8636 0 net47
rlabel metal1 20286 9622 20286 9622 0 net48
rlabel metal2 20746 12648 20746 12648 0 net49
rlabel metal1 23782 17646 23782 17646 0 net5
rlabel metal2 25162 7684 25162 7684 0 net50
rlabel metal2 23506 5712 23506 5712 0 net51
rlabel metal2 23000 7446 23000 7446 0 net52
rlabel metal1 5014 23834 5014 23834 0 net53
rlabel metal1 23966 11322 23966 11322 0 net54
rlabel metal1 25576 13974 25576 13974 0 net55
rlabel metal1 5336 25330 5336 25330 0 net56
rlabel metal1 22632 12954 22632 12954 0 net57
rlabel metal1 23966 19686 23966 19686 0 net58
rlabel metal2 21850 9316 21850 9316 0 net59
rlabel metal1 22356 25942 22356 25942 0 net6
rlabel metal2 18998 11594 18998 11594 0 net60
rlabel metal2 22494 17476 22494 17476 0 net61
rlabel metal2 23782 18088 23782 18088 0 net62
rlabel metal1 2852 6766 2852 6766 0 net63
rlabel metal1 20286 10710 20286 10710 0 net64
rlabel metal2 20746 22039 20746 22039 0 net65
rlabel metal2 22126 18734 22126 18734 0 net66
rlabel metal1 25668 9962 25668 9962 0 net67
rlabel metal1 24932 9554 24932 9554 0 net68
rlabel metal1 24242 19482 24242 19482 0 net69
rlabel metal1 20194 2618 20194 2618 0 net7
rlabel metal1 23230 18802 23230 18802 0 net70
rlabel metal1 21206 15878 21206 15878 0 net71
rlabel metal1 5750 13974 5750 13974 0 net72
rlabel metal1 16238 22984 16238 22984 0 net73
rlabel metal1 6900 20944 6900 20944 0 net74
rlabel metal1 24288 6970 24288 6970 0 net75
rlabel metal1 21666 6358 21666 6358 0 net76
rlabel metal1 6808 19482 6808 19482 0 net77
rlabel metal1 16192 18734 16192 18734 0 net78
rlabel metal1 11178 24174 11178 24174 0 net79
rlabel metal1 25714 16966 25714 16966 0 net8
rlabel metal1 18170 17680 18170 17680 0 net80
rlabel metal2 6946 16354 6946 16354 0 net81
rlabel metal1 12236 17578 12236 17578 0 net82
rlabel metal1 18814 24106 18814 24106 0 net83
rlabel metal1 7912 14926 7912 14926 0 net84
rlabel metal1 12144 21658 12144 21658 0 net85
rlabel metal1 17388 21930 17388 21930 0 net86
rlabel metal1 6946 23018 6946 23018 0 net87
rlabel metal2 11914 25568 11914 25568 0 net88
rlabel metal2 17434 25738 17434 25738 0 net89
rlabel metal1 19596 25330 19596 25330 0 net9
rlabel metal1 16560 26282 16560 26282 0 net90
rlabel metal1 15134 21658 15134 21658 0 net91
rlabel metal1 11960 22746 11960 22746 0 net92
rlabel metal1 13754 26282 13754 26282 0 net93
rlabel metal1 15364 22202 15364 22202 0 net94
rlabel metal1 18630 9044 18630 9044 0 net95
rlabel metal1 8947 17578 8947 17578 0 net96
rlabel metal1 17480 16490 17480 16490 0 net97
rlabel metal1 12282 16660 12282 16660 0 net98
rlabel metal1 9752 21930 9752 21930 0 net99
rlabel metal3 820 25228 820 25228 0 nrst
rlabel metal3 1004 8228 1004 8228 0 pb[0]
rlabel metal1 7268 26962 7268 26962 0 pb[1]
rlabel metal1 11684 26962 11684 26962 0 pb[2]
rlabel metal2 25990 8075 25990 8075 0 pb[3]
rlabel metal1 23506 27030 23506 27030 0 pb[4]
rlabel metal2 20010 823 20010 823 0 pb[5]
rlabel metal1 25990 17136 25990 17136 0 pb[6]
rlabel metal1 19412 26962 19412 26962 0 pb[7]
rlabel metal1 25392 2414 25392 2414 0 pb[8]
rlabel metal3 820 12308 820 12308 0 pb[9]
rlabel metal1 3588 27098 3588 27098 0 red
rlabel metal2 23874 1520 23874 1520 0 ss[0]
rlabel metal2 46 1554 46 1554 0 ss[10]
rlabel metal2 3910 959 3910 959 0 ss[11]
rlabel metal2 7774 1520 7774 1520 0 ss[12]
rlabel metal1 25944 4454 25944 4454 0 ss[13]
rlabel metal2 11638 959 11638 959 0 ss[1]
rlabel metal2 25898 21233 25898 21233 0 ss[2]
rlabel metal1 26128 25466 26128 25466 0 ss[3]
rlabel metal3 820 21148 820 21148 0 ss[4]
rlabel metal2 15778 27999 15778 27999 0 ss[5]
rlabel metal2 15502 959 15502 959 0 ss[6]
rlabel metal3 751 16388 751 16388 0 ss[7]
rlabel metal2 2806 28203 2806 28203 0 ss[8]
rlabel metal2 25898 13345 25898 13345 0 ss[9]
rlabel metal1 13570 12274 13570 12274 0 u1.keycode\[0\]
rlabel metal1 5290 13838 5290 13838 0 u1.keycode\[1\]
rlabel metal1 8142 15980 8142 15980 0 u1.keycode\[2\]
rlabel metal1 5106 15946 5106 15946 0 u1.keycode\[3\]
rlabel metal1 6256 14450 6256 14450 0 u1.keycode\[4\]
rlabel metal1 4784 17646 4784 17646 0 u1.keycode\[5\]
rlabel metal1 4278 17170 4278 17170 0 u1.keycode\[6\]
rlabel metal1 4278 17068 4278 17068 0 u1.keycode\[7\]
rlabel metal1 4508 20842 4508 20842 0 u1.keycode\[8\]
rlabel metal1 3772 13430 3772 13430 0 u1.keypad_async\[0\]
rlabel metal1 7452 26418 7452 26418 0 u1.keypad_async\[1\]
rlabel metal1 6716 24582 6716 24582 0 u1.keypad_i\[0\]
rlabel metal1 7222 24718 7222 24718 0 u1.keypad_i\[1\]
rlabel metal1 5382 22576 5382 22576 0 u1.keypad_sync\[0\]
rlabel metal2 5842 23392 5842 23392 0 u1.keypad_sync\[1\]
rlabel metal1 16882 25398 16882 25398 0 u1.s_e_detect_w.i_signal
rlabel metal1 20976 20230 20976 20230 0 u1.s_e_detect_w.p_signal
rlabel metal1 20470 20434 20470 20434 0 u1.s_e_detect_w.s_signal
rlabel metal1 25162 19346 25162 19346 0 u1.state\[0\]
rlabel metal2 22126 23902 22126 23902 0 u1.state\[10\]
rlabel metal1 24380 17170 24380 17170 0 u1.state\[11\]
rlabel metal1 22448 23562 22448 23562 0 u1.state\[12\]
rlabel metal1 21712 16014 21712 16014 0 u1.state\[13\]
rlabel metal1 22126 23528 22126 23528 0 u1.state\[14\]
rlabel metal1 22172 23086 22172 23086 0 u1.state\[1\]
rlabel metal1 22356 23222 22356 23222 0 u1.state\[2\]
rlabel metal1 18538 13974 18538 13974 0 u1.state\[3\]
rlabel metal1 22770 19856 22770 19856 0 u1.state\[4\]
rlabel metal1 20562 24038 20562 24038 0 u1.state\[6\]
rlabel metal1 24150 19822 24150 19822 0 u1.state\[7\]
rlabel metal2 23506 19108 23506 19108 0 u1.state\[8\]
rlabel metal2 20838 23222 20838 23222 0 u1.state\[9\]
rlabel metal1 21942 21488 21942 21488 0 u1.store_dig
rlabel metal1 22586 6766 22586 6766 0 u3.keypad_13\[0\]
rlabel metal1 22218 6800 22218 6800 0 u3.keypad_13\[1\]
rlabel metal1 24334 25330 24334 25330 0 u3.keypad_async\[0\]
rlabel metal1 21666 3570 21666 3570 0 u3.keypad_async\[1\]
rlabel metal2 22356 24582 22356 24582 0 u3.keypad_sync\[0\]
rlabel metal1 21666 6732 21666 6732 0 u3.keypad_sync\[1\]
rlabel metal2 21574 5916 21574 5916 0 u3.out\[1\]
rlabel metal2 17342 25806 17342 25806 0 u4.op1\[0\]
rlabel metal1 10212 18258 10212 18258 0 u4.op1\[1\]
rlabel metal1 7958 16082 7958 16082 0 u4.op1\[2\]
rlabel metal1 14950 21998 14950 21998 0 u4.op1\[3\]
rlabel metal1 11316 17306 11316 17306 0 u4.op1\[4\]
rlabel metal1 13202 19890 13202 19890 0 u4.op1\[5\]
rlabel metal1 8832 21454 8832 21454 0 u4.op1\[6\]
rlabel metal1 11086 24310 11086 24310 0 u4.op1\[7\]
rlabel metal1 9108 23698 9108 23698 0 u4.op1\[8\]
rlabel metal1 16238 10574 16238 10574 0 u4.result_ready
rlabel metal1 13386 13260 13386 13260 0 u4.ssdec\[0\]
rlabel metal1 14352 13294 14352 13294 0 u4.ssdec\[1\]
rlabel metal1 12880 12274 12880 12274 0 u4.ssdec\[2\]
rlabel metal1 13662 11016 13662 11016 0 u4.ssdec\[3\]
rlabel metal1 3864 12138 3864 12138 0 u4.ssdec\[4\]
rlabel metal1 4922 11594 4922 11594 0 u4.ssdec\[5\]
rlabel metal1 1518 10744 1518 10744 0 u4.ssdec\[6\]
rlabel metal1 4278 10064 4278 10064 0 u4.ssdec\[7\]
rlabel metal1 19826 24106 19826 24106 0 u5.reg1\[0\]
rlabel metal2 18906 18190 18906 18190 0 u5.reg1\[1\]
rlabel metal1 16864 16082 16864 16082 0 u5.reg1\[2\]
rlabel metal1 18584 21318 18584 21318 0 u5.reg1\[3\]
rlabel metal1 12512 16762 12512 16762 0 u5.reg1\[4\]
rlabel metal2 13294 19516 13294 19516 0 u5.reg1\[5\]
rlabel via1 13386 21522 13386 21522 0 u5.reg1\[6\]
rlabel metal1 12581 24242 12581 24242 0 u5.reg1\[7\]
rlabel viali 15686 24786 15686 24786 0 u5.reg1\[8\]
rlabel metal1 18952 24650 18952 24650 0 u5.reg2\[0\]
rlabel metal1 18906 18054 18906 18054 0 u5.reg2\[1\]
rlabel metal1 16790 16592 16790 16592 0 u5.reg2\[2\]
rlabel metal1 18584 20978 18584 20978 0 u5.reg2\[3\]
rlabel metal1 12926 17714 12926 17714 0 u5.reg2\[4\]
rlabel metal1 12880 19686 12880 19686 0 u5.reg2\[5\]
rlabel metal1 13064 21658 13064 21658 0 u5.reg2\[6\]
rlabel metal2 11822 25908 11822 25908 0 u5.reg2\[7\]
rlabel metal1 15180 24718 15180 24718 0 u5.reg2\[8\]
rlabel metal2 18446 26078 18446 26078 0 u5.reg3\[0\]
rlabel metal1 18538 19142 18538 19142 0 u5.reg3\[1\]
rlabel metal1 15594 18258 15594 18258 0 u5.reg3\[2\]
rlabel metal1 15916 21454 15916 21454 0 u5.reg3\[3\]
rlabel metal2 10902 17204 10902 17204 0 u5.reg3\[4\]
rlabel metal1 10764 20026 10764 20026 0 u5.reg3\[5\]
rlabel metal1 10212 21454 10212 21454 0 u5.reg3\[6\]
rlabel metal2 11362 26180 11362 26180 0 u5.reg3\[7\]
rlabel metal1 14306 26350 14306 26350 0 u5.reg3\[8\]
rlabel metal1 17572 26418 17572 26418 0 u5.reg4\[0\]
rlabel metal2 16514 19652 16514 19652 0 u5.reg4\[1\]
rlabel metal1 16192 18190 16192 18190 0 u5.reg4\[2\]
rlabel metal1 16008 21114 16008 21114 0 u5.reg4\[3\]
rlabel metal2 10166 17204 10166 17204 0 u5.reg4\[4\]
rlabel metal1 10488 19278 10488 19278 0 u5.reg4\[5\]
rlabel metal2 10028 21998 10028 21998 0 u5.reg4\[6\]
rlabel metal1 10718 26894 10718 26894 0 u5.reg4\[7\]
rlabel metal2 14582 25636 14582 25636 0 u5.reg4\[8\]
rlabel metal1 19320 14450 19320 14450 0 u5.reg_num\[0\]
rlabel metal1 18262 16048 18262 16048 0 u5.reg_num\[1\]
rlabel metal1 18216 15062 18216 15062 0 u5.reg_num\[2\]
rlabel metal1 18078 9350 18078 9350 0 u5.reg_val\[0\]
rlabel metal1 19044 12750 19044 12750 0 u5.reg_val\[1\]
rlabel metal1 17434 13498 17434 13498 0 u5.reg_val\[2\]
rlabel metal1 17388 9894 17388 9894 0 u5.reg_val\[3\]
rlabel via1 11638 14467 11638 14467 0 u5.reg_val\[4\]
rlabel metal1 13386 14790 13386 14790 0 u5.reg_val\[5\]
rlabel metal1 7774 13906 7774 13906 0 u5.reg_val\[6\]
rlabel metal1 10350 5746 10350 5746 0 u5.reg_val\[7\]
rlabel metal2 14490 14144 14490 14144 0 u5.reg_val\[8\]
rlabel metal1 21899 14042 21899 14042 0 u6.next_reg_num\[0\]
rlabel metal1 19918 13838 19918 13838 0 u6.next_reg_num\[1\]
rlabel metal1 20470 14042 20470 14042 0 u6.next_reg_num\[2\]
rlabel metal1 24242 15538 24242 15538 0 u6.reg_async\[0\]
rlabel metal1 22586 26282 22586 26282 0 u6.reg_async\[1\]
rlabel metal1 23644 6154 23644 6154 0 u6.reg_async\[2\]
rlabel metal1 5336 12954 5336 12954 0 u6.reg_async\[3\]
rlabel metal1 24288 14042 24288 14042 0 u6.reg_i\[0\]
rlabel metal1 24978 12954 24978 12954 0 u6.reg_i\[1\]
rlabel metal1 24886 11866 24886 11866 0 u6.reg_i\[2\]
rlabel metal2 24242 13940 24242 13940 0 u6.reg_i\[3\]
rlabel metal2 23414 14688 23414 14688 0 u6.reg_sync\[0\]
rlabel metal1 22586 26418 22586 26418 0 u6.reg_sync\[1\]
rlabel metal2 22494 14110 22494 14110 0 u6.reg_sync\[2\]
rlabel metal1 23046 14586 23046 14586 0 u6.reg_sync\[3\]
rlabel metal1 21252 9486 21252 9486 0 u7.assign_op1
rlabel metal1 21436 9894 21436 9894 0 u7.assign_op2
rlabel metal2 24978 8364 24978 8364 0 u7.s_e_detect.i_signal
rlabel metal1 25668 8602 25668 8602 0 u7.s_e_detect.p_signal
rlabel metal1 25392 9554 25392 9554 0 u7.s_e_detect.s_signal
rlabel metal1 24472 10574 24472 10574 0 u7.state\[0\]
rlabel metal1 20976 10982 20976 10982 0 u7.state\[4\]
rlabel metal2 21942 8704 21942 8704 0 u7.state\[5\]
rlabel metal1 20148 12750 20148 12750 0 u7.state\[6\]
rlabel metal1 15640 4658 15640 4658 0 u8.b_assign_op1
rlabel metal1 13846 4012 13846 4012 0 u8.b_assign_op2
rlabel metal1 14122 8466 14122 8466 0 u8.buff_opcode\[1\]
rlabel metal1 18124 7514 18124 7514 0 u8.new_op1\[0\]
rlabel metal1 16054 6834 16054 6834 0 u8.new_op1\[1\]
rlabel metal2 15962 4080 15962 4080 0 u8.new_op1\[2\]
rlabel metal1 15962 4182 15962 4182 0 u8.new_op1\[3\]
rlabel metal1 14720 9486 14720 9486 0 u8.new_op1\[8\]
rlabel metal2 9706 3672 9706 3672 0 u8.op1\[4\]
rlabel metal1 9246 4590 9246 4590 0 u8.op1\[5\]
rlabel metal2 7130 4352 7130 4352 0 u8.op1\[6\]
rlabel metal1 9982 6086 9982 6086 0 u8.op1\[7\]
rlabel metal1 16698 7786 16698 7786 0 u8.op2\[0\]
rlabel metal2 18722 5440 18722 5440 0 u8.op2\[1\]
rlabel metal2 17894 3638 17894 3638 0 u8.op2\[2\]
rlabel metal1 17572 4182 17572 4182 0 u8.op2\[3\]
rlabel metal1 12788 6902 12788 6902 0 u8.op2\[4\]
rlabel metal1 8418 5644 8418 5644 0 u8.op2\[5\]
rlabel metal1 12972 4658 12972 4658 0 u8.op2\[6\]
rlabel metal2 12374 4250 12374 4250 0 u8.op2\[7\]
rlabel metal1 15088 8466 15088 8466 0 u8.op2\[8\]
<< properties >>
string FIXED_BBOX 0 0 27465 29609
<< end >>
