// This is the unpowered netlist.
module Guitar_Villains (chip_select,
    clk,
    green_disp,
    n_rst,
    red_disp,
    bottom_row,
    button,
    ss0,
    ss1,
    top_row);
 input chip_select;
 input clk;
 output green_disp;
 input n_rst;
 output red_disp;
 output [6:0] bottom_row;
 input [3:0] button;
 output [6:0] ss0;
 output [6:0] ss1;
 output [6:0] top_row;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire \disp_song.display_note1[0] ;
 wire \disp_song.display_note1[1] ;
 wire \disp_song.display_note1[2] ;
 wire \disp_song.display_note1[3] ;
 wire \disp_song.display_note1[4] ;
 wire \disp_song.display_note1[5] ;
 wire \disp_song.display_note1[6] ;
 wire \disp_song.display_note2[0] ;
 wire \disp_song.display_note2[1] ;
 wire \disp_song.display_note2[2] ;
 wire \disp_song.display_note2[3] ;
 wire \disp_song.display_note2[4] ;
 wire \disp_song.display_note2[5] ;
 wire \disp_song.display_note2[6] ;
 wire \disp_song.mi6.in[0] ;
 wire \disp_song.mi6.in[1] ;
 wire \disp_song.mi6.in[2] ;
 wire \disp_song.mi6.in[3] ;
 wire \disp_song.mi6.in[4] ;
 wire \disp_song.next_green ;
 wire \disp_song.next_red ;
 wire \disp_song.note1[0] ;
 wire \disp_song.note1[10] ;
 wire \disp_song.note1[11] ;
 wire \disp_song.note1[12] ;
 wire \disp_song.note1[13] ;
 wire \disp_song.note1[14] ;
 wire \disp_song.note1[15] ;
 wire \disp_song.note1[16] ;
 wire \disp_song.note1[17] ;
 wire \disp_song.note1[18] ;
 wire \disp_song.note1[19] ;
 wire \disp_song.note1[1] ;
 wire \disp_song.note1[20] ;
 wire \disp_song.note1[21] ;
 wire \disp_song.note1[22] ;
 wire \disp_song.note1[23] ;
 wire \disp_song.note1[24] ;
 wire \disp_song.note1[25] ;
 wire \disp_song.note1[26] ;
 wire \disp_song.note1[27] ;
 wire \disp_song.note1[28] ;
 wire \disp_song.note1[29] ;
 wire \disp_song.note1[2] ;
 wire \disp_song.note1[30] ;
 wire \disp_song.note1[31] ;
 wire \disp_song.note1[3] ;
 wire \disp_song.note1[4] ;
 wire \disp_song.note1[5] ;
 wire \disp_song.note1[6] ;
 wire \disp_song.note1[7] ;
 wire \disp_song.note1[8] ;
 wire \disp_song.note1[9] ;
 wire \disp_song.note2[0] ;
 wire \disp_song.note2[10] ;
 wire \disp_song.note2[11] ;
 wire \disp_song.note2[12] ;
 wire \disp_song.note2[13] ;
 wire \disp_song.note2[14] ;
 wire \disp_song.note2[15] ;
 wire \disp_song.note2[16] ;
 wire \disp_song.note2[17] ;
 wire \disp_song.note2[18] ;
 wire \disp_song.note2[19] ;
 wire \disp_song.note2[1] ;
 wire \disp_song.note2[20] ;
 wire \disp_song.note2[21] ;
 wire \disp_song.note2[22] ;
 wire \disp_song.note2[23] ;
 wire \disp_song.note2[24] ;
 wire \disp_song.note2[25] ;
 wire \disp_song.note2[26] ;
 wire \disp_song.note2[27] ;
 wire \disp_song.note2[28] ;
 wire \disp_song.note2[29] ;
 wire \disp_song.note2[2] ;
 wire \disp_song.note2[30] ;
 wire \disp_song.note2[31] ;
 wire \disp_song.note2[3] ;
 wire \disp_song.note2[4] ;
 wire \disp_song.note2[5] ;
 wire \disp_song.note2[6] ;
 wire \disp_song.note2[7] ;
 wire \disp_song.note2[8] ;
 wire \disp_song.note2[9] ;
 wire \disp_song.toggle_green ;
 wire \disp_song.toggle_red ;
 wire \disp_song.toggle_state ;
 wire \disp_song.um.boton0e.edge_1 ;
 wire \disp_song.um.boton0e.edge_2 ;
 wire \disp_song.um.boton0e.sync_b ;
 wire \disp_song.um.boton1e.edge_1 ;
 wire \disp_song.um.boton1e.edge_2 ;
 wire \disp_song.um.boton1e.sync_b ;
 wire \disp_song.um.boton2e.edge_1 ;
 wire \disp_song.um.boton2e.edge_2 ;
 wire \disp_song.um.boton2e.sync_b ;
 wire \disp_song.um.drum.next_d1[0] ;
 wire \disp_song.um.drum.next_d1[1] ;
 wire \disp_song.um.drum.next_d1[2] ;
 wire \disp_song.um.drum.next_d1[3] ;
 wire \disp_song.um.drum.next_d1[4] ;
 wire \disp_song.um.drum.next_d1[5] ;
 wire \disp_song.um.drum.next_d1[6] ;
 wire \disp_song.um.drum.next_d2[0] ;
 wire \disp_song.um.drum.next_d2[1] ;
 wire \disp_song.um.drum.next_d2[2] ;
 wire \disp_song.um.drum.next_d2[3] ;
 wire \disp_song.um.drum.next_d2[4] ;
 wire \disp_song.um.drum.next_d2[5] ;
 wire \disp_song.um.drum.next_d2[6] ;
 wire \disp_song.um.drum.next_idx1[0] ;
 wire \disp_song.um.drum.next_idx1[1] ;
 wire \disp_song.um.drum.next_idx1[2] ;
 wire \disp_song.um.drum.next_idx1[3] ;
 wire \disp_song.um.drum.next_idx1[4] ;
 wire \disp_song.um.drum.next_idx2[0] ;
 wire \disp_song.um.drum.next_idx2[1] ;
 wire \disp_song.um.drum.next_idx2[2] ;
 wire \disp_song.um.drum.next_idx2[3] ;
 wire \disp_song.um.drum.next_idx2[4] ;
 wire \disp_song.um.drum.next_note1[0] ;
 wire \disp_song.um.drum.next_note1[10] ;
 wire \disp_song.um.drum.next_note1[11] ;
 wire \disp_song.um.drum.next_note1[12] ;
 wire \disp_song.um.drum.next_note1[13] ;
 wire \disp_song.um.drum.next_note1[14] ;
 wire \disp_song.um.drum.next_note1[15] ;
 wire \disp_song.um.drum.next_note1[16] ;
 wire \disp_song.um.drum.next_note1[17] ;
 wire \disp_song.um.drum.next_note1[18] ;
 wire \disp_song.um.drum.next_note1[19] ;
 wire \disp_song.um.drum.next_note1[1] ;
 wire \disp_song.um.drum.next_note1[20] ;
 wire \disp_song.um.drum.next_note1[21] ;
 wire \disp_song.um.drum.next_note1[22] ;
 wire \disp_song.um.drum.next_note1[23] ;
 wire \disp_song.um.drum.next_note1[24] ;
 wire \disp_song.um.drum.next_note1[25] ;
 wire \disp_song.um.drum.next_note1[26] ;
 wire \disp_song.um.drum.next_note1[27] ;
 wire \disp_song.um.drum.next_note1[28] ;
 wire \disp_song.um.drum.next_note1[29] ;
 wire \disp_song.um.drum.next_note1[2] ;
 wire \disp_song.um.drum.next_note1[30] ;
 wire \disp_song.um.drum.next_note1[31] ;
 wire \disp_song.um.drum.next_note1[3] ;
 wire \disp_song.um.drum.next_note1[4] ;
 wire \disp_song.um.drum.next_note1[5] ;
 wire \disp_song.um.drum.next_note1[6] ;
 wire \disp_song.um.drum.next_note1[7] ;
 wire \disp_song.um.drum.next_note1[8] ;
 wire \disp_song.um.drum.next_note1[9] ;
 wire \disp_song.um.drum.next_note2[0] ;
 wire \disp_song.um.drum.next_note2[10] ;
 wire \disp_song.um.drum.next_note2[11] ;
 wire \disp_song.um.drum.next_note2[12] ;
 wire \disp_song.um.drum.next_note2[13] ;
 wire \disp_song.um.drum.next_note2[14] ;
 wire \disp_song.um.drum.next_note2[15] ;
 wire \disp_song.um.drum.next_note2[16] ;
 wire \disp_song.um.drum.next_note2[17] ;
 wire \disp_song.um.drum.next_note2[18] ;
 wire \disp_song.um.drum.next_note2[19] ;
 wire \disp_song.um.drum.next_note2[1] ;
 wire \disp_song.um.drum.next_note2[20] ;
 wire \disp_song.um.drum.next_note2[21] ;
 wire \disp_song.um.drum.next_note2[22] ;
 wire \disp_song.um.drum.next_note2[23] ;
 wire \disp_song.um.drum.next_note2[24] ;
 wire \disp_song.um.drum.next_note2[25] ;
 wire \disp_song.um.drum.next_note2[26] ;
 wire \disp_song.um.drum.next_note2[27] ;
 wire \disp_song.um.drum.next_note2[28] ;
 wire \disp_song.um.drum.next_note2[29] ;
 wire \disp_song.um.drum.next_note2[2] ;
 wire \disp_song.um.drum.next_note2[30] ;
 wire \disp_song.um.drum.next_note2[31] ;
 wire \disp_song.um.drum.next_note2[3] ;
 wire \disp_song.um.drum.next_note2[4] ;
 wire \disp_song.um.drum.next_note2[5] ;
 wire \disp_song.um.drum.next_note2[6] ;
 wire \disp_song.um.drum.next_note2[7] ;
 wire \disp_song.um.drum.next_note2[8] ;
 wire \disp_song.um.drum.next_note2[9] ;
 wire \disp_song.um.idx_note1[0] ;
 wire \disp_song.um.idx_note1[1] ;
 wire \disp_song.um.idx_note1[2] ;
 wire \disp_song.um.idx_note1[3] ;
 wire \disp_song.um.idx_note1[4] ;
 wire \disp_song.um.idx_note2[0] ;
 wire \disp_song.um.idx_note2[1] ;
 wire \disp_song.um.idx_note2[2] ;
 wire \disp_song.um.idx_note2[3] ;
 wire \disp_song.um.idx_note2[4] ;
 wire \disp_song.um.next_position[0] ;
 wire \disp_song.um.next_position[1] ;
 wire \disp_song.um.next_position[2] ;
 wire \disp_song.um.next_position[3] ;
 wire \disp_song.um.next_position[4] ;
 wire \game.addhits.a[0] ;
 wire \game.addhits.a[10] ;
 wire \game.addhits.a[11] ;
 wire \game.addhits.a[12] ;
 wire \game.addhits.a[13] ;
 wire \game.addhits.a[14] ;
 wire \game.addhits.a[15] ;
 wire \game.addhits.a[1] ;
 wire \game.addhits.a[2] ;
 wire \game.addhits.a[3] ;
 wire \game.addhits.a[4] ;
 wire \game.addhits.a[5] ;
 wire \game.addhits.a[6] ;
 wire \game.addhits.a[7] ;
 wire \game.addhits.a[8] ;
 wire \game.addhits.a[9] ;
 wire \game.addhits.add1.b[0] ;
 wire \game.addhits.add1.b[1] ;
 wire \game.addhits.add1.b[2] ;
 wire \game.addhits.add1.b[3] ;
 wire \game.addhits.add2.b[0] ;
 wire \game.addhits.add2.b[1] ;
 wire \game.addhits.add2.b[2] ;
 wire \game.addhits.add2.b[3] ;
 wire \game.addhits.add3.b[0] ;
 wire \game.addhits.add3.b[1] ;
 wire \game.addhits.add3.b[2] ;
 wire \game.addhits.add3.b[3] ;
 wire \game.addhits.add4.b[0] ;
 wire \game.addhits.add4.b[1] ;
 wire \game.addhits.add4.b[2] ;
 wire \game.addhits.add4.b[3] ;
 wire \game.addmisses.a[0] ;
 wire \game.addmisses.a[10] ;
 wire \game.addmisses.a[11] ;
 wire \game.addmisses.a[12] ;
 wire \game.addmisses.a[13] ;
 wire \game.addmisses.a[14] ;
 wire \game.addmisses.a[15] ;
 wire \game.addmisses.a[1] ;
 wire \game.addmisses.a[2] ;
 wire \game.addmisses.a[3] ;
 wire \game.addmisses.a[4] ;
 wire \game.addmisses.a[5] ;
 wire \game.addmisses.a[6] ;
 wire \game.addmisses.a[7] ;
 wire \game.addmisses.a[8] ;
 wire \game.addmisses.a[9] ;
 wire \game.addmisses.add1.b[0] ;
 wire \game.addmisses.add1.b[1] ;
 wire \game.addmisses.add1.b[2] ;
 wire \game.addmisses.add1.b[3] ;
 wire \game.addmisses.add2.b[0] ;
 wire \game.addmisses.add2.b[1] ;
 wire \game.addmisses.add2.b[2] ;
 wire \game.addmisses.add2.b[3] ;
 wire \game.addmisses.add3.b[0] ;
 wire \game.addmisses.add3.b[1] ;
 wire \game.addmisses.add3.b[2] ;
 wire \game.addmisses.add3.b[3] ;
 wire \game.addmisses.add4.b[0] ;
 wire \game.addmisses.add4.b[1] ;
 wire \game.addmisses.add4.b[2] ;
 wire \game.addmisses.add4.b[3] ;
 wire \game.beat_clk ;
 wire \game.counter[0] ;
 wire \game.counter[10] ;
 wire \game.counter[11] ;
 wire \game.counter[12] ;
 wire \game.counter[13] ;
 wire \game.counter[14] ;
 wire \game.counter[15] ;
 wire \game.counter[16] ;
 wire \game.counter[17] ;
 wire \game.counter[18] ;
 wire \game.counter[19] ;
 wire \game.counter[1] ;
 wire \game.counter[20] ;
 wire \game.counter[21] ;
 wire \game.counter[22] ;
 wire \game.counter[2] ;
 wire \game.counter[3] ;
 wire \game.counter[4] ;
 wire \game.counter[5] ;
 wire \game.counter[6] ;
 wire \game.counter[7] ;
 wire \game.counter[8] ;
 wire \game.counter[9] ;
 wire \game.flash_counter[0] ;
 wire \game.flash_counter[10] ;
 wire \game.flash_counter[11] ;
 wire \game.flash_counter[12] ;
 wire \game.flash_counter[13] ;
 wire \game.flash_counter[14] ;
 wire \game.flash_counter[15] ;
 wire \game.flash_counter[16] ;
 wire \game.flash_counter[17] ;
 wire \game.flash_counter[18] ;
 wire \game.flash_counter[19] ;
 wire \game.flash_counter[1] ;
 wire \game.flash_counter[20] ;
 wire \game.flash_counter[21] ;
 wire \game.flash_counter[22] ;
 wire \game.flash_counter[23] ;
 wire \game.flash_counter[2] ;
 wire \game.flash_counter[3] ;
 wire \game.flash_counter[4] ;
 wire \game.flash_counter[5] ;
 wire \game.flash_counter[6] ;
 wire \game.flash_counter[7] ;
 wire \game.flash_counter[8] ;
 wire \game.flash_counter[9] ;
 wire \game.hit_1 ;
 wire \game.hit_2 ;
 wire \game.missed_1 ;
 wire \game.missed_2 ;
 wire \game.out[0] ;
 wire \game.out[10] ;
 wire \game.out[11] ;
 wire \game.out[12] ;
 wire \game.out[13] ;
 wire \game.out[1] ;
 wire \game.out[2] ;
 wire \game.out[3] ;
 wire \game.out[4] ;
 wire \game.out[5] ;
 wire \game.out[6] ;
 wire \game.out[7] ;
 wire \game.out[8] ;
 wire \game.out[9] ;
 wire \game.padded_notes1[0] ;
 wire \game.padded_notes1[10] ;
 wire \game.padded_notes1[11] ;
 wire \game.padded_notes1[12] ;
 wire \game.padded_notes1[13] ;
 wire \game.padded_notes1[14] ;
 wire \game.padded_notes1[15] ;
 wire \game.padded_notes1[16] ;
 wire \game.padded_notes1[17] ;
 wire \game.padded_notes1[18] ;
 wire \game.padded_notes1[19] ;
 wire \game.padded_notes1[1] ;
 wire \game.padded_notes1[20] ;
 wire \game.padded_notes1[21] ;
 wire \game.padded_notes1[22] ;
 wire \game.padded_notes1[23] ;
 wire \game.padded_notes1[24] ;
 wire \game.padded_notes1[25] ;
 wire \game.padded_notes1[26] ;
 wire \game.padded_notes1[27] ;
 wire \game.padded_notes1[28] ;
 wire \game.padded_notes1[29] ;
 wire \game.padded_notes1[2] ;
 wire \game.padded_notes1[30] ;
 wire \game.padded_notes1[31] ;
 wire \game.padded_notes1[3] ;
 wire \game.padded_notes1[4] ;
 wire \game.padded_notes1[5] ;
 wire \game.padded_notes1[6] ;
 wire \game.padded_notes1[7] ;
 wire \game.padded_notes1[8] ;
 wire \game.padded_notes1[9] ;
 wire \game.padded_notes2[0] ;
 wire \game.padded_notes2[10] ;
 wire \game.padded_notes2[11] ;
 wire \game.padded_notes2[12] ;
 wire \game.padded_notes2[13] ;
 wire \game.padded_notes2[14] ;
 wire \game.padded_notes2[15] ;
 wire \game.padded_notes2[16] ;
 wire \game.padded_notes2[17] ;
 wire \game.padded_notes2[18] ;
 wire \game.padded_notes2[19] ;
 wire \game.padded_notes2[1] ;
 wire \game.padded_notes2[20] ;
 wire \game.padded_notes2[21] ;
 wire \game.padded_notes2[22] ;
 wire \game.padded_notes2[23] ;
 wire \game.padded_notes2[24] ;
 wire \game.padded_notes2[25] ;
 wire \game.padded_notes2[26] ;
 wire \game.padded_notes2[27] ;
 wire \game.padded_notes2[28] ;
 wire \game.padded_notes2[29] ;
 wire \game.padded_notes2[2] ;
 wire \game.padded_notes2[30] ;
 wire \game.padded_notes2[31] ;
 wire \game.padded_notes2[3] ;
 wire \game.padded_notes2[4] ;
 wire \game.padded_notes2[5] ;
 wire \game.padded_notes2[6] ;
 wire \game.padded_notes2[7] ;
 wire \game.padded_notes2[8] ;
 wire \game.padded_notes2[9] ;
 wire \game.scoring_button_1.acc[1] ;
 wire \game.scoring_button_1.acc[2] ;
 wire \game.scoring_button_1.check_hit.edge_1 ;
 wire \game.scoring_button_1.check_hit.edge_2 ;
 wire \game.scoring_button_1.check_hit.in ;
 wire \game.scoring_button_1.counts[0] ;
 wire \game.scoring_button_1.counts[10] ;
 wire \game.scoring_button_1.counts[11] ;
 wire \game.scoring_button_1.counts[12] ;
 wire \game.scoring_button_1.counts[13] ;
 wire \game.scoring_button_1.counts[14] ;
 wire \game.scoring_button_1.counts[15] ;
 wire \game.scoring_button_1.counts[16] ;
 wire \game.scoring_button_1.counts[17] ;
 wire \game.scoring_button_1.counts[18] ;
 wire \game.scoring_button_1.counts[19] ;
 wire \game.scoring_button_1.counts[1] ;
 wire \game.scoring_button_1.counts[20] ;
 wire \game.scoring_button_1.counts[21] ;
 wire \game.scoring_button_1.counts[22] ;
 wire \game.scoring_button_1.counts[2] ;
 wire \game.scoring_button_1.counts[3] ;
 wire \game.scoring_button_1.counts[4] ;
 wire \game.scoring_button_1.counts[5] ;
 wire \game.scoring_button_1.counts[6] ;
 wire \game.scoring_button_1.counts[7] ;
 wire \game.scoring_button_1.counts[8] ;
 wire \game.scoring_button_1.counts[9] ;
 wire \game.scoring_button_1.flash_counter_1[0] ;
 wire \game.scoring_button_1.flash_counter_1[10] ;
 wire \game.scoring_button_1.flash_counter_1[11] ;
 wire \game.scoring_button_1.flash_counter_1[12] ;
 wire \game.scoring_button_1.flash_counter_1[13] ;
 wire \game.scoring_button_1.flash_counter_1[14] ;
 wire \game.scoring_button_1.flash_counter_1[15] ;
 wire \game.scoring_button_1.flash_counter_1[16] ;
 wire \game.scoring_button_1.flash_counter_1[17] ;
 wire \game.scoring_button_1.flash_counter_1[18] ;
 wire \game.scoring_button_1.flash_counter_1[19] ;
 wire \game.scoring_button_1.flash_counter_1[1] ;
 wire \game.scoring_button_1.flash_counter_1[20] ;
 wire \game.scoring_button_1.flash_counter_1[21] ;
 wire \game.scoring_button_1.flash_counter_1[22] ;
 wire \game.scoring_button_1.flash_counter_1[2] ;
 wire \game.scoring_button_1.flash_counter_1[3] ;
 wire \game.scoring_button_1.flash_counter_1[4] ;
 wire \game.scoring_button_1.flash_counter_1[5] ;
 wire \game.scoring_button_1.flash_counter_1[6] ;
 wire \game.scoring_button_1.flash_counter_1[7] ;
 wire \game.scoring_button_1.flash_counter_1[8] ;
 wire \game.scoring_button_1.flash_counter_1[9] ;
 wire \game.scoring_button_1.flash_counter_2[0] ;
 wire \game.scoring_button_1.flash_counter_2[10] ;
 wire \game.scoring_button_1.flash_counter_2[11] ;
 wire \game.scoring_button_1.flash_counter_2[12] ;
 wire \game.scoring_button_1.flash_counter_2[13] ;
 wire \game.scoring_button_1.flash_counter_2[14] ;
 wire \game.scoring_button_1.flash_counter_2[15] ;
 wire \game.scoring_button_1.flash_counter_2[16] ;
 wire \game.scoring_button_1.flash_counter_2[17] ;
 wire \game.scoring_button_1.flash_counter_2[18] ;
 wire \game.scoring_button_1.flash_counter_2[19] ;
 wire \game.scoring_button_1.flash_counter_2[1] ;
 wire \game.scoring_button_1.flash_counter_2[20] ;
 wire \game.scoring_button_1.flash_counter_2[21] ;
 wire \game.scoring_button_1.flash_counter_2[22] ;
 wire \game.scoring_button_1.flash_counter_2[2] ;
 wire \game.scoring_button_1.flash_counter_2[3] ;
 wire \game.scoring_button_1.flash_counter_2[4] ;
 wire \game.scoring_button_1.flash_counter_2[5] ;
 wire \game.scoring_button_1.flash_counter_2[6] ;
 wire \game.scoring_button_1.flash_counter_2[7] ;
 wire \game.scoring_button_1.flash_counter_2[8] ;
 wire \game.scoring_button_1.flash_counter_2[9] ;
 wire \game.scoring_button_1.hit ;
 wire \game.scoring_button_1.next_count[0] ;
 wire \game.scoring_button_1.next_count[10] ;
 wire \game.scoring_button_1.next_count[11] ;
 wire \game.scoring_button_1.next_count[12] ;
 wire \game.scoring_button_1.next_count[13] ;
 wire \game.scoring_button_1.next_count[14] ;
 wire \game.scoring_button_1.next_count[15] ;
 wire \game.scoring_button_1.next_count[16] ;
 wire \game.scoring_button_1.next_count[17] ;
 wire \game.scoring_button_1.next_count[18] ;
 wire \game.scoring_button_1.next_count[19] ;
 wire \game.scoring_button_1.next_count[1] ;
 wire \game.scoring_button_1.next_count[20] ;
 wire \game.scoring_button_1.next_count[21] ;
 wire \game.scoring_button_1.next_count[22] ;
 wire \game.scoring_button_1.next_count[2] ;
 wire \game.scoring_button_1.next_count[3] ;
 wire \game.scoring_button_1.next_count[4] ;
 wire \game.scoring_button_1.next_count[5] ;
 wire \game.scoring_button_1.next_count[6] ;
 wire \game.scoring_button_1.next_count[7] ;
 wire \game.scoring_button_1.next_count[8] ;
 wire \game.scoring_button_1.next_count[9] ;
 wire \game.scoring_button_1.next_flash_counter_1[0] ;
 wire \game.scoring_button_1.next_flash_counter_1[10] ;
 wire \game.scoring_button_1.next_flash_counter_1[11] ;
 wire \game.scoring_button_1.next_flash_counter_1[12] ;
 wire \game.scoring_button_1.next_flash_counter_1[13] ;
 wire \game.scoring_button_1.next_flash_counter_1[14] ;
 wire \game.scoring_button_1.next_flash_counter_1[15] ;
 wire \game.scoring_button_1.next_flash_counter_1[16] ;
 wire \game.scoring_button_1.next_flash_counter_1[17] ;
 wire \game.scoring_button_1.next_flash_counter_1[18] ;
 wire \game.scoring_button_1.next_flash_counter_1[19] ;
 wire \game.scoring_button_1.next_flash_counter_1[1] ;
 wire \game.scoring_button_1.next_flash_counter_1[20] ;
 wire \game.scoring_button_1.next_flash_counter_1[21] ;
 wire \game.scoring_button_1.next_flash_counter_1[22] ;
 wire \game.scoring_button_1.next_flash_counter_1[2] ;
 wire \game.scoring_button_1.next_flash_counter_1[3] ;
 wire \game.scoring_button_1.next_flash_counter_1[4] ;
 wire \game.scoring_button_1.next_flash_counter_1[5] ;
 wire \game.scoring_button_1.next_flash_counter_1[6] ;
 wire \game.scoring_button_1.next_flash_counter_1[7] ;
 wire \game.scoring_button_1.next_flash_counter_1[8] ;
 wire \game.scoring_button_1.next_flash_counter_1[9] ;
 wire \game.scoring_button_1.next_flash_counter_2[0] ;
 wire \game.scoring_button_1.next_flash_counter_2[10] ;
 wire \game.scoring_button_1.next_flash_counter_2[11] ;
 wire \game.scoring_button_1.next_flash_counter_2[12] ;
 wire \game.scoring_button_1.next_flash_counter_2[13] ;
 wire \game.scoring_button_1.next_flash_counter_2[14] ;
 wire \game.scoring_button_1.next_flash_counter_2[15] ;
 wire \game.scoring_button_1.next_flash_counter_2[16] ;
 wire \game.scoring_button_1.next_flash_counter_2[17] ;
 wire \game.scoring_button_1.next_flash_counter_2[18] ;
 wire \game.scoring_button_1.next_flash_counter_2[19] ;
 wire \game.scoring_button_1.next_flash_counter_2[1] ;
 wire \game.scoring_button_1.next_flash_counter_2[20] ;
 wire \game.scoring_button_1.next_flash_counter_2[21] ;
 wire \game.scoring_button_1.next_flash_counter_2[22] ;
 wire \game.scoring_button_1.next_flash_counter_2[2] ;
 wire \game.scoring_button_1.next_flash_counter_2[3] ;
 wire \game.scoring_button_1.next_flash_counter_2[4] ;
 wire \game.scoring_button_1.next_flash_counter_2[5] ;
 wire \game.scoring_button_1.next_flash_counter_2[6] ;
 wire \game.scoring_button_1.next_flash_counter_2[7] ;
 wire \game.scoring_button_1.next_flash_counter_2[8] ;
 wire \game.scoring_button_1.next_flash_counter_2[9] ;
 wire \game.scoring_button_1.next_good ;
 wire \game.scoring_button_1.next_missed ;
 wire \game.scoring_button_1.next_num_hits[0] ;
 wire \game.scoring_button_1.next_num_hits[10] ;
 wire \game.scoring_button_1.next_num_hits[11] ;
 wire \game.scoring_button_1.next_num_hits[12] ;
 wire \game.scoring_button_1.next_num_hits[13] ;
 wire \game.scoring_button_1.next_num_hits[14] ;
 wire \game.scoring_button_1.next_num_hits[15] ;
 wire \game.scoring_button_1.next_num_hits[1] ;
 wire \game.scoring_button_1.next_num_hits[2] ;
 wire \game.scoring_button_1.next_num_hits[3] ;
 wire \game.scoring_button_1.next_num_hits[4] ;
 wire \game.scoring_button_1.next_num_hits[5] ;
 wire \game.scoring_button_1.next_num_hits[6] ;
 wire \game.scoring_button_1.next_num_hits[7] ;
 wire \game.scoring_button_1.next_num_hits[8] ;
 wire \game.scoring_button_1.next_num_hits[9] ;
 wire \game.scoring_button_1.next_num_misses[0] ;
 wire \game.scoring_button_1.next_num_misses[10] ;
 wire \game.scoring_button_1.next_num_misses[11] ;
 wire \game.scoring_button_1.next_num_misses[12] ;
 wire \game.scoring_button_1.next_num_misses[13] ;
 wire \game.scoring_button_1.next_num_misses[14] ;
 wire \game.scoring_button_1.next_num_misses[15] ;
 wire \game.scoring_button_1.next_num_misses[1] ;
 wire \game.scoring_button_1.next_num_misses[2] ;
 wire \game.scoring_button_1.next_num_misses[3] ;
 wire \game.scoring_button_1.next_num_misses[4] ;
 wire \game.scoring_button_1.next_num_misses[5] ;
 wire \game.scoring_button_1.next_num_misses[6] ;
 wire \game.scoring_button_1.next_num_misses[7] ;
 wire \game.scoring_button_1.next_num_misses[8] ;
 wire \game.scoring_button_1.next_num_misses[9] ;
 wire \game.scoring_button_1.next_start_count ;
 wire \game.scoring_button_2.acc[1] ;
 wire \game.scoring_button_2.acc[2] ;
 wire \game.scoring_button_2.check_hit.edge_1 ;
 wire \game.scoring_button_2.check_hit.edge_2 ;
 wire \game.scoring_button_2.check_hit.in ;
 wire \game.scoring_button_2.counts[0] ;
 wire \game.scoring_button_2.counts[10] ;
 wire \game.scoring_button_2.counts[11] ;
 wire \game.scoring_button_2.counts[12] ;
 wire \game.scoring_button_2.counts[13] ;
 wire \game.scoring_button_2.counts[14] ;
 wire \game.scoring_button_2.counts[15] ;
 wire \game.scoring_button_2.counts[16] ;
 wire \game.scoring_button_2.counts[17] ;
 wire \game.scoring_button_2.counts[18] ;
 wire \game.scoring_button_2.counts[19] ;
 wire \game.scoring_button_2.counts[1] ;
 wire \game.scoring_button_2.counts[20] ;
 wire \game.scoring_button_2.counts[21] ;
 wire \game.scoring_button_2.counts[22] ;
 wire \game.scoring_button_2.counts[2] ;
 wire \game.scoring_button_2.counts[3] ;
 wire \game.scoring_button_2.counts[4] ;
 wire \game.scoring_button_2.counts[5] ;
 wire \game.scoring_button_2.counts[6] ;
 wire \game.scoring_button_2.counts[7] ;
 wire \game.scoring_button_2.counts[8] ;
 wire \game.scoring_button_2.counts[9] ;
 wire \game.scoring_button_2.flash_counter_1[0] ;
 wire \game.scoring_button_2.flash_counter_1[10] ;
 wire \game.scoring_button_2.flash_counter_1[11] ;
 wire \game.scoring_button_2.flash_counter_1[12] ;
 wire \game.scoring_button_2.flash_counter_1[13] ;
 wire \game.scoring_button_2.flash_counter_1[14] ;
 wire \game.scoring_button_2.flash_counter_1[15] ;
 wire \game.scoring_button_2.flash_counter_1[16] ;
 wire \game.scoring_button_2.flash_counter_1[17] ;
 wire \game.scoring_button_2.flash_counter_1[18] ;
 wire \game.scoring_button_2.flash_counter_1[19] ;
 wire \game.scoring_button_2.flash_counter_1[1] ;
 wire \game.scoring_button_2.flash_counter_1[20] ;
 wire \game.scoring_button_2.flash_counter_1[21] ;
 wire \game.scoring_button_2.flash_counter_1[22] ;
 wire \game.scoring_button_2.flash_counter_1[2] ;
 wire \game.scoring_button_2.flash_counter_1[3] ;
 wire \game.scoring_button_2.flash_counter_1[4] ;
 wire \game.scoring_button_2.flash_counter_1[5] ;
 wire \game.scoring_button_2.flash_counter_1[6] ;
 wire \game.scoring_button_2.flash_counter_1[7] ;
 wire \game.scoring_button_2.flash_counter_1[8] ;
 wire \game.scoring_button_2.flash_counter_1[9] ;
 wire \game.scoring_button_2.flash_counter_2[0] ;
 wire \game.scoring_button_2.flash_counter_2[10] ;
 wire \game.scoring_button_2.flash_counter_2[11] ;
 wire \game.scoring_button_2.flash_counter_2[12] ;
 wire \game.scoring_button_2.flash_counter_2[13] ;
 wire \game.scoring_button_2.flash_counter_2[14] ;
 wire \game.scoring_button_2.flash_counter_2[15] ;
 wire \game.scoring_button_2.flash_counter_2[16] ;
 wire \game.scoring_button_2.flash_counter_2[17] ;
 wire \game.scoring_button_2.flash_counter_2[18] ;
 wire \game.scoring_button_2.flash_counter_2[19] ;
 wire \game.scoring_button_2.flash_counter_2[1] ;
 wire \game.scoring_button_2.flash_counter_2[20] ;
 wire \game.scoring_button_2.flash_counter_2[21] ;
 wire \game.scoring_button_2.flash_counter_2[22] ;
 wire \game.scoring_button_2.flash_counter_2[2] ;
 wire \game.scoring_button_2.flash_counter_2[3] ;
 wire \game.scoring_button_2.flash_counter_2[4] ;
 wire \game.scoring_button_2.flash_counter_2[5] ;
 wire \game.scoring_button_2.flash_counter_2[6] ;
 wire \game.scoring_button_2.flash_counter_2[7] ;
 wire \game.scoring_button_2.flash_counter_2[8] ;
 wire \game.scoring_button_2.flash_counter_2[9] ;
 wire \game.scoring_button_2.hit ;
 wire \game.scoring_button_2.next_count[0] ;
 wire \game.scoring_button_2.next_count[10] ;
 wire \game.scoring_button_2.next_count[11] ;
 wire \game.scoring_button_2.next_count[12] ;
 wire \game.scoring_button_2.next_count[13] ;
 wire \game.scoring_button_2.next_count[14] ;
 wire \game.scoring_button_2.next_count[15] ;
 wire \game.scoring_button_2.next_count[16] ;
 wire \game.scoring_button_2.next_count[17] ;
 wire \game.scoring_button_2.next_count[18] ;
 wire \game.scoring_button_2.next_count[19] ;
 wire \game.scoring_button_2.next_count[1] ;
 wire \game.scoring_button_2.next_count[20] ;
 wire \game.scoring_button_2.next_count[21] ;
 wire \game.scoring_button_2.next_count[22] ;
 wire \game.scoring_button_2.next_count[2] ;
 wire \game.scoring_button_2.next_count[3] ;
 wire \game.scoring_button_2.next_count[4] ;
 wire \game.scoring_button_2.next_count[5] ;
 wire \game.scoring_button_2.next_count[6] ;
 wire \game.scoring_button_2.next_count[7] ;
 wire \game.scoring_button_2.next_count[8] ;
 wire \game.scoring_button_2.next_count[9] ;
 wire \game.scoring_button_2.next_flash_counter_1[0] ;
 wire \game.scoring_button_2.next_flash_counter_1[10] ;
 wire \game.scoring_button_2.next_flash_counter_1[11] ;
 wire \game.scoring_button_2.next_flash_counter_1[12] ;
 wire \game.scoring_button_2.next_flash_counter_1[13] ;
 wire \game.scoring_button_2.next_flash_counter_1[14] ;
 wire \game.scoring_button_2.next_flash_counter_1[15] ;
 wire \game.scoring_button_2.next_flash_counter_1[16] ;
 wire \game.scoring_button_2.next_flash_counter_1[17] ;
 wire \game.scoring_button_2.next_flash_counter_1[18] ;
 wire \game.scoring_button_2.next_flash_counter_1[19] ;
 wire \game.scoring_button_2.next_flash_counter_1[1] ;
 wire \game.scoring_button_2.next_flash_counter_1[20] ;
 wire \game.scoring_button_2.next_flash_counter_1[21] ;
 wire \game.scoring_button_2.next_flash_counter_1[22] ;
 wire \game.scoring_button_2.next_flash_counter_1[2] ;
 wire \game.scoring_button_2.next_flash_counter_1[3] ;
 wire \game.scoring_button_2.next_flash_counter_1[4] ;
 wire \game.scoring_button_2.next_flash_counter_1[5] ;
 wire \game.scoring_button_2.next_flash_counter_1[6] ;
 wire \game.scoring_button_2.next_flash_counter_1[7] ;
 wire \game.scoring_button_2.next_flash_counter_1[8] ;
 wire \game.scoring_button_2.next_flash_counter_1[9] ;
 wire \game.scoring_button_2.next_flash_counter_2[0] ;
 wire \game.scoring_button_2.next_flash_counter_2[10] ;
 wire \game.scoring_button_2.next_flash_counter_2[11] ;
 wire \game.scoring_button_2.next_flash_counter_2[12] ;
 wire \game.scoring_button_2.next_flash_counter_2[13] ;
 wire \game.scoring_button_2.next_flash_counter_2[14] ;
 wire \game.scoring_button_2.next_flash_counter_2[15] ;
 wire \game.scoring_button_2.next_flash_counter_2[16] ;
 wire \game.scoring_button_2.next_flash_counter_2[17] ;
 wire \game.scoring_button_2.next_flash_counter_2[18] ;
 wire \game.scoring_button_2.next_flash_counter_2[19] ;
 wire \game.scoring_button_2.next_flash_counter_2[1] ;
 wire \game.scoring_button_2.next_flash_counter_2[20] ;
 wire \game.scoring_button_2.next_flash_counter_2[21] ;
 wire \game.scoring_button_2.next_flash_counter_2[22] ;
 wire \game.scoring_button_2.next_flash_counter_2[2] ;
 wire \game.scoring_button_2.next_flash_counter_2[3] ;
 wire \game.scoring_button_2.next_flash_counter_2[4] ;
 wire \game.scoring_button_2.next_flash_counter_2[5] ;
 wire \game.scoring_button_2.next_flash_counter_2[6] ;
 wire \game.scoring_button_2.next_flash_counter_2[7] ;
 wire \game.scoring_button_2.next_flash_counter_2[8] ;
 wire \game.scoring_button_2.next_flash_counter_2[9] ;
 wire \game.scoring_button_2.next_good ;
 wire \game.scoring_button_2.next_missed ;
 wire \game.scoring_button_2.next_num_hits[0] ;
 wire \game.scoring_button_2.next_num_hits[10] ;
 wire \game.scoring_button_2.next_num_hits[11] ;
 wire \game.scoring_button_2.next_num_hits[12] ;
 wire \game.scoring_button_2.next_num_hits[13] ;
 wire \game.scoring_button_2.next_num_hits[14] ;
 wire \game.scoring_button_2.next_num_hits[15] ;
 wire \game.scoring_button_2.next_num_hits[1] ;
 wire \game.scoring_button_2.next_num_hits[2] ;
 wire \game.scoring_button_2.next_num_hits[3] ;
 wire \game.scoring_button_2.next_num_hits[4] ;
 wire \game.scoring_button_2.next_num_hits[5] ;
 wire \game.scoring_button_2.next_num_hits[6] ;
 wire \game.scoring_button_2.next_num_hits[7] ;
 wire \game.scoring_button_2.next_num_hits[8] ;
 wire \game.scoring_button_2.next_num_hits[9] ;
 wire \game.scoring_button_2.next_num_misses[0] ;
 wire \game.scoring_button_2.next_num_misses[10] ;
 wire \game.scoring_button_2.next_num_misses[11] ;
 wire \game.scoring_button_2.next_num_misses[12] ;
 wire \game.scoring_button_2.next_num_misses[13] ;
 wire \game.scoring_button_2.next_num_misses[14] ;
 wire \game.scoring_button_2.next_num_misses[15] ;
 wire \game.scoring_button_2.next_num_misses[1] ;
 wire \game.scoring_button_2.next_num_misses[2] ;
 wire \game.scoring_button_2.next_num_misses[3] ;
 wire \game.scoring_button_2.next_num_misses[4] ;
 wire \game.scoring_button_2.next_num_misses[5] ;
 wire \game.scoring_button_2.next_num_misses[6] ;
 wire \game.scoring_button_2.next_num_misses[7] ;
 wire \game.scoring_button_2.next_num_misses[8] ;
 wire \game.scoring_button_2.next_num_misses[9] ;
 wire \game.scoring_button_2.next_start_count ;
 wire \highest_score.highest_score[0] ;
 wire \highest_score.highest_score[1] ;
 wire \highest_score.highest_score[2] ;
 wire \highest_score.highest_score[3] ;
 wire \highest_score.highest_score[4] ;
 wire \highest_score.highest_score[5] ;
 wire \highest_score.highest_score[6] ;
 wire \highest_score.highest_score[7] ;
 wire \highest_score.nxt_mode[0] ;
 wire \highest_score.nxt_mode[1] ;
 wire \highest_score.score_mode[0] ;
 wire \highest_score.score_mode[1] ;
 wire \lvls.level[0] ;
 wire \lvls.level[1] ;
 wire \lvls.level[2] ;
 wire \modetrans.mode[0] ;
 wire \modetrans.mode[1] ;
 wire \modetrans.mode[2] ;
 wire \modetrans.mode[3] ;
 wire \modetrans.mode[4] ;
 wire \modetrans.mode[5] ;
 wire \modetrans.pushed_3 ;
 wire \modetrans.pushed_4 ;
 wire \modetrans.u2.Q1 ;
 wire \modetrans.u2.Q2 ;
 wire \modetrans.u2.sync_pb ;
 wire \modetrans.u3.Q1 ;
 wire \modetrans.u3.Q2 ;
 wire \modetrans.u3.sync_pb ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \pulseout.fin_pulse[0] ;
 wire \pulseout.fin_pulse[1] ;
 wire \pulseout.fin_pulse[2] ;
 wire \pulseout.fin_pulse[3] ;
 wire \pulseout.fin_pulse[4] ;
 wire \pulseout.fin_pulse[5] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net29));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_99 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__buf_6 _2680_ (.A(\modetrans.mode[2] ),
    .X(_2654_));
 sky130_fd_sc_hd__nand2b_4 _2681_ (.A_N(net148),
    .B(\disp_song.um.boton1e.edge_1 ),
    .Y(_2655_));
 sky130_fd_sc_hd__nor2b_4 _2682_ (.A(\disp_song.um.boton0e.edge_2 ),
    .B_N(\disp_song.um.boton0e.edge_1 ),
    .Y(_2656_));
 sky130_fd_sc_hd__nor2_4 _2683_ (.A(_2655_),
    .B(_2656_),
    .Y(_2657_));
 sky130_fd_sc_hd__nor2b_4 _2684_ (.A(net148),
    .B_N(\disp_song.um.boton1e.edge_1 ),
    .Y(_2658_));
 sky130_fd_sc_hd__or2b_4 _2685_ (.A(\disp_song.um.boton0e.edge_2 ),
    .B_N(\disp_song.um.boton0e.edge_1 ),
    .X(_2659_));
 sky130_fd_sc_hd__nor2_4 _2686_ (.A(_2658_),
    .B(_2659_),
    .Y(_2660_));
 sky130_fd_sc_hd__clkbuf_8 _2687_ (.A(\disp_song.toggle_state ),
    .X(_2661_));
 sky130_fd_sc_hd__o21ai_4 _2688_ (.A1(_2657_),
    .A2(_2660_),
    .B1(_2661_),
    .Y(_2662_));
 sky130_fd_sc_hd__or2_1 _2689_ (.A(\disp_song.um.idx_note2[0] ),
    .B(_2662_),
    .X(_2663_));
 sky130_fd_sc_hd__xor2_2 _2690_ (.A(\disp_song.um.idx_note2[1] ),
    .B(_2663_),
    .X(_2664_));
 sky130_fd_sc_hd__and2_1 _2691_ (.A(_2654_),
    .B(_2664_),
    .X(_2665_));
 sky130_fd_sc_hd__clkbuf_8 _2692_ (.A(_2665_),
    .X(_2666_));
 sky130_fd_sc_hd__inv_2 _2693_ (.A(_2666_),
    .Y(_2667_));
 sky130_fd_sc_hd__clkbuf_8 _2694_ (.A(_2667_),
    .X(\disp_song.um.drum.next_idx2[1] ));
 sky130_fd_sc_hd__nand2_1 _2695_ (.A(_2654_),
    .B(_2663_),
    .Y(_2668_));
 sky130_fd_sc_hd__a21oi_4 _2696_ (.A1(\disp_song.um.idx_note2[0] ),
    .A2(_2662_),
    .B1(_2668_),
    .Y(_2669_));
 sky130_fd_sc_hd__inv_2 _2697_ (.A(_2669_),
    .Y(_2670_));
 sky130_fd_sc_hd__clkbuf_8 _2698_ (.A(_2670_),
    .X(\disp_song.um.drum.next_idx2[0] ));
 sky130_fd_sc_hd__inv_2 _2699_ (.A(\disp_song.um.idx_note2[3] ),
    .Y(_2671_));
 sky130_fd_sc_hd__or3_2 _2700_ (.A(\disp_song.um.idx_note2[1] ),
    .B(\disp_song.um.idx_note2[0] ),
    .C(\disp_song.um.idx_note2[2] ),
    .X(_2672_));
 sky130_fd_sc_hd__nor2_1 _2701_ (.A(\disp_song.um.idx_note2[3] ),
    .B(_2672_),
    .Y(_2673_));
 sky130_fd_sc_hd__and2_1 _2702_ (.A(\disp_song.um.idx_note2[3] ),
    .B(_2672_),
    .X(_2674_));
 sky130_fd_sc_hd__nor2_1 _2703_ (.A(_2673_),
    .B(_2674_),
    .Y(_2675_));
 sky130_fd_sc_hd__o21a_1 _2704_ (.A1(_2657_),
    .A2(_2660_),
    .B1(_2661_),
    .X(_2676_));
 sky130_fd_sc_hd__mux2_2 _2705_ (.A0(_2671_),
    .A1(_2675_),
    .S(_2676_),
    .X(_2677_));
 sky130_fd_sc_hd__and2_1 _2706_ (.A(_2654_),
    .B(_2677_),
    .X(_2678_));
 sky130_fd_sc_hd__clkbuf_4 _2707_ (.A(_2678_),
    .X(_2679_));
 sky130_fd_sc_hd__inv_2 _2708_ (.A(_2679_),
    .Y(\disp_song.um.drum.next_idx2[3] ));
 sky130_fd_sc_hd__inv_2 _2709_ (.A(\disp_song.um.idx_note2[4] ),
    .Y(_0156_));
 sky130_fd_sc_hd__or2_1 _2710_ (.A(\disp_song.um.idx_note2[3] ),
    .B(_2672_),
    .X(_0157_));
 sky130_fd_sc_hd__nor2_2 _2711_ (.A(\disp_song.um.idx_note2[4] ),
    .B(_0157_),
    .Y(_0158_));
 sky130_fd_sc_hd__nor2_1 _2712_ (.A(_0156_),
    .B(_2673_),
    .Y(_0159_));
 sky130_fd_sc_hd__nor2_1 _2713_ (.A(_0158_),
    .B(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__and3_1 _2714_ (.A(_2654_),
    .B(_2676_),
    .C(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__a31o_4 _2715_ (.A1(_2654_),
    .A2(_0156_),
    .A3(_2662_),
    .B1(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__inv_2 _2716_ (.A(_0162_),
    .Y(\disp_song.um.drum.next_idx2[4] ));
 sky130_fd_sc_hd__or3b_4 _2717_ (.A(\disp_song.um.idx_note2[1] ),
    .B(\disp_song.um.idx_note2[0] ),
    .C_N(\disp_song.um.idx_note2[2] ),
    .X(_0163_));
 sky130_fd_sc_hd__inv_2 _2718_ (.A(_0163_),
    .Y(_0164_));
 sky130_fd_sc_hd__o21ba_1 _2719_ (.A1(\disp_song.um.idx_note2[1] ),
    .A2(\disp_song.um.idx_note2[0] ),
    .B1_N(\disp_song.um.idx_note2[2] ),
    .X(_0165_));
 sky130_fd_sc_hd__or2_2 _2720_ (.A(_0164_),
    .B(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__nand2_1 _2721_ (.A(\disp_song.um.idx_note2[2] ),
    .B(_2662_),
    .Y(_0167_));
 sky130_fd_sc_hd__o211a_1 _2722_ (.A1(_2662_),
    .A2(_0166_),
    .B1(_0167_),
    .C1(_2654_),
    .X(_0168_));
 sky130_fd_sc_hd__clkbuf_8 _2723_ (.A(_0168_),
    .X(_0169_));
 sky130_fd_sc_hd__inv_4 _2724_ (.A(_0169_),
    .Y(\disp_song.um.drum.next_idx2[2] ));
 sky130_fd_sc_hd__o21bai_4 _2725_ (.A1(_2657_),
    .A2(_2660_),
    .B1_N(\disp_song.toggle_state ),
    .Y(_0170_));
 sky130_fd_sc_hd__nor2_1 _2726_ (.A(\disp_song.um.idx_note1[0] ),
    .B(_0170_),
    .Y(_0171_));
 sky130_fd_sc_hd__and2_1 _2727_ (.A(\disp_song.um.idx_note1[0] ),
    .B(_0170_),
    .X(_0172_));
 sky130_fd_sc_hd__nor2_1 _2728_ (.A(_0171_),
    .B(_0172_),
    .Y(_0173_));
 sky130_fd_sc_hd__and2_1 _2729_ (.A(_2654_),
    .B(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__buf_4 _2730_ (.A(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__inv_2 _2731_ (.A(_0175_),
    .Y(_0176_));
 sky130_fd_sc_hd__clkbuf_8 _2732_ (.A(_0176_),
    .X(\disp_song.um.drum.next_idx1[0] ));
 sky130_fd_sc_hd__inv_2 _2733_ (.A(\disp_song.um.idx_note1[3] ),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _2734_ (.A(\disp_song.um.idx_note1[2] ),
    .Y(_0178_));
 sky130_fd_sc_hd__clkbuf_8 _2735_ (.A(\disp_song.um.idx_note1[1] ),
    .X(_0179_));
 sky130_fd_sc_hd__nor2_2 _2736_ (.A(\disp_song.um.idx_note1[0] ),
    .B(_0179_),
    .Y(_0180_));
 sky130_fd_sc_hd__and2_1 _2737_ (.A(_0178_),
    .B(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__nand2_1 _2738_ (.A(_0177_),
    .B(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__or2_1 _2739_ (.A(\disp_song.um.idx_note1[4] ),
    .B(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__o21ai_1 _2740_ (.A1(_0170_),
    .A2(_0182_),
    .B1(\disp_song.um.idx_note1[4] ),
    .Y(_0184_));
 sky130_fd_sc_hd__o211a_4 _2741_ (.A1(_0170_),
    .A2(_0183_),
    .B1(_0184_),
    .C1(_2654_),
    .X(_0185_));
 sky130_fd_sc_hd__inv_2 _2742_ (.A(_0185_),
    .Y(\disp_song.um.drum.next_idx1[4] ));
 sky130_fd_sc_hd__nand2_1 _2743_ (.A(_0178_),
    .B(_0180_),
    .Y(_0186_));
 sky130_fd_sc_hd__or2_1 _2744_ (.A(_0178_),
    .B(_0180_),
    .X(_0187_));
 sky130_fd_sc_hd__a21oi_1 _2745_ (.A1(_0186_),
    .A2(_0187_),
    .B1(_0170_),
    .Y(_0188_));
 sky130_fd_sc_hd__a21oi_1 _2746_ (.A1(\disp_song.um.idx_note1[2] ),
    .A2(_0170_),
    .B1(_0188_),
    .Y(_0189_));
 sky130_fd_sc_hd__and2_1 _2747_ (.A(_2654_),
    .B(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__buf_4 _2748_ (.A(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__clkinv_4 _2749_ (.A(_0191_),
    .Y(\disp_song.um.drum.next_idx1[2] ));
 sky130_fd_sc_hd__nand2_1 _2750_ (.A(\disp_song.um.idx_note1[3] ),
    .B(_0186_),
    .Y(_0192_));
 sky130_fd_sc_hd__and2_1 _2751_ (.A(_0182_),
    .B(_0192_),
    .X(_0193_));
 sky130_fd_sc_hd__buf_2 _2752_ (.A(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _2753_ (.A0(_0194_),
    .A1(_0177_),
    .S(_0170_),
    .X(_0195_));
 sky130_fd_sc_hd__and2_1 _2754_ (.A(\modetrans.mode[2] ),
    .B(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__buf_4 _2755_ (.A(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__inv_2 _2756_ (.A(_0197_),
    .Y(\disp_song.um.drum.next_idx1[3] ));
 sky130_fd_sc_hd__xnor2_2 _2757_ (.A(_0179_),
    .B(_0171_),
    .Y(_0198_));
 sky130_fd_sc_hd__and2_2 _2758_ (.A(_2654_),
    .B(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__inv_6 _2759_ (.A(_0199_),
    .Y(\disp_song.um.drum.next_idx1[1] ));
 sky130_fd_sc_hd__and2_1 _2760_ (.A(\modetrans.mode[5] ),
    .B(_2658_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _2761_ (.A0(\lvls.level[0] ),
    .A1(\lvls.level[2] ),
    .S(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__clkbuf_1 _2762_ (.A(_0201_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _2763_ (.A0(\lvls.level[2] ),
    .A1(\lvls.level[1] ),
    .S(_0200_),
    .X(_0202_));
 sky130_fd_sc_hd__clkbuf_1 _2764_ (.A(_0202_),
    .X(_0002_));
 sky130_fd_sc_hd__and2b_1 _2765_ (.A_N(\modetrans.u3.Q2 ),
    .B(\modetrans.u3.Q1 ),
    .X(_0203_));
 sky130_fd_sc_hd__inv_2 _2766_ (.A(\pulseout.fin_pulse[5] ),
    .Y(_0204_));
 sky130_fd_sc_hd__or3b_1 _2767_ (.A(\pulseout.fin_pulse[2] ),
    .B(\pulseout.fin_pulse[4] ),
    .C_N(\pulseout.fin_pulse[3] ),
    .X(_0205_));
 sky130_fd_sc_hd__or4b_4 _2768_ (.A(\pulseout.fin_pulse[1] ),
    .B(_0204_),
    .C(_0205_),
    .D_N(\pulseout.fin_pulse[0] ),
    .X(_0206_));
 sky130_fd_sc_hd__nor2_1 _2769_ (.A(_0203_),
    .B(_0206_),
    .Y(_0207_));
 sky130_fd_sc_hd__clkbuf_16 _2770_ (.A(\modetrans.mode[0] ),
    .X(_0208_));
 sky130_fd_sc_hd__buf_8 _2771_ (.A(\modetrans.mode[1] ),
    .X(_0209_));
 sky130_fd_sc_hd__or2_4 _2772_ (.A(_0209_),
    .B(\modetrans.mode[4] ),
    .X(_0210_));
 sky130_fd_sc_hd__buf_8 _2773_ (.A(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__o31a_1 _2774_ (.A1(\modetrans.mode[5] ),
    .A2(_0208_),
    .A3(_0211_),
    .B1(_0203_),
    .X(_0212_));
 sky130_fd_sc_hd__or2b_1 _2775_ (.A(net114),
    .B_N(\modetrans.u2.Q1 ),
    .X(_0213_));
 sky130_fd_sc_hd__o31a_1 _2776_ (.A1(\modetrans.mode[3] ),
    .A2(_0207_),
    .A3(_0212_),
    .B1(_0213_),
    .X(_0006_));
 sky130_fd_sc_hd__buf_6 _2777_ (.A(_2654_),
    .X(_0214_));
 sky130_fd_sc_hd__nand2_1 _2778_ (.A(_0214_),
    .B(_0213_),
    .Y(_0215_));
 sky130_fd_sc_hd__and2b_1 _2779_ (.A_N(\modetrans.u2.Q2 ),
    .B(\modetrans.u2.Q1 ),
    .X(_0216_));
 sky130_fd_sc_hd__clkbuf_2 _2780_ (.A(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__a2bb2o_1 _2781_ (.A1_N(_0207_),
    .A2_N(_0215_),
    .B1(_0208_),
    .B2(_0217_),
    .X(_0005_));
 sky130_fd_sc_hd__nor3b_2 _2782_ (.A(_0217_),
    .B(_0203_),
    .C_N(_0206_),
    .Y(_0218_));
 sky130_fd_sc_hd__a22o_1 _2783_ (.A1(_0214_),
    .A2(_0217_),
    .B1(_0218_),
    .B2(\modetrans.mode[5] ),
    .X(_0008_));
 sky130_fd_sc_hd__buf_8 _2784_ (.A(_0209_),
    .X(_0219_));
 sky130_fd_sc_hd__or2_1 _2785_ (.A(\modetrans.mode[5] ),
    .B(net270),
    .X(_0220_));
 sky130_fd_sc_hd__a22o_1 _2786_ (.A1(_0219_),
    .A2(_0218_),
    .B1(_0220_),
    .B2(_0217_),
    .X(_0004_));
 sky130_fd_sc_hd__a22o_1 _2787_ (.A1(\modetrans.mode[3] ),
    .A2(_0217_),
    .B1(_0218_),
    .B2(_0208_),
    .X(_0003_));
 sky130_fd_sc_hd__a22o_1 _2788_ (.A1(_0219_),
    .A2(_0217_),
    .B1(_0218_),
    .B2(net164),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _2789_ (.A0(\lvls.level[1] ),
    .A1(\lvls.level[0] ),
    .S(_0200_),
    .X(_0221_));
 sky130_fd_sc_hd__clkbuf_1 _2790_ (.A(_0221_),
    .X(_0001_));
 sky130_fd_sc_hd__nor2b_2 _2791_ (.A(\lvls.level[0] ),
    .B_N(\lvls.level[1] ),
    .Y(_0222_));
 sky130_fd_sc_hd__nand2_1 _2792_ (.A(\game.counter[20] ),
    .B(_0222_),
    .Y(_0223_));
 sky130_fd_sc_hd__or2_1 _2793_ (.A(\game.counter[20] ),
    .B(_0222_),
    .X(_0224_));
 sky130_fd_sc_hd__o21a_1 _2794_ (.A1(\game.counter[14] ),
    .A2(_0223_),
    .B1(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__or3b_1 _2795_ (.A(\lvls.level[0] ),
    .B(\lvls.level[1] ),
    .C_N(\lvls.level[2] ),
    .X(_0226_));
 sky130_fd_sc_hd__clkbuf_4 _2796_ (.A(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__xor2_1 _2797_ (.A(\game.counter[11] ),
    .B(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__xor2_1 _2798_ (.A(\game.counter[8] ),
    .B(_0227_),
    .X(_0229_));
 sky130_fd_sc_hd__xor2_1 _2799_ (.A(\game.counter[10] ),
    .B(_0227_),
    .X(_0230_));
 sky130_fd_sc_hd__or4b_1 _2800_ (.A(_0225_),
    .B(_0228_),
    .C(_0229_),
    .D_N(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__clkbuf_2 _2801_ (.A(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__nor2_1 _2802_ (.A(\game.counter[6] ),
    .B(_0222_),
    .Y(_0233_));
 sky130_fd_sc_hd__and2_1 _2803_ (.A(\game.counter[6] ),
    .B(_0222_),
    .X(_0234_));
 sky130_fd_sc_hd__xnor2_1 _2804_ (.A(\game.counter[7] ),
    .B(_0227_),
    .Y(_0235_));
 sky130_fd_sc_hd__or3_1 _2805_ (.A(_0233_),
    .B(_0234_),
    .C(_0235_),
    .X(_0236_));
 sky130_fd_sc_hd__inv_2 _2806_ (.A(\game.counter[14] ),
    .Y(_0237_));
 sky130_fd_sc_hd__or4b_1 _2807_ (.A(\game.counter[5] ),
    .B(\game.counter[13] ),
    .C(\game.counter[12] ),
    .D_N(_0209_),
    .X(_0238_));
 sky130_fd_sc_hd__a221o_1 _2808_ (.A1(\game.counter[9] ),
    .A2(_0237_),
    .B1(\game.counter[15] ),
    .B2(_0227_),
    .C1(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__inv_2 _2809_ (.A(\game.counter[15] ),
    .Y(_0240_));
 sky130_fd_sc_hd__inv_2 _2810_ (.A(_0227_),
    .Y(_0241_));
 sky130_fd_sc_hd__nor2_1 _2811_ (.A(\lvls.level[2] ),
    .B(\lvls.level[1] ),
    .Y(_0242_));
 sky130_fd_sc_hd__or2_1 _2812_ (.A(\lvls.level[0] ),
    .B(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__a22o_1 _2813_ (.A1(_0240_),
    .A2(_0241_),
    .B1(_0243_),
    .B2(\game.counter[21] ),
    .X(_0244_));
 sky130_fd_sc_hd__nor2_1 _2814_ (.A(\lvls.level[0] ),
    .B(_0242_),
    .Y(_0245_));
 sky130_fd_sc_hd__o21a_1 _2815_ (.A1(\game.counter[16] ),
    .A2(_0245_),
    .B1(\game.counter[22] ),
    .X(_0246_));
 sky130_fd_sc_hd__a21oi_1 _2816_ (.A1(\game.counter[16] ),
    .A2(\game.counter[21] ),
    .B1(\game.counter[22] ),
    .Y(_0247_));
 sky130_fd_sc_hd__or2_1 _2817_ (.A(\game.counter[1] ),
    .B(\game.counter[0] ),
    .X(_0248_));
 sky130_fd_sc_hd__or3_1 _2818_ (.A(\game.counter[3] ),
    .B(\game.counter[2] ),
    .C(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__nor2_1 _2819_ (.A(\game.counter[4] ),
    .B(\game.counter[17] ),
    .Y(_0250_));
 sky130_fd_sc_hd__o2111a_1 _2820_ (.A1(\game.counter[9] ),
    .A2(_0222_),
    .B1(_0250_),
    .C1(\game.counter[19] ),
    .D1(\game.counter[18] ),
    .X(_0251_));
 sky130_fd_sc_hd__or4b_1 _2821_ (.A(_0246_),
    .B(_0247_),
    .C(_0249_),
    .D_N(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__or4_1 _2822_ (.A(_0236_),
    .B(_0239_),
    .C(_0244_),
    .D(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__clkbuf_2 _2823_ (.A(_0253_),
    .X(_0254_));
 sky130_fd_sc_hd__nor2_4 _2824_ (.A(_0232_),
    .B(_0254_),
    .Y(_0032_));
 sky130_fd_sc_hd__clkbuf_8 _2825_ (.A(\highest_score.score_mode[0] ),
    .X(_0255_));
 sky130_fd_sc_hd__nand2_1 _2826_ (.A(_0255_),
    .B(_2659_),
    .Y(_0256_));
 sky130_fd_sc_hd__or2_1 _2827_ (.A(_0255_),
    .B(_2659_),
    .X(_0257_));
 sky130_fd_sc_hd__nand2_1 _2828_ (.A(_0256_),
    .B(_0257_),
    .Y(\highest_score.nxt_mode[0] ));
 sky130_fd_sc_hd__clkbuf_8 _2829_ (.A(\highest_score.score_mode[1] ),
    .X(_0258_));
 sky130_fd_sc_hd__nor2_4 _2830_ (.A(_0255_),
    .B(_0258_),
    .Y(_0259_));
 sky130_fd_sc_hd__and2_1 _2831_ (.A(_0255_),
    .B(_0258_),
    .X(_0260_));
 sky130_fd_sc_hd__buf_2 _2832_ (.A(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__nor2_1 _2833_ (.A(_0259_),
    .B(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__xnor2_1 _2834_ (.A(_0256_),
    .B(_0262_),
    .Y(\highest_score.nxt_mode[1] ));
 sky130_fd_sc_hd__and3_1 _2835_ (.A(\modetrans.mode[2] ),
    .B(_2658_),
    .C(_2659_),
    .X(_0263_));
 sky130_fd_sc_hd__buf_2 _2836_ (.A(_0263_),
    .X(_0264_));
 sky130_fd_sc_hd__nand2_2 _2837_ (.A(_2654_),
    .B(_2660_),
    .Y(_0265_));
 sky130_fd_sc_hd__nand2_1 _2838_ (.A(_2661_),
    .B(_0158_),
    .Y(_0266_));
 sky130_fd_sc_hd__o21a_1 _2839_ (.A1(_0265_),
    .A2(_0266_),
    .B1(\disp_song.note2[0] ),
    .X(_0267_));
 sky130_fd_sc_hd__a31o_1 _2840_ (.A1(_2661_),
    .A2(_0158_),
    .A3(_0264_),
    .B1(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2841_ (.A(_0268_),
    .X(\disp_song.um.drum.next_note2[0] ));
 sky130_fd_sc_hd__clkbuf_8 _2842_ (.A(_2657_),
    .X(_0269_));
 sky130_fd_sc_hd__or3b_2 _2843_ (.A(\disp_song.um.idx_note2[1] ),
    .B(\disp_song.um.idx_note2[2] ),
    .C_N(\disp_song.um.idx_note2[0] ),
    .X(_0270_));
 sky130_fd_sc_hd__inv_2 _2844_ (.A(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__and4_1 _2845_ (.A(_2654_),
    .B(_0156_),
    .C(_2676_),
    .D(_2675_),
    .X(_0272_));
 sky130_fd_sc_hd__clkbuf_2 _2846_ (.A(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__nand2_1 _2847_ (.A(_0271_),
    .B(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__mux2_1 _2848_ (.A0(_0269_),
    .A1(\disp_song.note2[1] ),
    .S(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__buf_1 _2849_ (.A(_0275_),
    .X(\disp_song.um.drum.next_note2[1] ));
 sky130_fd_sc_hd__or3b_2 _2850_ (.A(\disp_song.um.idx_note2[0] ),
    .B(\disp_song.um.idx_note2[2] ),
    .C_N(\disp_song.um.idx_note2[1] ),
    .X(_0276_));
 sky130_fd_sc_hd__or3b_1 _2851_ (.A(_0276_),
    .B(\disp_song.um.idx_note2[3] ),
    .C_N(_0161_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _2852_ (.A0(_0269_),
    .A1(\disp_song.note2[2] ),
    .S(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__buf_1 _2853_ (.A(_0278_),
    .X(\disp_song.um.drum.next_note2[2] ));
 sky130_fd_sc_hd__nand3_2 _2854_ (.A(\disp_song.um.idx_note2[1] ),
    .B(\disp_song.um.idx_note2[0] ),
    .C(_0166_),
    .Y(_0279_));
 sky130_fd_sc_hd__or3b_1 _2855_ (.A(_0279_),
    .B(\disp_song.um.idx_note2[3] ),
    .C_N(_0161_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _2856_ (.A0(_0269_),
    .A1(\disp_song.note2[3] ),
    .S(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__buf_1 _2857_ (.A(_0281_),
    .X(\disp_song.um.drum.next_note2[3] ));
 sky130_fd_sc_hd__or3b_1 _2858_ (.A(\disp_song.um.idx_note2[3] ),
    .B(\disp_song.um.idx_note2[4] ),
    .C_N(_2661_),
    .X(_0282_));
 sky130_fd_sc_hd__nor2_1 _2859_ (.A(_0163_),
    .B(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__or3_1 _2860_ (.A(_0163_),
    .B(_0265_),
    .C(_0282_),
    .X(_0284_));
 sky130_fd_sc_hd__a22o_1 _2861_ (.A1(_0264_),
    .A2(_0283_),
    .B1(_0284_),
    .B2(\disp_song.note2[4] ),
    .X(\disp_song.um.drum.next_note2[4] ));
 sky130_fd_sc_hd__and3b_1 _2862_ (.A_N(\disp_song.um.idx_note2[1] ),
    .B(\disp_song.um.idx_note2[0] ),
    .C(\disp_song.um.idx_note2[2] ),
    .X(_0285_));
 sky130_fd_sc_hd__nand2_1 _2863_ (.A(_0273_),
    .B(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__mux2_1 _2864_ (.A0(_0269_),
    .A1(\disp_song.note2[5] ),
    .S(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__buf_1 _2865_ (.A(_0287_),
    .X(\disp_song.um.drum.next_note2[5] ));
 sky130_fd_sc_hd__and3b_1 _2866_ (.A_N(\disp_song.um.idx_note2[0] ),
    .B(\disp_song.um.idx_note2[2] ),
    .C(\disp_song.um.idx_note2[1] ),
    .X(_0288_));
 sky130_fd_sc_hd__nand2_1 _2867_ (.A(_0273_),
    .B(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__mux2_1 _2868_ (.A0(_0269_),
    .A1(\disp_song.note2[6] ),
    .S(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__buf_1 _2869_ (.A(_0290_),
    .X(\disp_song.um.drum.next_note2[6] ));
 sky130_fd_sc_hd__and3_1 _2870_ (.A(\disp_song.um.idx_note2[1] ),
    .B(\disp_song.um.idx_note2[0] ),
    .C(\disp_song.um.idx_note2[2] ),
    .X(_0291_));
 sky130_fd_sc_hd__nand2_1 _2871_ (.A(_0273_),
    .B(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__mux2_1 _2872_ (.A0(_0269_),
    .A1(\disp_song.note2[7] ),
    .S(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__buf_1 _2873_ (.A(_0293_),
    .X(\disp_song.um.drum.next_note2[7] ));
 sky130_fd_sc_hd__nor2_1 _2874_ (.A(_2672_),
    .B(_0158_),
    .Y(_0294_));
 sky130_fd_sc_hd__nand2_1 _2875_ (.A(_0273_),
    .B(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__mux2_1 _2876_ (.A0(_0269_),
    .A1(\disp_song.note2[8] ),
    .S(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__clkbuf_1 _2877_ (.A(_0296_),
    .X(\disp_song.um.drum.next_note2[8] ));
 sky130_fd_sc_hd__or2_1 _2878_ (.A(_2673_),
    .B(_2674_),
    .X(_0297_));
 sky130_fd_sc_hd__nand2_2 _2879_ (.A(_0297_),
    .B(_0161_),
    .Y(_0298_));
 sky130_fd_sc_hd__nor2_1 _2880_ (.A(_0270_),
    .B(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__mux2_1 _2881_ (.A0(\disp_song.note2[9] ),
    .A1(_0269_),
    .S(_0299_),
    .X(_0300_));
 sky130_fd_sc_hd__buf_1 _2882_ (.A(_0300_),
    .X(\disp_song.um.drum.next_note2[9] ));
 sky130_fd_sc_hd__nor2_1 _2883_ (.A(_0276_),
    .B(_0298_),
    .Y(_0301_));
 sky130_fd_sc_hd__mux2_1 _2884_ (.A0(\disp_song.note2[10] ),
    .A1(_0269_),
    .S(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__buf_1 _2885_ (.A(_0302_),
    .X(\disp_song.um.drum.next_note2[10] ));
 sky130_fd_sc_hd__nor2_1 _2886_ (.A(_0279_),
    .B(_0298_),
    .Y(_0303_));
 sky130_fd_sc_hd__mux2_1 _2887_ (.A0(\disp_song.note2[11] ),
    .A1(_0269_),
    .S(_0303_),
    .X(_0304_));
 sky130_fd_sc_hd__buf_1 _2888_ (.A(_0304_),
    .X(\disp_song.um.drum.next_note2[11] ));
 sky130_fd_sc_hd__nor2_1 _2889_ (.A(_0163_),
    .B(_0298_),
    .Y(_0305_));
 sky130_fd_sc_hd__mux2_1 _2890_ (.A0(\disp_song.note2[12] ),
    .A1(_0269_),
    .S(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__buf_1 _2891_ (.A(_0306_),
    .X(\disp_song.um.drum.next_note2[12] ));
 sky130_fd_sc_hd__or3b_1 _2892_ (.A(_0166_),
    .B(\disp_song.um.idx_note2[1] ),
    .C_N(\disp_song.um.idx_note2[0] ),
    .X(_0307_));
 sky130_fd_sc_hd__nor2_1 _2893_ (.A(_0307_),
    .B(_0298_),
    .Y(_0308_));
 sky130_fd_sc_hd__mux2_1 _2894_ (.A0(\disp_song.note2[13] ),
    .A1(_0269_),
    .S(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__buf_1 _2895_ (.A(_0309_),
    .X(\disp_song.um.drum.next_note2[13] ));
 sky130_fd_sc_hd__or3b_1 _2896_ (.A(\disp_song.um.idx_note2[0] ),
    .B(_0166_),
    .C_N(\disp_song.um.idx_note2[1] ),
    .X(_0310_));
 sky130_fd_sc_hd__nor2_1 _2897_ (.A(_0310_),
    .B(_0298_),
    .Y(_0311_));
 sky130_fd_sc_hd__mux2_1 _2898_ (.A0(\disp_song.note2[14] ),
    .A1(_0269_),
    .S(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__buf_1 _2899_ (.A(_0312_),
    .X(\disp_song.um.drum.next_note2[14] ));
 sky130_fd_sc_hd__nand3_1 _2900_ (.A(\disp_song.um.idx_note2[1] ),
    .B(\disp_song.um.idx_note2[0] ),
    .C(\disp_song.um.idx_note2[2] ),
    .Y(_0313_));
 sky130_fd_sc_hd__nor2_1 _2901_ (.A(_0313_),
    .B(_0298_),
    .Y(_0314_));
 sky130_fd_sc_hd__mux2_1 _2902_ (.A0(\disp_song.note2[15] ),
    .A1(_2657_),
    .S(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__buf_1 _2903_ (.A(_0315_),
    .X(\disp_song.um.drum.next_note2[15] ));
 sky130_fd_sc_hd__nand2_1 _2904_ (.A(_2661_),
    .B(\disp_song.um.idx_note2[4] ),
    .Y(_0316_));
 sky130_fd_sc_hd__o31a_1 _2905_ (.A1(_0157_),
    .A2(_0265_),
    .A3(_0316_),
    .B1(\disp_song.note2[16] ),
    .X(_0317_));
 sky130_fd_sc_hd__a41o_1 _2906_ (.A1(_2661_),
    .A2(\disp_song.um.idx_note2[4] ),
    .A3(_2673_),
    .A4(_0264_),
    .B1(_0317_),
    .X(\disp_song.um.drum.next_note2[16] ));
 sky130_fd_sc_hd__nand2_1 _2907_ (.A(_2654_),
    .B(_2676_),
    .Y(_0318_));
 sky130_fd_sc_hd__or4_1 _2908_ (.A(_0156_),
    .B(_0297_),
    .C(_0318_),
    .D(_0270_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _2909_ (.A0(_2657_),
    .A1(\disp_song.note2[17] ),
    .S(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__clkbuf_1 _2910_ (.A(_0320_),
    .X(\disp_song.um.drum.next_note2[17] ));
 sky130_fd_sc_hd__or4_1 _2911_ (.A(\disp_song.um.idx_note2[3] ),
    .B(_0318_),
    .C(_0160_),
    .D(_0276_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _2912_ (.A0(_0269_),
    .A1(\disp_song.note2[18] ),
    .S(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__buf_1 _2913_ (.A(_0322_),
    .X(\disp_song.um.drum.next_note2[18] ));
 sky130_fd_sc_hd__or4_1 _2914_ (.A(\disp_song.um.idx_note2[3] ),
    .B(_0318_),
    .C(_0160_),
    .D(_0279_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _2915_ (.A0(_0269_),
    .A1(\disp_song.note2[19] ),
    .S(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__buf_1 _2916_ (.A(_0324_),
    .X(\disp_song.um.drum.next_note2[19] ));
 sky130_fd_sc_hd__nand2_2 _2917_ (.A(_2661_),
    .B(\modetrans.mode[2] ),
    .Y(_0325_));
 sky130_fd_sc_hd__nor2_1 _2918_ (.A(_0160_),
    .B(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__inv_2 _2919_ (.A(_0325_),
    .Y(\disp_song.next_red ));
 sky130_fd_sc_hd__nand4_2 _2920_ (.A(\disp_song.um.idx_note2[4] ),
    .B(_2660_),
    .C(_2675_),
    .D(\disp_song.next_red ),
    .Y(_0327_));
 sky130_fd_sc_hd__o21a_1 _2921_ (.A1(_0163_),
    .A2(_0327_),
    .B1(\disp_song.note2[20] ),
    .X(_0328_));
 sky130_fd_sc_hd__a41o_1 _2922_ (.A1(_2671_),
    .A2(_0269_),
    .A3(_0164_),
    .A4(_0326_),
    .B1(_0328_),
    .X(\disp_song.um.drum.next_note2[20] ));
 sky130_fd_sc_hd__or2_1 _2923_ (.A(_0307_),
    .B(_0327_),
    .X(_0329_));
 sky130_fd_sc_hd__and4_2 _2924_ (.A(\disp_song.um.idx_note2[4] ),
    .B(_0269_),
    .C(_2675_),
    .D(\disp_song.next_red ),
    .X(_0330_));
 sky130_fd_sc_hd__a22o_1 _2925_ (.A1(\disp_song.note2[21] ),
    .A2(_0329_),
    .B1(_0330_),
    .B2(_0285_),
    .X(\disp_song.um.drum.next_note2[21] ));
 sky130_fd_sc_hd__or2_1 _2926_ (.A(_0310_),
    .B(_0327_),
    .X(_0331_));
 sky130_fd_sc_hd__a22o_1 _2927_ (.A1(_0288_),
    .A2(_0330_),
    .B1(_0331_),
    .B2(net191),
    .X(\disp_song.um.drum.next_note2[22] ));
 sky130_fd_sc_hd__or2_1 _2928_ (.A(_0313_),
    .B(_0327_),
    .X(_0332_));
 sky130_fd_sc_hd__a22o_1 _2929_ (.A1(_0291_),
    .A2(_0330_),
    .B1(_0332_),
    .B2(net236),
    .X(\disp_song.um.drum.next_note2[23] ));
 sky130_fd_sc_hd__or3_1 _2930_ (.A(_2672_),
    .B(_0158_),
    .C(_0327_),
    .X(_0333_));
 sky130_fd_sc_hd__a22o_1 _2931_ (.A1(_0294_),
    .A2(_0330_),
    .B1(_0333_),
    .B2(\disp_song.note2[24] ),
    .X(\disp_song.um.drum.next_note2[24] ));
 sky130_fd_sc_hd__and3_1 _2932_ (.A(\disp_song.um.idx_note2[3] ),
    .B(\disp_song.um.idx_note2[4] ),
    .C(\disp_song.next_red ),
    .X(_0334_));
 sky130_fd_sc_hd__nand2_1 _2933_ (.A(_0297_),
    .B(_0326_),
    .Y(_0335_));
 sky130_fd_sc_hd__or2_1 _2934_ (.A(_2659_),
    .B(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__or2_2 _2935_ (.A(_2658_),
    .B(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__o21a_1 _2936_ (.A1(_0270_),
    .A2(_0337_),
    .B1(\disp_song.note2[25] ),
    .X(_0338_));
 sky130_fd_sc_hd__a31o_1 _2937_ (.A1(_0269_),
    .A2(_0271_),
    .A3(_0334_),
    .B1(_0338_),
    .X(\disp_song.um.drum.next_note2[25] ));
 sky130_fd_sc_hd__or2_1 _2938_ (.A(_2656_),
    .B(_0335_),
    .X(_0339_));
 sky130_fd_sc_hd__o21ba_1 _2939_ (.A1(_0276_),
    .A2(_0339_),
    .B1_N(\disp_song.note2[26] ),
    .X(_0340_));
 sky130_fd_sc_hd__o21ai_1 _2940_ (.A1(_0276_),
    .A2(_0336_),
    .B1(\disp_song.note2[26] ),
    .Y(_0341_));
 sky130_fd_sc_hd__o21ai_2 _2941_ (.A1(_2655_),
    .A2(_0340_),
    .B1(_0341_),
    .Y(\disp_song.um.drum.next_note2[26] ));
 sky130_fd_sc_hd__o21ai_1 _2942_ (.A1(_0279_),
    .A2(_0337_),
    .B1(\disp_song.note2[27] ),
    .Y(_0342_));
 sky130_fd_sc_hd__o31a_1 _2943_ (.A1(_2655_),
    .A2(_0279_),
    .A3(_0339_),
    .B1(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__inv_2 _2944_ (.A(_0343_),
    .Y(\disp_song.um.drum.next_note2[27] ));
 sky130_fd_sc_hd__o21a_1 _2945_ (.A1(_0163_),
    .A2(_0337_),
    .B1(\disp_song.note2[28] ),
    .X(_0344_));
 sky130_fd_sc_hd__a31o_1 _2946_ (.A1(_0269_),
    .A2(_0164_),
    .A3(_0334_),
    .B1(_0344_),
    .X(\disp_song.um.drum.next_note2[28] ));
 sky130_fd_sc_hd__nor2_1 _2947_ (.A(_2655_),
    .B(_0339_),
    .Y(_0345_));
 sky130_fd_sc_hd__or2_1 _2948_ (.A(_0307_),
    .B(_0337_),
    .X(_0346_));
 sky130_fd_sc_hd__a22o_1 _2949_ (.A1(_0285_),
    .A2(_0345_),
    .B1(_0346_),
    .B2(net244),
    .X(\disp_song.um.drum.next_note2[29] ));
 sky130_fd_sc_hd__or2_1 _2950_ (.A(_0310_),
    .B(_0337_),
    .X(_0347_));
 sky130_fd_sc_hd__a22o_1 _2951_ (.A1(_0288_),
    .A2(_0345_),
    .B1(_0347_),
    .B2(net200),
    .X(\disp_song.um.drum.next_note2[30] ));
 sky130_fd_sc_hd__or2_1 _2952_ (.A(_0313_),
    .B(_0337_),
    .X(_0348_));
 sky130_fd_sc_hd__a22o_1 _2953_ (.A1(_0291_),
    .A2(_0345_),
    .B1(_0348_),
    .B2(net255),
    .X(\disp_song.um.drum.next_note2[31] ));
 sky130_fd_sc_hd__or3_1 _2954_ (.A(_2661_),
    .B(_0183_),
    .C(_0265_),
    .X(_0349_));
 sky130_fd_sc_hd__or3b_1 _2955_ (.A(_2661_),
    .B(_0183_),
    .C_N(_0264_),
    .X(_0350_));
 sky130_fd_sc_hd__a21bo_1 _2956_ (.A1(\disp_song.note1[0] ),
    .A2(_0349_),
    .B1_N(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_2 _2957_ (.A(_0351_),
    .X(\disp_song.um.drum.next_note1[0] ));
 sky130_fd_sc_hd__clkinv_4 _2958_ (.A(\modetrans.mode[2] ),
    .Y(_0352_));
 sky130_fd_sc_hd__or3b_2 _2959_ (.A(\disp_song.um.idx_note1[2] ),
    .B(_0179_),
    .C_N(\disp_song.um.idx_note1[0] ),
    .X(_0353_));
 sky130_fd_sc_hd__or2_1 _2960_ (.A(_0352_),
    .B(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__or3b_1 _2961_ (.A(_0354_),
    .B(_2661_),
    .C_N(_0194_),
    .X(_0355_));
 sky130_fd_sc_hd__nand2_1 _2962_ (.A(\disp_song.um.idx_note1[4] ),
    .B(_0182_),
    .Y(_0356_));
 sky130_fd_sc_hd__and2_2 _2963_ (.A(_0183_),
    .B(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__nand2_1 _2964_ (.A(_2657_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__nand2_2 _2965_ (.A(_2660_),
    .B(_0357_),
    .Y(_0359_));
 sky130_fd_sc_hd__or2_1 _2966_ (.A(_0359_),
    .B(_0355_),
    .X(_0360_));
 sky130_fd_sc_hd__a2bb2o_1 _2967_ (.A1_N(_0355_),
    .A2_N(_0358_),
    .B1(_0360_),
    .B2(\disp_song.note1[1] ),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_2 _2968_ (.A(_0361_),
    .X(\disp_song.um.drum.next_note1[1] ));
 sky130_fd_sc_hd__or3b_2 _2969_ (.A(\disp_song.um.idx_note1[0] ),
    .B(\disp_song.um.idx_note1[2] ),
    .C_N(_0179_),
    .X(_0362_));
 sky130_fd_sc_hd__inv_2 _2970_ (.A(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__nand2_2 _2971_ (.A(_0194_),
    .B(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__or2_1 _2972_ (.A(_2661_),
    .B(_0352_),
    .X(_0365_));
 sky130_fd_sc_hd__clkbuf_4 _2973_ (.A(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__or2_2 _2974_ (.A(_0358_),
    .B(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__or2_2 _2975_ (.A(_0359_),
    .B(_0366_),
    .X(_0368_));
 sky130_fd_sc_hd__o21ai_1 _2976_ (.A1(_0368_),
    .A2(_0364_),
    .B1(\disp_song.note1[2] ),
    .Y(_0369_));
 sky130_fd_sc_hd__o21ai_2 _2977_ (.A1(_0364_),
    .A2(_0367_),
    .B1(_0369_),
    .Y(\disp_song.um.drum.next_note1[2] ));
 sky130_fd_sc_hd__nand3_2 _2978_ (.A(\disp_song.um.idx_note1[0] ),
    .B(_0178_),
    .C(_0179_),
    .Y(_0370_));
 sky130_fd_sc_hd__or2_1 _2979_ (.A(\disp_song.um.idx_note1[3] ),
    .B(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__o21ai_1 _2980_ (.A1(_0368_),
    .A2(_0371_),
    .B1(\disp_song.note1[3] ),
    .Y(_0372_));
 sky130_fd_sc_hd__o21a_1 _2981_ (.A1(_0367_),
    .A2(_0371_),
    .B1(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__inv_2 _2982_ (.A(_0373_),
    .Y(\disp_song.um.drum.next_note1[3] ));
 sky130_fd_sc_hd__nand2_2 _2983_ (.A(\disp_song.um.idx_note1[2] ),
    .B(_0180_),
    .Y(_0374_));
 sky130_fd_sc_hd__or2_2 _2984_ (.A(\disp_song.um.idx_note1[3] ),
    .B(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__o21ai_1 _2985_ (.A1(_0368_),
    .A2(_0375_),
    .B1(\disp_song.note1[4] ),
    .Y(_0376_));
 sky130_fd_sc_hd__o21ai_2 _2986_ (.A1(_0367_),
    .A2(_0375_),
    .B1(_0376_),
    .Y(\disp_song.um.drum.next_note1[4] ));
 sky130_fd_sc_hd__or4bb_2 _2987_ (.A(\disp_song.um.idx_note1[3] ),
    .B(_0179_),
    .C_N(\disp_song.um.idx_note1[0] ),
    .D_N(\disp_song.um.idx_note1[2] ),
    .X(_0377_));
 sky130_fd_sc_hd__or2_1 _2988_ (.A(_0368_),
    .B(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__a2bb2o_1 _2989_ (.A1_N(_0367_),
    .A2_N(_0377_),
    .B1(_0378_),
    .B2(\disp_song.note1[5] ),
    .X(_0379_));
 sky130_fd_sc_hd__clkbuf_2 _2990_ (.A(_0379_),
    .X(\disp_song.um.drum.next_note1[5] ));
 sky130_fd_sc_hd__nor2_2 _2991_ (.A(_0358_),
    .B(_0366_),
    .Y(_0380_));
 sky130_fd_sc_hd__and4b_1 _2992_ (.A_N(\disp_song.um.idx_note1[0] ),
    .B(\disp_song.um.idx_note1[2] ),
    .C(_0177_),
    .D(_0179_),
    .X(_0381_));
 sky130_fd_sc_hd__nor2_2 _2993_ (.A(_0359_),
    .B(_0366_),
    .Y(_0382_));
 sky130_fd_sc_hd__nand2_1 _2994_ (.A(_0382_),
    .B(_0381_),
    .Y(_0383_));
 sky130_fd_sc_hd__a22o_1 _2995_ (.A1(_0380_),
    .A2(_0381_),
    .B1(_0383_),
    .B2(net262),
    .X(\disp_song.um.drum.next_note1[6] ));
 sky130_fd_sc_hd__and4_1 _2996_ (.A(\disp_song.um.idx_note1[0] ),
    .B(\disp_song.um.idx_note1[2] ),
    .C(_0177_),
    .D(_0179_),
    .X(_0384_));
 sky130_fd_sc_hd__nand2_1 _2997_ (.A(_0382_),
    .B(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__a22o_1 _2998_ (.A1(_0380_),
    .A2(_0384_),
    .B1(_0385_),
    .B2(net268),
    .X(\disp_song.um.drum.next_note1[7] ));
 sky130_fd_sc_hd__nand2_1 _2999_ (.A(\disp_song.um.idx_note1[3] ),
    .B(_0181_),
    .Y(_0386_));
 sky130_fd_sc_hd__o21ai_1 _3000_ (.A1(_0368_),
    .A2(_0386_),
    .B1(net247),
    .Y(_0387_));
 sky130_fd_sc_hd__o21ai_1 _3001_ (.A1(_0367_),
    .A2(_0386_),
    .B1(_0387_),
    .Y(\disp_song.um.drum.next_note1[8] ));
 sky130_fd_sc_hd__and3b_1 _3002_ (.A_N(_0179_),
    .B(\disp_song.um.idx_note1[0] ),
    .C(_0178_),
    .X(_0388_));
 sky130_fd_sc_hd__nor3_1 _3003_ (.A(_2661_),
    .B(_0194_),
    .C(_0358_),
    .Y(_0389_));
 sky130_fd_sc_hd__or4_1 _3004_ (.A(_2661_),
    .B(_0194_),
    .C(_0359_),
    .D(_0354_),
    .X(_0390_));
 sky130_fd_sc_hd__a32o_1 _3005_ (.A1(_2654_),
    .A2(_0388_),
    .A3(_0389_),
    .B1(_0390_),
    .B2(\disp_song.note1[9] ),
    .X(_0391_));
 sky130_fd_sc_hd__clkbuf_2 _3006_ (.A(_0391_),
    .X(\disp_song.um.drum.next_note1[9] ));
 sky130_fd_sc_hd__nor4_1 _3007_ (.A(_2661_),
    .B(_0352_),
    .C(_0194_),
    .D(_0359_),
    .Y(_0392_));
 sky130_fd_sc_hd__nand2_1 _3008_ (.A(_0363_),
    .B(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__and2_1 _3009_ (.A(_2654_),
    .B(_0389_),
    .X(_0394_));
 sky130_fd_sc_hd__a22o_1 _3010_ (.A1(\disp_song.note1[10] ),
    .A2(_0393_),
    .B1(_0394_),
    .B2(_0363_),
    .X(\disp_song.um.drum.next_note1[10] ));
 sky130_fd_sc_hd__o41a_1 _3011_ (.A1(_0194_),
    .A2(_0359_),
    .A3(_0366_),
    .A4(_0370_),
    .B1(\disp_song.note1[11] ),
    .X(_0395_));
 sky130_fd_sc_hd__a41o_1 _3012_ (.A1(\disp_song.um.idx_note1[0] ),
    .A2(_0178_),
    .A3(_0179_),
    .A4(_0394_),
    .B1(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_2 _3013_ (.A(_0396_),
    .X(\disp_song.um.drum.next_note1[11] ));
 sky130_fd_sc_hd__or2b_1 _3014_ (.A(_0374_),
    .B_N(_0392_),
    .X(_0397_));
 sky130_fd_sc_hd__a32o_1 _3015_ (.A1(\disp_song.um.idx_note1[2] ),
    .A2(_0180_),
    .A3(_0394_),
    .B1(_0397_),
    .B2(net183),
    .X(\disp_song.um.drum.next_note1[12] ));
 sky130_fd_sc_hd__and4b_1 _3016_ (.A_N(_0179_),
    .B(\disp_song.um.idx_note1[3] ),
    .C(\disp_song.um.idx_note1[2] ),
    .D(\disp_song.um.idx_note1[0] ),
    .X(_0398_));
 sky130_fd_sc_hd__nand2_1 _3017_ (.A(_0382_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__a22o_1 _3018_ (.A1(_0380_),
    .A2(_0398_),
    .B1(_0399_),
    .B2(net246),
    .X(\disp_song.um.drum.next_note1[13] ));
 sky130_fd_sc_hd__and4b_2 _3019_ (.A_N(\disp_song.um.idx_note1[0] ),
    .B(\disp_song.um.idx_note1[2] ),
    .C(\disp_song.um.idx_note1[3] ),
    .D(_0179_),
    .X(_0400_));
 sky130_fd_sc_hd__nand2_1 _3020_ (.A(_0382_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__a22o_1 _3021_ (.A1(_0380_),
    .A2(_0400_),
    .B1(_0401_),
    .B2(net250),
    .X(\disp_song.um.drum.next_note1[14] ));
 sky130_fd_sc_hd__and4_1 _3022_ (.A(\disp_song.um.idx_note1[0] ),
    .B(\disp_song.um.idx_note1[2] ),
    .C(\disp_song.um.idx_note1[3] ),
    .D(_0179_),
    .X(_0402_));
 sky130_fd_sc_hd__nand2_1 _3023_ (.A(_0382_),
    .B(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__a22o_1 _3024_ (.A1(_0380_),
    .A2(_0402_),
    .B1(_0403_),
    .B2(net237),
    .X(\disp_song.um.drum.next_note1[15] ));
 sky130_fd_sc_hd__inv_2 _3025_ (.A(\disp_song.um.idx_note1[4] ),
    .Y(_0404_));
 sky130_fd_sc_hd__nor2_1 _3026_ (.A(_2661_),
    .B(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__o41a_1 _3027_ (.A1(_2661_),
    .A2(_0404_),
    .A3(_0182_),
    .A4(_0265_),
    .B1(\disp_song.note1[16] ),
    .X(_0406_));
 sky130_fd_sc_hd__a41o_1 _3028_ (.A1(_0177_),
    .A2(_0181_),
    .A3(_0264_),
    .A4(_0405_),
    .B1(_0406_),
    .X(\disp_song.um.drum.next_note1[16] ));
 sky130_fd_sc_hd__nor2_1 _3029_ (.A(_0357_),
    .B(_0355_),
    .Y(_0407_));
 sky130_fd_sc_hd__nand2_1 _3030_ (.A(_2660_),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__a22o_1 _3031_ (.A1(_0269_),
    .A2(_0407_),
    .B1(_0408_),
    .B2(\disp_song.note1[17] ),
    .X(\disp_song.um.drum.next_note1[17] ));
 sky130_fd_sc_hd__nor2_1 _3032_ (.A(_2661_),
    .B(_0357_),
    .Y(_0409_));
 sky130_fd_sc_hd__nand2_2 _3033_ (.A(_0264_),
    .B(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__or3_1 _3034_ (.A(_2661_),
    .B(_0265_),
    .C(_0357_),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_2 _3035_ (.A(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__o21ai_1 _3036_ (.A1(_0364_),
    .A2(_0412_),
    .B1(net240),
    .Y(_0413_));
 sky130_fd_sc_hd__o21ai_1 _3037_ (.A1(_0364_),
    .A2(_0410_),
    .B1(_0413_),
    .Y(\disp_song.um.drum.next_note1[18] ));
 sky130_fd_sc_hd__or2_1 _3038_ (.A(_0371_),
    .B(_0412_),
    .X(_0414_));
 sky130_fd_sc_hd__o2bb2a_1 _3039_ (.A1_N(\disp_song.note1[19] ),
    .A2_N(_0414_),
    .B1(_0410_),
    .B2(_0371_),
    .X(_0415_));
 sky130_fd_sc_hd__inv_2 _3040_ (.A(_0415_),
    .Y(\disp_song.um.drum.next_note1[19] ));
 sky130_fd_sc_hd__o21ai_1 _3041_ (.A1(_0375_),
    .A2(_0412_),
    .B1(net163),
    .Y(_0416_));
 sky130_fd_sc_hd__o21ai_1 _3042_ (.A1(_0375_),
    .A2(_0410_),
    .B1(_0416_),
    .Y(\disp_song.um.drum.next_note1[20] ));
 sky130_fd_sc_hd__o21ai_1 _3043_ (.A1(_0377_),
    .A2(_0412_),
    .B1(net245),
    .Y(_0417_));
 sky130_fd_sc_hd__o21ai_2 _3044_ (.A1(_0377_),
    .A2(_0410_),
    .B1(_0417_),
    .Y(\disp_song.um.drum.next_note1[21] ));
 sky130_fd_sc_hd__and2_1 _3045_ (.A(_0264_),
    .B(_0409_),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_2 _3046_ (.A(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__and3_1 _3047_ (.A(_2654_),
    .B(_2660_),
    .C(_0409_),
    .X(_0420_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3048_ (.A(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__nand2_1 _3049_ (.A(_0381_),
    .B(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__a22o_1 _3050_ (.A1(_0381_),
    .A2(_0419_),
    .B1(_0422_),
    .B2(net205),
    .X(\disp_song.um.drum.next_note1[22] ));
 sky130_fd_sc_hd__nand2_1 _3051_ (.A(_0384_),
    .B(_0421_),
    .Y(_0423_));
 sky130_fd_sc_hd__a22o_1 _3052_ (.A1(_0384_),
    .A2(_0419_),
    .B1(_0423_),
    .B2(net204),
    .X(\disp_song.um.drum.next_note1[23] ));
 sky130_fd_sc_hd__o21ai_1 _3053_ (.A1(_0386_),
    .A2(_0412_),
    .B1(net259),
    .Y(_0424_));
 sky130_fd_sc_hd__o21ai_1 _3054_ (.A1(_0386_),
    .A2(_0410_),
    .B1(_0424_),
    .Y(\disp_song.um.drum.next_note1[24] ));
 sky130_fd_sc_hd__or2_2 _3055_ (.A(_0194_),
    .B(_0410_),
    .X(_0425_));
 sky130_fd_sc_hd__or2_2 _3056_ (.A(_0194_),
    .B(_0412_),
    .X(_0426_));
 sky130_fd_sc_hd__o21ai_1 _3057_ (.A1(_0353_),
    .A2(_0426_),
    .B1(net150),
    .Y(_0427_));
 sky130_fd_sc_hd__o21ai_2 _3058_ (.A1(_0353_),
    .A2(_0425_),
    .B1(_0427_),
    .Y(\disp_song.um.drum.next_note1[25] ));
 sky130_fd_sc_hd__o21ai_1 _3059_ (.A1(_0362_),
    .A2(_0426_),
    .B1(net154),
    .Y(_0428_));
 sky130_fd_sc_hd__o21ai_1 _3060_ (.A1(_0362_),
    .A2(_0425_),
    .B1(_0428_),
    .Y(\disp_song.um.drum.next_note1[26] ));
 sky130_fd_sc_hd__o21ai_1 _3061_ (.A1(_0370_),
    .A2(_0426_),
    .B1(\disp_song.note1[27] ),
    .Y(_0429_));
 sky130_fd_sc_hd__o21a_1 _3062_ (.A1(_0370_),
    .A2(_0425_),
    .B1(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__inv_2 _3063_ (.A(_0430_),
    .Y(\disp_song.um.drum.next_note1[27] ));
 sky130_fd_sc_hd__o21ai_1 _3064_ (.A1(_0374_),
    .A2(_0426_),
    .B1(net122),
    .Y(_0431_));
 sky130_fd_sc_hd__o21ai_2 _3065_ (.A1(_0374_),
    .A2(_0425_),
    .B1(_0431_),
    .Y(\disp_song.um.drum.next_note1[28] ));
 sky130_fd_sc_hd__nand2_1 _3066_ (.A(_0398_),
    .B(_0421_),
    .Y(_0432_));
 sky130_fd_sc_hd__a22o_1 _3067_ (.A1(_0398_),
    .A2(_0419_),
    .B1(_0432_),
    .B2(net165),
    .X(\disp_song.um.drum.next_note1[29] ));
 sky130_fd_sc_hd__nand2_1 _3068_ (.A(_0400_),
    .B(_0421_),
    .Y(_0433_));
 sky130_fd_sc_hd__a22o_1 _3069_ (.A1(_0400_),
    .A2(_0419_),
    .B1(_0433_),
    .B2(net197),
    .X(\disp_song.um.drum.next_note1[30] ));
 sky130_fd_sc_hd__nand2_1 _3070_ (.A(_0402_),
    .B(_0421_),
    .Y(_0434_));
 sky130_fd_sc_hd__a22o_1 _3071_ (.A1(_0402_),
    .A2(_0419_),
    .B1(_0434_),
    .B2(net160),
    .X(\disp_song.um.drum.next_note1[31] ));
 sky130_fd_sc_hd__and2_1 _3072_ (.A(\game.addmisses.a[12] ),
    .B(\game.addmisses.add4.b[0] ),
    .X(_0435_));
 sky130_fd_sc_hd__nor2_1 _3073_ (.A(\game.addmisses.a[12] ),
    .B(\game.addmisses.add4.b[0] ),
    .Y(_0436_));
 sky130_fd_sc_hd__nor2_1 _3074_ (.A(_0435_),
    .B(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__nand2_1 _3075_ (.A(\game.addmisses.a[9] ),
    .B(\game.addmisses.add3.b[1] ),
    .Y(_0438_));
 sky130_fd_sc_hd__or2_1 _3076_ (.A(\game.addmisses.a[9] ),
    .B(\game.addmisses.add3.b[1] ),
    .X(_0439_));
 sky130_fd_sc_hd__nand2_1 _3077_ (.A(_0438_),
    .B(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__nand2_1 _3078_ (.A(\game.addmisses.a[8] ),
    .B(\game.addmisses.add3.b[0] ),
    .Y(_0441_));
 sky130_fd_sc_hd__or2_1 _3079_ (.A(\game.addmisses.a[8] ),
    .B(\game.addmisses.add3.b[0] ),
    .X(_0442_));
 sky130_fd_sc_hd__nand2_2 _3080_ (.A(_0441_),
    .B(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__nand2_1 _3081_ (.A(\game.addmisses.a[5] ),
    .B(\game.addmisses.add2.b[1] ),
    .Y(_0444_));
 sky130_fd_sc_hd__or2_1 _3082_ (.A(\game.addmisses.a[5] ),
    .B(\game.addmisses.add2.b[1] ),
    .X(_0445_));
 sky130_fd_sc_hd__nand2_2 _3083_ (.A(_0444_),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__nand2_1 _3084_ (.A(\game.addmisses.a[4] ),
    .B(\game.addmisses.add2.b[0] ),
    .Y(_0447_));
 sky130_fd_sc_hd__or2_1 _3085_ (.A(\game.addmisses.a[4] ),
    .B(\game.addmisses.add2.b[0] ),
    .X(_0448_));
 sky130_fd_sc_hd__nand2_2 _3086_ (.A(_0447_),
    .B(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__nand2_2 _3087_ (.A(\game.addmisses.add1.b[0] ),
    .B(\game.addmisses.a[0] ),
    .Y(_0450_));
 sky130_fd_sc_hd__nand2_1 _3088_ (.A(\game.addmisses.a[1] ),
    .B(\game.addmisses.add1.b[1] ),
    .Y(_0451_));
 sky130_fd_sc_hd__or2_1 _3089_ (.A(\game.addmisses.a[1] ),
    .B(\game.addmisses.add1.b[1] ),
    .X(_0452_));
 sky130_fd_sc_hd__nand2_2 _3090_ (.A(_0451_),
    .B(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__xor2_4 _3091_ (.A(_0450_),
    .B(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__nor2_1 _3092_ (.A(\game.addmisses.a[1] ),
    .B(\game.addmisses.add1.b[1] ),
    .Y(_0455_));
 sky130_fd_sc_hd__o21a_2 _3093_ (.A1(_0450_),
    .A2(_0455_),
    .B1(_0451_),
    .X(_0456_));
 sky130_fd_sc_hd__nor2_1 _3094_ (.A(\game.addmisses.a[2] ),
    .B(\game.addmisses.add1.b[2] ),
    .Y(_0457_));
 sky130_fd_sc_hd__nand2_1 _3095_ (.A(\game.addmisses.a[2] ),
    .B(\game.addmisses.add1.b[2] ),
    .Y(_0458_));
 sky130_fd_sc_hd__and2b_1 _3096_ (.A_N(_0457_),
    .B(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__xnor2_4 _3097_ (.A(_0456_),
    .B(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__nor2_1 _3098_ (.A(_0454_),
    .B(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__nor2_1 _3099_ (.A(\game.addmisses.a[3] ),
    .B(\game.addmisses.add1.b[3] ),
    .Y(_0462_));
 sky130_fd_sc_hd__nand2_1 _3100_ (.A(\game.addmisses.a[3] ),
    .B(\game.addmisses.add1.b[3] ),
    .Y(_0463_));
 sky130_fd_sc_hd__or2b_2 _3101_ (.A(_0462_),
    .B_N(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__o21a_2 _3102_ (.A1(_0456_),
    .A2(_0457_),
    .B1(_0458_),
    .X(_0465_));
 sky130_fd_sc_hd__xnor2_4 _3103_ (.A(_0464_),
    .B(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__o21a_1 _3104_ (.A1(_0462_),
    .A2(_0465_),
    .B1(_0463_),
    .X(_0467_));
 sky130_fd_sc_hd__o21a_4 _3105_ (.A1(_0461_),
    .A2(_0466_),
    .B1(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__nor3_1 _3106_ (.A(_0461_),
    .B(_0463_),
    .C(_0465_),
    .Y(_0469_));
 sky130_fd_sc_hd__o31a_2 _3107_ (.A1(_0449_),
    .A2(_0468_),
    .A3(_0469_),
    .B1(_0447_),
    .X(_0470_));
 sky130_fd_sc_hd__xnor2_4 _3108_ (.A(_0446_),
    .B(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__o21a_1 _3109_ (.A1(_0446_),
    .A2(_0470_),
    .B1(_0444_),
    .X(_0472_));
 sky130_fd_sc_hd__nor2_1 _3110_ (.A(\game.addmisses.a[6] ),
    .B(\game.addmisses.add2.b[2] ),
    .Y(_0473_));
 sky130_fd_sc_hd__nand2_1 _3111_ (.A(\game.addmisses.a[6] ),
    .B(\game.addmisses.add2.b[2] ),
    .Y(_0474_));
 sky130_fd_sc_hd__or2b_1 _3112_ (.A(_0473_),
    .B_N(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__xnor2_2 _3113_ (.A(_0472_),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__and2_1 _3114_ (.A(_0471_),
    .B(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__nor2_1 _3115_ (.A(\game.addmisses.a[7] ),
    .B(\game.addmisses.add2.b[3] ),
    .Y(_0478_));
 sky130_fd_sc_hd__nand2_1 _3116_ (.A(\game.addmisses.a[7] ),
    .B(\game.addmisses.add2.b[3] ),
    .Y(_0479_));
 sky130_fd_sc_hd__or2b_1 _3117_ (.A(_0478_),
    .B_N(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__o21a_1 _3118_ (.A1(_0472_),
    .A2(_0473_),
    .B1(_0474_),
    .X(_0481_));
 sky130_fd_sc_hd__xnor2_1 _3119_ (.A(_0480_),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__o21ai_2 _3120_ (.A1(_0478_),
    .A2(_0481_),
    .B1(_0479_),
    .Y(_0483_));
 sky130_fd_sc_hd__o21ba_2 _3121_ (.A1(_0477_),
    .A2(_0482_),
    .B1_N(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__nor3_2 _3122_ (.A(_0477_),
    .B(_0479_),
    .C(_0481_),
    .Y(_0485_));
 sky130_fd_sc_hd__o31ai_4 _3123_ (.A1(_0443_),
    .A2(_0484_),
    .A3(_0485_),
    .B1(_0441_),
    .Y(_0486_));
 sky130_fd_sc_hd__xor2_2 _3124_ (.A(_0440_),
    .B(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__a21boi_2 _3125_ (.A1(_0439_),
    .A2(_0486_),
    .B1_N(_0438_),
    .Y(_0488_));
 sky130_fd_sc_hd__nor2_1 _3126_ (.A(\game.addmisses.a[10] ),
    .B(\game.addmisses.add3.b[2] ),
    .Y(_0489_));
 sky130_fd_sc_hd__nand2_1 _3127_ (.A(\game.addmisses.a[10] ),
    .B(\game.addmisses.add3.b[2] ),
    .Y(_0490_));
 sky130_fd_sc_hd__or2b_1 _3128_ (.A(_0489_),
    .B_N(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__xnor2_2 _3129_ (.A(_0488_),
    .B(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__nand2_1 _3130_ (.A(_0487_),
    .B(_0492_),
    .Y(_0493_));
 sky130_fd_sc_hd__nor2_1 _3131_ (.A(\game.addmisses.a[11] ),
    .B(\game.addmisses.add3.b[3] ),
    .Y(_0494_));
 sky130_fd_sc_hd__nand2_1 _3132_ (.A(\game.addmisses.a[11] ),
    .B(\game.addmisses.add3.b[3] ),
    .Y(_0495_));
 sky130_fd_sc_hd__or2b_1 _3133_ (.A(_0494_),
    .B_N(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__o21a_1 _3134_ (.A1(_0488_),
    .A2(_0489_),
    .B1(_0490_),
    .X(_0497_));
 sky130_fd_sc_hd__xor2_2 _3135_ (.A(_0496_),
    .B(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__o21ai_1 _3136_ (.A1(_0494_),
    .A2(_0497_),
    .B1(_0495_),
    .Y(_0499_));
 sky130_fd_sc_hd__a21o_1 _3137_ (.A1(_0493_),
    .A2(_0498_),
    .B1(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__or3b_1 _3138_ (.A(_0495_),
    .B(_0497_),
    .C_N(_0493_),
    .X(_0501_));
 sky130_fd_sc_hd__and3_1 _3139_ (.A(_0437_),
    .B(_0500_),
    .C(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__a21oi_1 _3140_ (.A1(_0500_),
    .A2(_0501_),
    .B1(_0437_),
    .Y(_0503_));
 sky130_fd_sc_hd__or2_1 _3141_ (.A(_0502_),
    .B(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__a31o_1 _3142_ (.A1(_0437_),
    .A2(_0500_),
    .A3(_0501_),
    .B1(_0435_),
    .X(_0505_));
 sky130_fd_sc_hd__or2_1 _3143_ (.A(\game.addmisses.a[13] ),
    .B(\game.addmisses.add4.b[1] ),
    .X(_0506_));
 sky130_fd_sc_hd__and2_1 _3144_ (.A(\game.addmisses.a[13] ),
    .B(\game.addmisses.add4.b[1] ),
    .X(_0507_));
 sky130_fd_sc_hd__a21oi_2 _3145_ (.A1(_0505_),
    .A2(_0506_),
    .B1(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__and2_1 _3146_ (.A(\game.addmisses.a[14] ),
    .B(\game.addmisses.add4.b[2] ),
    .X(_0509_));
 sky130_fd_sc_hd__nor2_1 _3147_ (.A(\game.addmisses.a[14] ),
    .B(\game.addmisses.add4.b[2] ),
    .Y(_0510_));
 sky130_fd_sc_hd__nor2_1 _3148_ (.A(_0509_),
    .B(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__xnor2_2 _3149_ (.A(_0508_),
    .B(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__or2b_1 _3150_ (.A(_0507_),
    .B_N(_0506_),
    .X(_0513_));
 sky130_fd_sc_hd__xnor2_2 _3151_ (.A(_0505_),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__nor2_1 _3152_ (.A(_0514_),
    .B(_0512_),
    .Y(_0515_));
 sky130_fd_sc_hd__o21ba_1 _3153_ (.A1(_0508_),
    .A2(_0510_),
    .B1_N(_0509_),
    .X(_0516_));
 sky130_fd_sc_hd__nand2_1 _3154_ (.A(\game.addmisses.a[15] ),
    .B(\game.addmisses.add4.b[3] ),
    .Y(_0517_));
 sky130_fd_sc_hd__or2_1 _3155_ (.A(\game.addmisses.a[15] ),
    .B(\game.addmisses.add4.b[3] ),
    .X(_0518_));
 sky130_fd_sc_hd__nand2_1 _3156_ (.A(_0517_),
    .B(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__xnor2_1 _3157_ (.A(_0516_),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__nor2_1 _3158_ (.A(\game.addmisses.a[15] ),
    .B(\game.addmisses.add4.b[3] ),
    .Y(_0521_));
 sky130_fd_sc_hd__o21ai_1 _3159_ (.A1(_0521_),
    .A2(_0516_),
    .B1(_0517_),
    .Y(_0522_));
 sky130_fd_sc_hd__o21ba_1 _3160_ (.A1(_0515_),
    .A2(_0520_),
    .B1_N(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__xnor2_2 _3161_ (.A(_0514_),
    .B(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__or2_1 _3162_ (.A(_0514_),
    .B(_0512_),
    .X(_0525_));
 sky130_fd_sc_hd__nand2_1 _3163_ (.A(_0525_),
    .B(_0522_),
    .Y(_0526_));
 sky130_fd_sc_hd__mux2_2 _3164_ (.A0(_0525_),
    .A1(_0526_),
    .S(_0520_),
    .X(_0527_));
 sky130_fd_sc_hd__o21bai_1 _3165_ (.A1(_0512_),
    .A2(_0524_),
    .B1_N(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__and2_1 _3166_ (.A(\game.addhits.a[12] ),
    .B(\game.addhits.add4.b[0] ),
    .X(_0529_));
 sky130_fd_sc_hd__nor2_1 _3167_ (.A(\game.addhits.a[12] ),
    .B(\game.addhits.add4.b[0] ),
    .Y(_0530_));
 sky130_fd_sc_hd__nor2_1 _3168_ (.A(_0529_),
    .B(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__nand2_1 _3169_ (.A(\game.addhits.a[9] ),
    .B(\game.addhits.add3.b[1] ),
    .Y(_0532_));
 sky130_fd_sc_hd__or2_1 _3170_ (.A(\game.addhits.a[9] ),
    .B(\game.addhits.add3.b[1] ),
    .X(_0533_));
 sky130_fd_sc_hd__nand2_1 _3171_ (.A(_0532_),
    .B(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__and2_1 _3172_ (.A(\game.addhits.a[8] ),
    .B(\game.addhits.add3.b[0] ),
    .X(_0535_));
 sky130_fd_sc_hd__nor2_1 _3173_ (.A(\game.addhits.a[8] ),
    .B(\game.addhits.add3.b[0] ),
    .Y(_0536_));
 sky130_fd_sc_hd__nor2_1 _3174_ (.A(_0535_),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__nand2_1 _3175_ (.A(\game.addhits.a[5] ),
    .B(\game.addhits.add2.b[1] ),
    .Y(_0538_));
 sky130_fd_sc_hd__or2_1 _3176_ (.A(\game.addhits.a[5] ),
    .B(\game.addhits.add2.b[1] ),
    .X(_0539_));
 sky130_fd_sc_hd__nand2_2 _3177_ (.A(_0538_),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__and2_1 _3178_ (.A(\game.addhits.a[4] ),
    .B(\game.addhits.add2.b[0] ),
    .X(_0541_));
 sky130_fd_sc_hd__nor2_1 _3179_ (.A(\game.addhits.a[4] ),
    .B(\game.addhits.add2.b[0] ),
    .Y(_0542_));
 sky130_fd_sc_hd__nor2_1 _3180_ (.A(_0541_),
    .B(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__nand2_2 _3181_ (.A(\game.addhits.add1.b[0] ),
    .B(\game.addhits.a[0] ),
    .Y(_0544_));
 sky130_fd_sc_hd__xor2_4 _3182_ (.A(\game.addhits.a[1] ),
    .B(\game.addhits.add1.b[1] ),
    .X(_0545_));
 sky130_fd_sc_hd__xnor2_4 _3183_ (.A(_0544_),
    .B(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__and2_1 _3184_ (.A(\game.addhits.a[1] ),
    .B(\game.addhits.add1.b[1] ),
    .X(_0547_));
 sky130_fd_sc_hd__a31oi_4 _3185_ (.A1(\game.addhits.add1.b[0] ),
    .A2(\game.addhits.a[0] ),
    .A3(_0545_),
    .B1(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__nor2_1 _3186_ (.A(\game.addhits.a[2] ),
    .B(\game.addhits.add1.b[2] ),
    .Y(_0549_));
 sky130_fd_sc_hd__nand2_1 _3187_ (.A(\game.addhits.a[2] ),
    .B(\game.addhits.add1.b[2] ),
    .Y(_0550_));
 sky130_fd_sc_hd__and2b_1 _3188_ (.A_N(_0549_),
    .B(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__xnor2_2 _3189_ (.A(_0548_),
    .B(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__nor2_2 _3190_ (.A(_0546_),
    .B(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__nor2_1 _3191_ (.A(\game.addhits.a[3] ),
    .B(\game.addhits.add1.b[3] ),
    .Y(_0554_));
 sky130_fd_sc_hd__nand2_1 _3192_ (.A(\game.addhits.a[3] ),
    .B(\game.addhits.add1.b[3] ),
    .Y(_0555_));
 sky130_fd_sc_hd__or2b_1 _3193_ (.A(_0554_),
    .B_N(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__o21a_1 _3194_ (.A1(_0548_),
    .A2(_0549_),
    .B1(_0550_),
    .X(_0557_));
 sky130_fd_sc_hd__xnor2_2 _3195_ (.A(_0556_),
    .B(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__o21a_1 _3196_ (.A1(_0554_),
    .A2(_0557_),
    .B1(_0555_),
    .X(_0559_));
 sky130_fd_sc_hd__o21ai_4 _3197_ (.A1(_0553_),
    .A2(_0558_),
    .B1(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__or3_2 _3198_ (.A(_0553_),
    .B(_0555_),
    .C(_0557_),
    .X(_0561_));
 sky130_fd_sc_hd__a31oi_4 _3199_ (.A1(_0543_),
    .A2(_0560_),
    .A3(_0561_),
    .B1(_0541_),
    .Y(_0562_));
 sky130_fd_sc_hd__xor2_4 _3200_ (.A(_0540_),
    .B(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__nor2_1 _3201_ (.A(\game.addhits.a[6] ),
    .B(\game.addhits.add2.b[2] ),
    .Y(_0564_));
 sky130_fd_sc_hd__nand2_1 _3202_ (.A(\game.addhits.a[6] ),
    .B(\game.addhits.add2.b[2] ),
    .Y(_0565_));
 sky130_fd_sc_hd__or2b_1 _3203_ (.A(_0564_),
    .B_N(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__o21a_1 _3204_ (.A1(_0540_),
    .A2(_0562_),
    .B1(_0538_),
    .X(_0567_));
 sky130_fd_sc_hd__xor2_1 _3205_ (.A(_0566_),
    .B(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__nor2_2 _3206_ (.A(_0563_),
    .B(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__nor2_1 _3207_ (.A(\game.addhits.a[7] ),
    .B(\game.addhits.add2.b[3] ),
    .Y(_0570_));
 sky130_fd_sc_hd__nand2_1 _3208_ (.A(\game.addhits.a[7] ),
    .B(\game.addhits.add2.b[3] ),
    .Y(_0571_));
 sky130_fd_sc_hd__or2b_1 _3209_ (.A(_0570_),
    .B_N(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__o21a_1 _3210_ (.A1(_0564_),
    .A2(_0567_),
    .B1(_0565_),
    .X(_0573_));
 sky130_fd_sc_hd__xnor2_2 _3211_ (.A(_0572_),
    .B(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__o21ai_1 _3212_ (.A1(_0570_),
    .A2(_0573_),
    .B1(_0571_),
    .Y(_0575_));
 sky130_fd_sc_hd__o21bai_4 _3213_ (.A1(_0569_),
    .A2(_0574_),
    .B1_N(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__or3_1 _3214_ (.A(_0569_),
    .B(_0571_),
    .C(_0573_),
    .X(_0577_));
 sky130_fd_sc_hd__a31o_1 _3215_ (.A1(_0537_),
    .A2(_0576_),
    .A3(_0577_),
    .B1(_0535_),
    .X(_0578_));
 sky130_fd_sc_hd__xnor2_1 _3216_ (.A(_0534_),
    .B(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__a21boi_1 _3217_ (.A1(_0533_),
    .A2(_0578_),
    .B1_N(_0532_),
    .Y(_0580_));
 sky130_fd_sc_hd__nor2_1 _3218_ (.A(\game.addhits.a[10] ),
    .B(\game.addhits.add3.b[2] ),
    .Y(_0581_));
 sky130_fd_sc_hd__nand2_1 _3219_ (.A(\game.addhits.a[10] ),
    .B(\game.addhits.add3.b[2] ),
    .Y(_0582_));
 sky130_fd_sc_hd__and2b_1 _3220_ (.A_N(_0581_),
    .B(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__xnor2_1 _3221_ (.A(_0580_),
    .B(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__nor2_1 _3222_ (.A(_0579_),
    .B(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__nor2_1 _3223_ (.A(\game.addhits.a[11] ),
    .B(\game.addhits.add3.b[3] ),
    .Y(_0586_));
 sky130_fd_sc_hd__nand2_1 _3224_ (.A(\game.addhits.a[11] ),
    .B(\game.addhits.add3.b[3] ),
    .Y(_0587_));
 sky130_fd_sc_hd__or2b_1 _3225_ (.A(_0586_),
    .B_N(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__o21a_1 _3226_ (.A1(_0580_),
    .A2(_0581_),
    .B1(_0582_),
    .X(_0589_));
 sky130_fd_sc_hd__xnor2_1 _3227_ (.A(_0588_),
    .B(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__nor2_2 _3228_ (.A(_0585_),
    .B(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__o21ai_2 _3229_ (.A1(_0586_),
    .A2(_0589_),
    .B1(_0587_),
    .Y(_0592_));
 sky130_fd_sc_hd__xor2_2 _3230_ (.A(_0591_),
    .B(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__xor2_1 _3231_ (.A(_0531_),
    .B(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__a21oi_2 _3232_ (.A1(_0504_),
    .A2(_0528_),
    .B1(_0594_),
    .Y(_0595_));
 sky130_fd_sc_hd__nor2_1 _3233_ (.A(_0484_),
    .B(_0485_),
    .Y(_0596_));
 sky130_fd_sc_hd__xnor2_2 _3234_ (.A(_0443_),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__xor2_1 _3235_ (.A(_0487_),
    .B(_0500_),
    .X(_0598_));
 sky130_fd_sc_hd__a21oi_1 _3236_ (.A1(_0493_),
    .A2(_0499_),
    .B1(_0498_),
    .Y(_0599_));
 sky130_fd_sc_hd__a21oi_2 _3237_ (.A1(_0493_),
    .A2(_0498_),
    .B1(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__a21boi_1 _3238_ (.A1(_0492_),
    .A2(_0598_),
    .B1_N(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__and3_1 _3239_ (.A(_0537_),
    .B(_0576_),
    .C(_0577_),
    .X(_0602_));
 sky130_fd_sc_hd__a21oi_1 _3240_ (.A1(_0576_),
    .A2(_0577_),
    .B1(_0537_),
    .Y(_0603_));
 sky130_fd_sc_hd__nor2_1 _3241_ (.A(_0602_),
    .B(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__inv_2 _3242_ (.A(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__o21a_1 _3243_ (.A1(_0597_),
    .A2(_0601_),
    .B1(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__or2b_1 _3244_ (.A(_0563_),
    .B_N(_0576_),
    .X(_0607_));
 sky130_fd_sc_hd__a22o_2 _3245_ (.A1(_0569_),
    .A2(_0575_),
    .B1(_0607_),
    .B2(_0568_),
    .X(_0608_));
 sky130_fd_sc_hd__xnor2_2 _3246_ (.A(_0471_),
    .B(_0484_),
    .Y(_0609_));
 sky130_fd_sc_hd__nand2_1 _3247_ (.A(_0471_),
    .B(_0476_),
    .Y(_0610_));
 sky130_fd_sc_hd__inv_2 _3248_ (.A(_0483_),
    .Y(_0611_));
 sky130_fd_sc_hd__inv_2 _3249_ (.A(_0471_),
    .Y(_0612_));
 sky130_fd_sc_hd__nor2_1 _3250_ (.A(_0612_),
    .B(_0484_),
    .Y(_0613_));
 sky130_fd_sc_hd__o22a_1 _3251_ (.A1(_0610_),
    .A2(_0611_),
    .B1(_0613_),
    .B2(_0476_),
    .X(_0614_));
 sky130_fd_sc_hd__nand2_1 _3252_ (.A(_0476_),
    .B(_0609_),
    .Y(_0615_));
 sky130_fd_sc_hd__and2_1 _3253_ (.A(_0610_),
    .B(_0483_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_2 _3254_ (.A0(_0477_),
    .A1(_0616_),
    .S(_0482_),
    .X(_0617_));
 sky130_fd_sc_hd__inv_2 _3255_ (.A(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__o211a_1 _3256_ (.A1(_0609_),
    .A2(_0614_),
    .B1(_0615_),
    .C1(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__nand2_1 _3257_ (.A(_0608_),
    .B(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__or2_1 _3258_ (.A(_0608_),
    .B(_0619_),
    .X(_0621_));
 sky130_fd_sc_hd__nand2_1 _3259_ (.A(_0620_),
    .B(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__nor2_1 _3260_ (.A(_0553_),
    .B(_0559_),
    .Y(_0623_));
 sky130_fd_sc_hd__mux2_1 _3261_ (.A0(_0553_),
    .A1(_0623_),
    .S(_0558_),
    .X(_0624_));
 sky130_fd_sc_hd__inv_2 _3262_ (.A(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__or2_1 _3263_ (.A(_0461_),
    .B(_0467_),
    .X(_0626_));
 sky130_fd_sc_hd__nor2_1 _3264_ (.A(_0461_),
    .B(_0466_),
    .Y(_0627_));
 sky130_fd_sc_hd__a21o_1 _3265_ (.A1(_0466_),
    .A2(_0626_),
    .B1(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__xnor2_4 _3266_ (.A(_0454_),
    .B(_0468_),
    .Y(_0629_));
 sky130_fd_sc_hd__nor2_1 _3267_ (.A(_0460_),
    .B(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__nand2_1 _3268_ (.A(_0628_),
    .B(_0630_),
    .Y(_0631_));
 sky130_fd_sc_hd__xnor2_1 _3269_ (.A(_0624_),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__a21oi_4 _3270_ (.A1(_0466_),
    .A2(_0626_),
    .B1(_0627_),
    .Y(_0633_));
 sky130_fd_sc_hd__o21ai_4 _3271_ (.A1(_0460_),
    .A2(_0629_),
    .B1(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__or2_1 _3272_ (.A(\game.addmisses.add1.b[0] ),
    .B(\game.addmisses.a[0] ),
    .X(_0635_));
 sky130_fd_sc_hd__nand2_2 _3273_ (.A(_0450_),
    .B(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__or2_1 _3274_ (.A(\game.addhits.add1.b[0] ),
    .B(\game.addhits.a[0] ),
    .X(_0637_));
 sky130_fd_sc_hd__nand2_2 _3275_ (.A(_0544_),
    .B(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__inv_2 _3276_ (.A(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__a21oi_4 _3277_ (.A1(_0634_),
    .A2(_0636_),
    .B1(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__xor2_2 _3278_ (.A(_0454_),
    .B(_0468_),
    .X(_0641_));
 sky130_fd_sc_hd__xor2_4 _3279_ (.A(_0546_),
    .B(_0560_),
    .X(_0642_));
 sky130_fd_sc_hd__or3b_1 _3280_ (.A(_0633_),
    .B(_0641_),
    .C_N(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__a21o_1 _3281_ (.A1(_0628_),
    .A2(_0629_),
    .B1(_0642_),
    .X(_0644_));
 sky130_fd_sc_hd__nand2_1 _3282_ (.A(_0643_),
    .B(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__o21ai_1 _3283_ (.A1(_0640_),
    .A2(_0645_),
    .B1(_0643_),
    .Y(_0646_));
 sky130_fd_sc_hd__or2b_1 _3284_ (.A(_0546_),
    .B_N(_0560_),
    .X(_0647_));
 sky130_fd_sc_hd__and2b_1 _3285_ (.A_N(_0559_),
    .B(_0553_),
    .X(_0648_));
 sky130_fd_sc_hd__a21o_1 _3286_ (.A1(_0552_),
    .A2(_0647_),
    .B1(_0648_),
    .X(_0649_));
 sky130_fd_sc_hd__or2_1 _3287_ (.A(_0460_),
    .B(_0629_),
    .X(_0650_));
 sky130_fd_sc_hd__o21ai_1 _3288_ (.A1(_0454_),
    .A2(_0468_),
    .B1(_0460_),
    .Y(_0651_));
 sky130_fd_sc_hd__or3_1 _3289_ (.A(_0454_),
    .B(_0460_),
    .C(_0467_),
    .X(_0652_));
 sky130_fd_sc_hd__a21o_1 _3290_ (.A1(_0651_),
    .A2(_0652_),
    .B1(_0641_),
    .X(_0653_));
 sky130_fd_sc_hd__and3_1 _3291_ (.A(_0628_),
    .B(_0650_),
    .C(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__xor2_1 _3292_ (.A(_0649_),
    .B(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__and2_1 _3293_ (.A(_0649_),
    .B(_0654_),
    .X(_0656_));
 sky130_fd_sc_hd__a21o_1 _3294_ (.A1(_0646_),
    .A2(_0655_),
    .B1(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__nand2_1 _3295_ (.A(_0632_),
    .B(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__o21ai_1 _3296_ (.A1(_0625_),
    .A2(_0631_),
    .B1(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__xnor2_1 _3297_ (.A(_0632_),
    .B(_0657_),
    .Y(_0660_));
 sky130_fd_sc_hd__xnor2_2 _3298_ (.A(_0640_),
    .B(_0645_),
    .Y(_0661_));
 sky130_fd_sc_hd__xnor2_1 _3299_ (.A(_0646_),
    .B(_0655_),
    .Y(_0662_));
 sky130_fd_sc_hd__nand2_1 _3300_ (.A(_0661_),
    .B(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__and2b_1 _3301_ (.A_N(_0660_),
    .B(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__or2_2 _3302_ (.A(_0659_),
    .B(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__nor2_2 _3303_ (.A(_0468_),
    .B(_0469_),
    .Y(_0666_));
 sky130_fd_sc_hd__xnor2_4 _3304_ (.A(_0449_),
    .B(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__a21boi_1 _3305_ (.A1(_0476_),
    .A2(_0609_),
    .B1_N(_0617_),
    .Y(_0668_));
 sky130_fd_sc_hd__and3_1 _3306_ (.A(_0543_),
    .B(_0560_),
    .C(_0561_),
    .X(_0669_));
 sky130_fd_sc_hd__a21oi_1 _3307_ (.A1(_0560_),
    .A2(_0561_),
    .B1(_0543_),
    .Y(_0670_));
 sky130_fd_sc_hd__or2_2 _3308_ (.A(_0669_),
    .B(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__o21ai_1 _3309_ (.A1(_0667_),
    .A2(_0668_),
    .B1(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__or3_1 _3310_ (.A(_0671_),
    .B(_0667_),
    .C(_0668_),
    .X(_0673_));
 sky130_fd_sc_hd__a21bo_1 _3311_ (.A1(_0665_),
    .A2(_0672_),
    .B1_N(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__xor2_4 _3312_ (.A(_0563_),
    .B(_0576_),
    .X(_0675_));
 sky130_fd_sc_hd__nor2_1 _3313_ (.A(_0617_),
    .B(_0609_),
    .Y(_0676_));
 sky130_fd_sc_hd__or2_1 _3314_ (.A(_0675_),
    .B(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__and2_1 _3315_ (.A(_0675_),
    .B(_0676_),
    .X(_0678_));
 sky130_fd_sc_hd__a21oi_2 _3316_ (.A1(_0674_),
    .A2(_0677_),
    .B1(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__xor2_2 _3317_ (.A(_0622_),
    .B(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__and2b_1 _3318_ (.A_N(_0678_),
    .B(_0677_),
    .X(_0681_));
 sky130_fd_sc_hd__xnor2_2 _3319_ (.A(_0674_),
    .B(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__and2b_1 _3320_ (.A_N(_0680_),
    .B(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__o21ai_1 _3321_ (.A1(_0622_),
    .A2(_0679_),
    .B1(_0620_),
    .Y(_0684_));
 sky130_fd_sc_hd__and2b_1 _3322_ (.A_N(_0569_),
    .B(_0575_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _3323_ (.A0(_0569_),
    .A1(_0685_),
    .S(_0574_),
    .X(_0686_));
 sky130_fd_sc_hd__nor2_1 _3324_ (.A(_0617_),
    .B(_0615_),
    .Y(_0687_));
 sky130_fd_sc_hd__and2_1 _3325_ (.A(_0686_),
    .B(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__or2_1 _3326_ (.A(_0686_),
    .B(_0687_),
    .X(_0689_));
 sky130_fd_sc_hd__and2b_1 _3327_ (.A_N(_0688_),
    .B(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__xnor2_1 _3328_ (.A(_0684_),
    .B(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__a21o_1 _3329_ (.A1(_0684_),
    .A2(_0689_),
    .B1(_0688_),
    .X(_0692_));
 sky130_fd_sc_hd__o21ba_2 _3330_ (.A1(_0683_),
    .A2(_0691_),
    .B1_N(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__or3_1 _3331_ (.A(_0605_),
    .B(_0597_),
    .C(_0601_),
    .X(_0694_));
 sky130_fd_sc_hd__o21ai_1 _3332_ (.A1(_0606_),
    .A2(_0693_),
    .B1(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__nor2_1 _3333_ (.A(_0591_),
    .B(_0592_),
    .Y(_0696_));
 sky130_fd_sc_hd__xnor2_1 _3334_ (.A(_0579_),
    .B(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__nor2_1 _3335_ (.A(_0600_),
    .B(_0598_),
    .Y(_0698_));
 sky130_fd_sc_hd__and2_1 _3336_ (.A(_0697_),
    .B(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__nor2_1 _3337_ (.A(_0697_),
    .B(_0698_),
    .Y(_0700_));
 sky130_fd_sc_hd__nor2_1 _3338_ (.A(_0699_),
    .B(_0700_),
    .Y(_0701_));
 sky130_fd_sc_hd__xor2_1 _3339_ (.A(_0695_),
    .B(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__or2_1 _3340_ (.A(_0579_),
    .B(_0696_),
    .X(_0703_));
 sky130_fd_sc_hd__a22o_1 _3341_ (.A1(_0585_),
    .A2(_0592_),
    .B1(_0703_),
    .B2(_0584_),
    .X(_0704_));
 sky130_fd_sc_hd__or2_1 _3342_ (.A(_0487_),
    .B(_0500_),
    .X(_0705_));
 sky130_fd_sc_hd__xnor2_1 _3343_ (.A(_0492_),
    .B(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__nor2_1 _3344_ (.A(_0600_),
    .B(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__xnor2_2 _3345_ (.A(_0704_),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__a21o_1 _3346_ (.A1(_0695_),
    .A2(_0701_),
    .B1(_0699_),
    .X(_0709_));
 sky130_fd_sc_hd__xnor2_1 _3347_ (.A(_0708_),
    .B(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__or2_2 _3348_ (.A(_0702_),
    .B(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__inv_2 _3349_ (.A(_0708_),
    .Y(_0712_));
 sky130_fd_sc_hd__and2_1 _3350_ (.A(_0704_),
    .B(_0707_),
    .X(_0713_));
 sky130_fd_sc_hd__a21o_1 _3351_ (.A1(_0712_),
    .A2(_0709_),
    .B1(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__or2b_1 _3352_ (.A(_0585_),
    .B_N(_0592_),
    .X(_0715_));
 sky130_fd_sc_hd__a21o_1 _3353_ (.A1(_0590_),
    .A2(_0715_),
    .B1(_0591_),
    .X(_0716_));
 sky130_fd_sc_hd__nand3b_1 _3354_ (.A_N(_0600_),
    .B(_0598_),
    .C(_0492_),
    .Y(_0717_));
 sky130_fd_sc_hd__nor2_1 _3355_ (.A(_0716_),
    .B(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__and2_1 _3356_ (.A(_0716_),
    .B(_0717_),
    .X(_0719_));
 sky130_fd_sc_hd__nor2_1 _3357_ (.A(_0718_),
    .B(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__xor2_2 _3358_ (.A(_0714_),
    .B(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__a21o_1 _3359_ (.A1(_0714_),
    .A2(_0720_),
    .B1(_0718_),
    .X(_0722_));
 sky130_fd_sc_hd__a21oi_4 _3360_ (.A1(_0711_),
    .A2(_0721_),
    .B1(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__and3_1 _3361_ (.A(_0594_),
    .B(_0504_),
    .C(_0528_),
    .X(_0724_));
 sky130_fd_sc_hd__o21bai_4 _3362_ (.A1(_0595_),
    .A2(_0723_),
    .B1_N(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__nand2_1 _3363_ (.A(\game.addhits.a[13] ),
    .B(\game.addhits.add4.b[1] ),
    .Y(_0726_));
 sky130_fd_sc_hd__or2_1 _3364_ (.A(\game.addhits.a[13] ),
    .B(\game.addhits.add4.b[1] ),
    .X(_0727_));
 sky130_fd_sc_hd__nand2_1 _3365_ (.A(_0726_),
    .B(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__a21oi_2 _3366_ (.A1(_0531_),
    .A2(_0593_),
    .B1(_0529_),
    .Y(_0729_));
 sky130_fd_sc_hd__xnor2_2 _3367_ (.A(_0728_),
    .B(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__o21a_1 _3368_ (.A1(_0728_),
    .A2(_0729_),
    .B1(_0726_),
    .X(_0731_));
 sky130_fd_sc_hd__nor2_1 _3369_ (.A(\game.addhits.a[14] ),
    .B(\game.addhits.add4.b[2] ),
    .Y(_0732_));
 sky130_fd_sc_hd__nand2_1 _3370_ (.A(\game.addhits.a[14] ),
    .B(\game.addhits.add4.b[2] ),
    .Y(_0733_));
 sky130_fd_sc_hd__o21ai_1 _3371_ (.A1(_0731_),
    .A2(_0732_),
    .B1(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__o21ai_1 _3372_ (.A1(\game.addhits.a[15] ),
    .A2(\game.addhits.add4.b[3] ),
    .B1(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__or2_1 _3373_ (.A(\game.addhits.a[14] ),
    .B(\game.addhits.add4.b[2] ),
    .X(_0736_));
 sky130_fd_sc_hd__nand2_1 _3374_ (.A(_0733_),
    .B(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__xnor2_2 _3375_ (.A(_0731_),
    .B(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__nand2_1 _3376_ (.A(_0738_),
    .B(_0730_),
    .Y(_0739_));
 sky130_fd_sc_hd__nor2_1 _3377_ (.A(\game.addhits.a[15] ),
    .B(\game.addhits.add4.b[3] ),
    .Y(_0740_));
 sky130_fd_sc_hd__inv_2 _3378_ (.A(\game.addhits.a[15] ),
    .Y(_0741_));
 sky130_fd_sc_hd__inv_2 _3379_ (.A(\game.addhits.add4.b[3] ),
    .Y(_0742_));
 sky130_fd_sc_hd__nor2_1 _3380_ (.A(_0741_),
    .B(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__or2_1 _3381_ (.A(_0740_),
    .B(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__xnor2_1 _3382_ (.A(_0734_),
    .B(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__a21oi_1 _3383_ (.A1(_0739_),
    .A2(_0745_),
    .B1(_0743_),
    .Y(_0746_));
 sky130_fd_sc_hd__and2_1 _3384_ (.A(_0735_),
    .B(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__xor2_1 _3385_ (.A(_0730_),
    .B(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__and3_1 _3386_ (.A(_0527_),
    .B(_0748_),
    .C(_0524_),
    .X(_0749_));
 sky130_fd_sc_hd__a21o_1 _3387_ (.A1(_0527_),
    .A2(_0524_),
    .B1(_0748_),
    .X(_0750_));
 sky130_fd_sc_hd__and2b_1 _3388_ (.A_N(_0749_),
    .B(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__xnor2_4 _3389_ (.A(_0725_),
    .B(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__a21boi_1 _3390_ (.A1(_0735_),
    .A2(_0746_),
    .B1_N(_0730_),
    .Y(_0753_));
 sky130_fd_sc_hd__xnor2_1 _3391_ (.A(_0738_),
    .B(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__nand2_1 _3392_ (.A(_0514_),
    .B(_0523_),
    .Y(_0755_));
 sky130_fd_sc_hd__xnor2_1 _3393_ (.A(_0512_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__and2_1 _3394_ (.A(_0527_),
    .B(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__nor2_1 _3395_ (.A(_0754_),
    .B(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__nand2_1 _3396_ (.A(_0754_),
    .B(_0757_),
    .Y(_0759_));
 sky130_fd_sc_hd__or2b_2 _3397_ (.A(_0758_),
    .B_N(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__a21oi_4 _3398_ (.A1(_0725_),
    .A2(_0750_),
    .B1(_0749_),
    .Y(_0761_));
 sky130_fd_sc_hd__xnor2_4 _3399_ (.A(_0760_),
    .B(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__nand2_2 _3400_ (.A(_0762_),
    .B(_0752_),
    .Y(_0763_));
 sky130_fd_sc_hd__o21ai_4 _3401_ (.A1(_0758_),
    .A2(_0761_),
    .B1(_0759_),
    .Y(_0764_));
 sky130_fd_sc_hd__a21o_1 _3402_ (.A1(_0738_),
    .A2(_0730_),
    .B1(_0747_),
    .X(_0765_));
 sky130_fd_sc_hd__mux2_1 _3403_ (.A0(_0765_),
    .A1(_0739_),
    .S(_0745_),
    .X(_0766_));
 sky130_fd_sc_hd__or3b_2 _3404_ (.A(_0512_),
    .B(_0524_),
    .C_N(_0527_),
    .X(_0767_));
 sky130_fd_sc_hd__and2_1 _3405_ (.A(_0766_),
    .B(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__nor2_1 _3406_ (.A(_0766_),
    .B(_0767_),
    .Y(_0769_));
 sky130_fd_sc_hd__nor2_2 _3407_ (.A(_0768_),
    .B(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__xor2_4 _3408_ (.A(_0764_),
    .B(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__a21o_1 _3409_ (.A1(_0764_),
    .A2(_0770_),
    .B1(_0769_),
    .X(_0772_));
 sky130_fd_sc_hd__a21o_1 _3410_ (.A1(_0763_),
    .A2(_0771_),
    .B1(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__inv_2 _3411_ (.A(_0762_),
    .Y(_0774_));
 sky130_fd_sc_hd__a21o_1 _3412_ (.A1(_0752_),
    .A2(_0773_),
    .B1(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__a211o_1 _3413_ (.A1(_0763_),
    .A2(_0771_),
    .B1(_0772_),
    .C1(_0752_),
    .X(_0776_));
 sky130_fd_sc_hd__and2_1 _3414_ (.A(_0763_),
    .B(_0771_),
    .X(_0777_));
 sky130_fd_sc_hd__a21oi_2 _3415_ (.A1(_0763_),
    .A2(_0772_),
    .B1(_0771_),
    .Y(_0778_));
 sky130_fd_sc_hd__inv_2 _3416_ (.A(_0683_),
    .Y(_0779_));
 sky130_fd_sc_hd__and2_1 _3417_ (.A(_0692_),
    .B(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__mux2_2 _3418_ (.A0(_0683_),
    .A1(_0780_),
    .S(_0691_),
    .X(_0781_));
 sky130_fd_sc_hd__and3_1 _3419_ (.A(_0673_),
    .B(_0665_),
    .C(_0672_),
    .X(_0782_));
 sky130_fd_sc_hd__a21oi_1 _3420_ (.A1(_0673_),
    .A2(_0672_),
    .B1(_0665_),
    .Y(_0783_));
 sky130_fd_sc_hd__nor2_1 _3421_ (.A(_0782_),
    .B(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__nand2_1 _3422_ (.A(_0659_),
    .B(_0663_),
    .Y(_0785_));
 sky130_fd_sc_hd__a21o_1 _3423_ (.A1(_0660_),
    .A2(_0785_),
    .B1(_0664_),
    .X(_0786_));
 sky130_fd_sc_hd__nor2_1 _3424_ (.A(_0661_),
    .B(_0665_),
    .Y(_0787_));
 sky130_fd_sc_hd__a21bo_1 _3425_ (.A1(_0661_),
    .A2(_0665_),
    .B1_N(_0662_),
    .X(_0788_));
 sky130_fd_sc_hd__nor2_1 _3426_ (.A(_0787_),
    .B(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__nor2_1 _3427_ (.A(_0786_),
    .B(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__xnor2_2 _3428_ (.A(_0682_),
    .B(_0693_),
    .Y(_0791_));
 sky130_fd_sc_hd__inv_2 _3429_ (.A(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__or2_1 _3430_ (.A(_0680_),
    .B(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__a21o_1 _3431_ (.A1(_0784_),
    .A2(_0790_),
    .B1(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__a221o_1 _3432_ (.A1(_0702_),
    .A2(_0723_),
    .B1(_0781_),
    .B2(_0794_),
    .C1(_0710_),
    .X(_0795_));
 sky130_fd_sc_hd__o21bai_1 _3433_ (.A1(_0702_),
    .A2(_0723_),
    .B1_N(_0795_),
    .Y(_0796_));
 sky130_fd_sc_hd__or2_1 _3434_ (.A(_0724_),
    .B(_0595_),
    .X(_0797_));
 sky130_fd_sc_hd__xnor2_1 _3435_ (.A(_0797_),
    .B(_0723_),
    .Y(_0798_));
 sky130_fd_sc_hd__o21ai_1 _3436_ (.A1(_0597_),
    .A2(_0601_),
    .B1(_0605_),
    .Y(_0799_));
 sky130_fd_sc_hd__and2_1 _3437_ (.A(_0694_),
    .B(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__xnor2_1 _3438_ (.A(_0800_),
    .B(_0693_),
    .Y(_0801_));
 sky130_fd_sc_hd__a21oi_1 _3439_ (.A1(_0722_),
    .A2(_0711_),
    .B1(_0721_),
    .Y(_0802_));
 sky130_fd_sc_hd__a21oi_1 _3440_ (.A1(_0711_),
    .A2(_0721_),
    .B1(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__or2_1 _3441_ (.A(_0781_),
    .B(_0793_),
    .X(_0804_));
 sky130_fd_sc_hd__and3_1 _3442_ (.A(_0544_),
    .B(_0637_),
    .C(_0636_),
    .X(_0805_));
 sky130_fd_sc_hd__a21oi_4 _3443_ (.A1(_0634_),
    .A2(_0805_),
    .B1(_0640_),
    .Y(_0806_));
 sky130_fd_sc_hd__and2_1 _3444_ (.A(_0786_),
    .B(_0789_),
    .X(_0807_));
 sky130_fd_sc_hd__nand2_1 _3445_ (.A(_0806_),
    .B(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__or3_1 _3446_ (.A(_0784_),
    .B(_0804_),
    .C(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__and4b_1 _3447_ (.A_N(_0798_),
    .B(_0801_),
    .C(_0803_),
    .D(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__nor4b_1 _3448_ (.A(_0777_),
    .B(_0778_),
    .C(_0796_),
    .D_N(_0810_),
    .Y(_0811_));
 sky130_fd_sc_hd__a21o_1 _3449_ (.A1(_0781_),
    .A2(_0793_),
    .B1(_0784_),
    .X(_0812_));
 sky130_fd_sc_hd__or2_1 _3450_ (.A(_0808_),
    .B(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__or3_2 _3451_ (.A(_0781_),
    .B(_0791_),
    .C(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__inv_2 _3452_ (.A(_0693_),
    .Y(_0815_));
 sky130_fd_sc_hd__nand2_1 _3453_ (.A(_0682_),
    .B(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__a22oi_2 _3454_ (.A1(_0692_),
    .A2(_0683_),
    .B1(_0816_),
    .B2(_0680_),
    .Y(_0817_));
 sky130_fd_sc_hd__o21ai_1 _3455_ (.A1(_0791_),
    .A2(_0817_),
    .B1(_0793_),
    .Y(_0818_));
 sky130_fd_sc_hd__nor2_1 _3456_ (.A(_0781_),
    .B(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__xnor2_1 _3457_ (.A(_0814_),
    .B(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__and4b_1 _3458_ (.A_N(_0775_),
    .B(_0776_),
    .C(net43),
    .D(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__inv_2 _3459_ (.A(_0752_),
    .Y(_0822_));
 sky130_fd_sc_hd__a21oi_2 _3460_ (.A1(_0763_),
    .A2(_0771_),
    .B1(_0772_),
    .Y(_0823_));
 sky130_fd_sc_hd__nor2_2 _3461_ (.A(_0822_),
    .B(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__and2_2 _3462_ (.A(_0776_),
    .B(_0798_),
    .X(_0825_));
 sky130_fd_sc_hd__o32a_4 _3463_ (.A1(_0774_),
    .A2(_0822_),
    .A3(_0823_),
    .B1(_0778_),
    .B2(_0777_),
    .X(_0826_));
 sky130_fd_sc_hd__inv_2 _3464_ (.A(_0817_),
    .Y(_0827_));
 sky130_fd_sc_hd__o311a_1 _3465_ (.A1(_0762_),
    .A2(_0824_),
    .A3(_0825_),
    .B1(_0826_),
    .C1(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__o31a_1 _3466_ (.A1(_0762_),
    .A2(_0824_),
    .A3(_0825_),
    .B1(_0826_),
    .X(_0829_));
 sky130_fd_sc_hd__clkbuf_4 _3467_ (.A(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__nor2_1 _3468_ (.A(_0752_),
    .B(_0773_),
    .Y(_0831_));
 sky130_fd_sc_hd__or4b_1 _3469_ (.A(_0796_),
    .B(_0801_),
    .C(_0803_),
    .D_N(_0798_),
    .X(_0832_));
 sky130_fd_sc_hd__or3_1 _3470_ (.A(_0775_),
    .B(_0831_),
    .C(_0832_),
    .X(_0833_));
 sky130_fd_sc_hd__buf_2 _3471_ (.A(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__a2bb2o_1 _3472_ (.A1_N(_0821_),
    .A2_N(_0828_),
    .B1(_0830_),
    .B2(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__o21ai_1 _3473_ (.A1(_0781_),
    .A2(_0791_),
    .B1(_0813_),
    .Y(_0836_));
 sky130_fd_sc_hd__and3_1 _3474_ (.A(_0804_),
    .B(_0814_),
    .C(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__and4b_1 _3475_ (.A_N(_0775_),
    .B(_0776_),
    .C(_0811_),
    .D(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__o311a_1 _3476_ (.A1(_0762_),
    .A2(_0824_),
    .A3(_0825_),
    .B1(_0826_),
    .C1(_0792_),
    .X(_0839_));
 sky130_fd_sc_hd__a2bb2o_2 _3477_ (.A1_N(_0838_),
    .A2_N(_0839_),
    .B1(_0830_),
    .B2(_0834_),
    .X(_0840_));
 sky130_fd_sc_hd__nand2_1 _3478_ (.A(_0830_),
    .B(_0834_),
    .Y(_0841_));
 sky130_fd_sc_hd__o31ai_4 _3479_ (.A1(_0762_),
    .A2(_0824_),
    .A3(_0825_),
    .B1(_0826_),
    .Y(_0842_));
 sky130_fd_sc_hd__o31ai_1 _3480_ (.A1(_0781_),
    .A2(_0814_),
    .A3(_0818_),
    .B1(_0804_),
    .Y(_0843_));
 sky130_fd_sc_hd__or4b_2 _3481_ (.A(_0777_),
    .B(_0778_),
    .C(_0796_),
    .D_N(_0810_),
    .X(_0844_));
 sky130_fd_sc_hd__a2111o_1 _3482_ (.A1(_0809_),
    .A2(_0843_),
    .B1(_0844_),
    .C1(_0775_),
    .D1(_0831_),
    .X(_0845_));
 sky130_fd_sc_hd__o311a_1 _3483_ (.A1(_0762_),
    .A2(_0824_),
    .A3(_0825_),
    .B1(_0826_),
    .C1(_0781_),
    .X(_0846_));
 sky130_fd_sc_hd__a21oi_2 _3484_ (.A1(net42),
    .A2(_0845_),
    .B1(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__and2_1 _3485_ (.A(_0841_),
    .B(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__o21ai_1 _3486_ (.A1(_0835_),
    .A2(_0840_),
    .B1(_0848_),
    .Y(_0849_));
 sky130_fd_sc_hd__and3_1 _3487_ (.A(_0841_),
    .B(_0847_),
    .C(_0835_),
    .X(_0850_));
 sky130_fd_sc_hd__nand2_1 _3488_ (.A(_0808_),
    .B(_0812_),
    .Y(_0851_));
 sky130_fd_sc_hd__a2111oi_1 _3489_ (.A1(_0813_),
    .A2(_0851_),
    .B1(_0775_),
    .C1(_0831_),
    .D1(_0844_),
    .Y(_0852_));
 sky130_fd_sc_hd__inv_2 _3490_ (.A(_0784_),
    .Y(_0853_));
 sky130_fd_sc_hd__o311a_1 _3491_ (.A1(_0762_),
    .A2(_0824_),
    .A3(_0825_),
    .B1(_0826_),
    .C1(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__o2bb2a_2 _3492_ (.A1_N(_0830_),
    .A2_N(_0834_),
    .B1(net40),
    .B2(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__and3_1 _3493_ (.A(_0840_),
    .B(_0850_),
    .C(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__and2_1 _3494_ (.A(_0830_),
    .B(_0834_),
    .X(_0857_));
 sky130_fd_sc_hd__o2bb2a_1 _3495_ (.A1_N(_0830_),
    .A2_N(_0834_),
    .B1(_0821_),
    .B2(_0828_),
    .X(_0858_));
 sky130_fd_sc_hd__or3b_1 _3496_ (.A(_0857_),
    .B(_0858_),
    .C_N(_0847_),
    .X(_0859_));
 sky130_fd_sc_hd__or3b_1 _3497_ (.A(_0855_),
    .B(_0835_),
    .C_N(_0840_),
    .X(_0860_));
 sky130_fd_sc_hd__o21ai_1 _3498_ (.A1(_0840_),
    .A2(_0859_),
    .B1(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__o211a_1 _3499_ (.A1(\game.flash_counter[6] ),
    .A2(\game.flash_counter[7] ),
    .B1(\game.flash_counter[9] ),
    .C1(\game.flash_counter[8] ),
    .X(_0862_));
 sky130_fd_sc_hd__o21a_1 _3500_ (.A1(\game.flash_counter[10] ),
    .A2(_0862_),
    .B1(\game.flash_counter[11] ),
    .X(_0863_));
 sky130_fd_sc_hd__o31a_1 _3501_ (.A1(\game.flash_counter[12] ),
    .A2(\game.flash_counter[13] ),
    .A3(_0863_),
    .B1(\game.flash_counter[14] ),
    .X(_0864_));
 sky130_fd_sc_hd__or4_1 _3502_ (.A(\game.flash_counter[17] ),
    .B(\game.flash_counter[16] ),
    .C(\game.flash_counter[15] ),
    .D(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__a31o_1 _3503_ (.A1(\game.flash_counter[19] ),
    .A2(\game.flash_counter[18] ),
    .A3(_0865_),
    .B1(\game.flash_counter[21] ),
    .X(_0866_));
 sky130_fd_sc_hd__o21a_1 _3504_ (.A1(\game.flash_counter[20] ),
    .A2(_0866_),
    .B1(\game.flash_counter[22] ),
    .X(_0867_));
 sky130_fd_sc_hd__and3_1 _3505_ (.A(\game.flash_counter[3] ),
    .B(\game.flash_counter[2] ),
    .C(\game.flash_counter[4] ),
    .X(_0868_));
 sky130_fd_sc_hd__and3_1 _3506_ (.A(\game.flash_counter[1] ),
    .B(\game.flash_counter[0] ),
    .C(\game.flash_counter[5] ),
    .X(_0869_));
 sky130_fd_sc_hd__and3_1 _3507_ (.A(\game.flash_counter[9] ),
    .B(\game.flash_counter[8] ),
    .C(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__nand2_1 _3508_ (.A(\game.flash_counter[19] ),
    .B(\game.flash_counter[18] ),
    .Y(_0871_));
 sky130_fd_sc_hd__or4_1 _3509_ (.A(\game.flash_counter[17] ),
    .B(\game.flash_counter[16] ),
    .C(\game.flash_counter[6] ),
    .D(\game.flash_counter[7] ),
    .X(_0872_));
 sky130_fd_sc_hd__or4_1 _3510_ (.A(\game.flash_counter[20] ),
    .B(\game.flash_counter[21] ),
    .C(_0871_),
    .D(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__or4bb_1 _3511_ (.A(\game.flash_counter[15] ),
    .B(\game.flash_counter[12] ),
    .C_N(\game.flash_counter[14] ),
    .D_N(\game.flash_counter[22] ),
    .X(_0874_));
 sky130_fd_sc_hd__or4b_1 _3512_ (.A(\game.flash_counter[13] ),
    .B(\game.flash_counter[10] ),
    .C(_0874_),
    .D_N(\game.flash_counter[11] ),
    .X(_0875_));
 sky130_fd_sc_hd__nor2_1 _3513_ (.A(_0873_),
    .B(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__and3_1 _3514_ (.A(_0868_),
    .B(_0870_),
    .C(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__o31ai_1 _3515_ (.A1(\game.flash_counter[23] ),
    .A2(_0867_),
    .A3(_0877_),
    .B1(_0842_),
    .Y(_0878_));
 sky130_fd_sc_hd__nor2_2 _3516_ (.A(_0209_),
    .B(\modetrans.mode[4] ),
    .Y(_0879_));
 sky130_fd_sc_hd__or2_1 _3517_ (.A(_0552_),
    .B(_0642_),
    .X(_0880_));
 sky130_fd_sc_hd__and3b_1 _3518_ (.A_N(_0671_),
    .B(_0624_),
    .C(_0880_),
    .X(_0881_));
 sky130_fd_sc_hd__o31a_1 _3519_ (.A1(_0608_),
    .A2(_0675_),
    .A3(_0881_),
    .B1(_0686_),
    .X(_0882_));
 sky130_fd_sc_hd__or4b_1 _3520_ (.A(_0697_),
    .B(_0604_),
    .C(_0882_),
    .D_N(_0716_),
    .X(_0883_));
 sky130_fd_sc_hd__or4_1 _3521_ (.A(_0748_),
    .B(_0594_),
    .C(_0704_),
    .D(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__nor3b_1 _3522_ (.A(_0754_),
    .B(_0884_),
    .C_N(_0766_),
    .Y(_0885_));
 sky130_fd_sc_hd__nand2b_1 _3523_ (.A_N(_0686_),
    .B(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__a21oi_1 _3524_ (.A1(_0608_),
    .A2(_0675_),
    .B1(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__or2b_1 _3525_ (.A(_0675_),
    .B_N(_0671_),
    .X(_0888_));
 sky130_fd_sc_hd__nor2_1 _3526_ (.A(_0608_),
    .B(_0886_),
    .Y(_0889_));
 sky130_fd_sc_hd__or2b_1 _3527_ (.A(_0886_),
    .B_N(_0608_),
    .X(_0890_));
 sky130_fd_sc_hd__nor2_1 _3528_ (.A(_0675_),
    .B(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__a21o_1 _3529_ (.A1(_0675_),
    .A2(_0889_),
    .B1(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__nor3_1 _3530_ (.A(_0608_),
    .B(_0886_),
    .C(_0888_),
    .Y(_0893_));
 sky130_fd_sc_hd__a21oi_1 _3531_ (.A1(_0888_),
    .A2(_0892_),
    .B1(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__inv_2 _3532_ (.A(_0258_),
    .Y(_0895_));
 sky130_fd_sc_hd__or2_2 _3533_ (.A(_0255_),
    .B(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__a21o_1 _3534_ (.A1(_0887_),
    .A2(_0894_),
    .B1(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__inv_2 _3535_ (.A(\highest_score.highest_score[5] ),
    .Y(_0898_));
 sky130_fd_sc_hd__inv_2 _3536_ (.A(net152),
    .Y(_0899_));
 sky130_fd_sc_hd__nand2_1 _3537_ (.A(_0899_),
    .B(\highest_score.highest_score[6] ),
    .Y(_0900_));
 sky130_fd_sc_hd__or3_1 _3538_ (.A(_0899_),
    .B(\highest_score.highest_score[6] ),
    .C(\highest_score.highest_score[5] ),
    .X(_0901_));
 sky130_fd_sc_hd__o21a_1 _3539_ (.A1(_0898_),
    .A2(_0900_),
    .B1(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__o31ai_1 _3540_ (.A1(\highest_score.highest_score[6] ),
    .A2(\highest_score.highest_score[5] ),
    .A3(\highest_score.highest_score[4] ),
    .B1(_0899_),
    .Y(_0903_));
 sky130_fd_sc_hd__nand2_1 _3541_ (.A(_0901_),
    .B(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__or3b_1 _3542_ (.A(_0900_),
    .B(\highest_score.highest_score[5] ),
    .C_N(\highest_score.highest_score[4] ),
    .X(_0905_));
 sky130_fd_sc_hd__or3_2 _3543_ (.A(\highest_score.highest_score[7] ),
    .B(\highest_score.highest_score[6] ),
    .C(_0898_),
    .X(_0906_));
 sky130_fd_sc_hd__and4_1 _3544_ (.A(_0255_),
    .B(_0904_),
    .C(_0905_),
    .D(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__a21o_1 _3545_ (.A1(_0902_),
    .A2(_0907_),
    .B1(_0258_),
    .X(_0908_));
 sky130_fd_sc_hd__a31o_2 _3546_ (.A1(_0612_),
    .A2(_0482_),
    .A3(_0611_),
    .B1(_0613_),
    .X(_0909_));
 sky130_fd_sc_hd__a31o_1 _3547_ (.A1(_0667_),
    .A2(_0633_),
    .A3(_0650_),
    .B1(_0615_),
    .X(_0910_));
 sky130_fd_sc_hd__a21o_1 _3548_ (.A1(_0617_),
    .A2(_0910_),
    .B1(_0597_),
    .X(_0911_));
 sky130_fd_sc_hd__or4b_4 _3549_ (.A(_0717_),
    .B(_0767_),
    .C(_0911_),
    .D_N(_0504_),
    .X(_0912_));
 sky130_fd_sc_hd__and3b_1 _3550_ (.A_N(_0912_),
    .B(_0618_),
    .C(_0614_),
    .X(_0913_));
 sky130_fd_sc_hd__or2_1 _3551_ (.A(_0617_),
    .B(_0912_),
    .X(_0914_));
 sky130_fd_sc_hd__nor3_1 _3552_ (.A(_0909_),
    .B(_0614_),
    .C(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__a22o_1 _3553_ (.A1(_0909_),
    .A2(_0913_),
    .B1(_0915_),
    .B2(_0667_),
    .X(_0916_));
 sky130_fd_sc_hd__and2_1 _3554_ (.A(_0609_),
    .B(_0667_),
    .X(_0917_));
 sky130_fd_sc_hd__a21o_1 _3555_ (.A1(_0909_),
    .A2(_0913_),
    .B1(_0915_),
    .X(_0918_));
 sky130_fd_sc_hd__a21oi_1 _3556_ (.A1(_0913_),
    .A2(_0917_),
    .B1(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__o21ai_1 _3557_ (.A1(_0916_),
    .A2(_0919_),
    .B1(_0261_),
    .Y(_0920_));
 sky130_fd_sc_hd__inv_2 _3558_ (.A(\modetrans.mode[3] ),
    .Y(_0921_));
 sky130_fd_sc_hd__a31o_1 _3559_ (.A1(_0897_),
    .A2(_0908_),
    .A3(_0920_),
    .B1(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__nand2_1 _3560_ (.A(_0879_),
    .B(_0922_),
    .Y(_0923_));
 sky130_fd_sc_hd__o311a_1 _3561_ (.A1(_0849_),
    .A2(_0856_),
    .A3(_0861_),
    .B1(net39),
    .C1(_0923_),
    .X(_0924_));
 sky130_fd_sc_hd__buf_4 _3562_ (.A(\disp_song.mi6.in[4] ),
    .X(_0925_));
 sky130_fd_sc_hd__clkbuf_4 _3563_ (.A(\disp_song.mi6.in[1] ),
    .X(_0926_));
 sky130_fd_sc_hd__o21a_1 _3564_ (.A1(\disp_song.mi6.in[2] ),
    .A2(_0926_),
    .B1(\disp_song.mi6.in[3] ),
    .X(_0927_));
 sky130_fd_sc_hd__nor2_1 _3565_ (.A(_0925_),
    .B(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__o21ai_1 _3566_ (.A1(\disp_song.mi6.in[3] ),
    .A2(\disp_song.mi6.in[2] ),
    .B1(_0925_),
    .Y(_0929_));
 sky130_fd_sc_hd__nor2_1 _3567_ (.A(_0352_),
    .B(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__a21o_1 _3568_ (.A1(_0214_),
    .A2(_0928_),
    .B1(_0930_),
    .X(_0931_));
 sky130_fd_sc_hd__nor2_1 _3569_ (.A(_0259_),
    .B(_0922_),
    .Y(_0932_));
 sky130_fd_sc_hd__inv_12 _3570_ (.A(net5),
    .Y(_0933_));
 sky130_fd_sc_hd__o41a_1 _3571_ (.A1(_2654_),
    .A2(\modetrans.mode[5] ),
    .A3(\modetrans.mode[3] ),
    .A4(_0210_),
    .B1(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__buf_4 _3572_ (.A(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__o31a_1 _3573_ (.A1(_0924_),
    .A2(_0931_),
    .A3(_0932_),
    .B1(_0935_),
    .X(net23));
 sky130_fd_sc_hd__nor2_1 _3574_ (.A(_0667_),
    .B(_0912_),
    .Y(_0936_));
 sky130_fd_sc_hd__a21oi_1 _3575_ (.A1(_0909_),
    .A2(_0936_),
    .B1(_0917_),
    .Y(_0937_));
 sky130_fd_sc_hd__o31a_1 _3576_ (.A1(_0614_),
    .A2(_0914_),
    .A3(_0937_),
    .B1(_0261_),
    .X(_0938_));
 sky130_fd_sc_hd__nand2_1 _3577_ (.A(_0671_),
    .B(net44),
    .Y(_0939_));
 sky130_fd_sc_hd__mux2_1 _3578_ (.A0(_0671_),
    .A1(_0939_),
    .S(_0675_),
    .X(_0940_));
 sky130_fd_sc_hd__nor2_2 _3579_ (.A(_0255_),
    .B(_0895_),
    .Y(_0941_));
 sky130_fd_sc_hd__o21a_1 _3580_ (.A1(_0890_),
    .A2(_0940_),
    .B1(_0941_),
    .X(_0942_));
 sky130_fd_sc_hd__a21oi_1 _3581_ (.A1(\highest_score.highest_score[5] ),
    .A2(\highest_score.highest_score[4] ),
    .B1(_0900_),
    .Y(_0943_));
 sky130_fd_sc_hd__o211a_1 _3582_ (.A1(\highest_score.highest_score[5] ),
    .A2(\highest_score.highest_score[4] ),
    .B1(_0255_),
    .C1(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__nor2_1 _3583_ (.A(_0258_),
    .B(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hd__a2bb2o_1 _3584_ (.A1_N(net40),
    .A2_N(_0854_),
    .B1(_0830_),
    .B2(_0834_),
    .X(_0946_));
 sky130_fd_sc_hd__xnor2_1 _3585_ (.A(_0840_),
    .B(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__nand2_1 _3586_ (.A(_0858_),
    .B(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__or2_2 _3587_ (.A(_0255_),
    .B(_0258_),
    .X(_0949_));
 sky130_fd_sc_hd__a21o_1 _3588_ (.A1(net39),
    .A2(_0948_),
    .B1(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__o311a_1 _3589_ (.A1(_0938_),
    .A2(_0942_),
    .A3(_0945_),
    .B1(_0950_),
    .C1(\modetrans.mode[3] ),
    .X(_0951_));
 sky130_fd_sc_hd__or2_1 _3590_ (.A(\lvls.level[2] ),
    .B(\lvls.level[0] ),
    .X(_0952_));
 sky130_fd_sc_hd__o21a_2 _3591_ (.A1(\lvls.level[1] ),
    .A2(_0952_),
    .B1(\modetrans.mode[5] ),
    .X(_0953_));
 sky130_fd_sc_hd__a311o_1 _3592_ (.A1(_0211_),
    .A2(net39),
    .A3(_0948_),
    .B1(_0953_),
    .C1(_0214_),
    .X(_0954_));
 sky130_fd_sc_hd__o21a_1 _3593_ (.A1(_0951_),
    .A2(_0954_),
    .B1(_0935_),
    .X(net24));
 sky130_fd_sc_hd__nand2_2 _3594_ (.A(_0255_),
    .B(_0258_),
    .Y(_0955_));
 sky130_fd_sc_hd__and3_1 _3595_ (.A(_0909_),
    .B(_0913_),
    .C(_0936_),
    .X(_0956_));
 sky130_fd_sc_hd__or2_1 _3596_ (.A(_0955_),
    .B(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__o21ai_1 _3597_ (.A1(\highest_score.highest_score[4] ),
    .A2(_0906_),
    .B1(_0895_),
    .Y(_0958_));
 sky130_fd_sc_hd__and3b_1 _3598_ (.A_N(_0939_),
    .B(_0675_),
    .C(_0889_),
    .X(_0959_));
 sky130_fd_sc_hd__a22o_1 _3599_ (.A1(_0255_),
    .A2(_0958_),
    .B1(_0959_),
    .B2(_0258_),
    .X(_0960_));
 sky130_fd_sc_hd__a21oi_1 _3600_ (.A1(_0957_),
    .A2(_0960_),
    .B1(_0921_),
    .Y(_0961_));
 sky130_fd_sc_hd__or3_1 _3601_ (.A(_0840_),
    .B(_0859_),
    .C(_0946_),
    .X(_0962_));
 sky130_fd_sc_hd__o211a_1 _3602_ (.A1(_0211_),
    .A2(_0961_),
    .B1(_0962_),
    .C1(net39),
    .X(_0963_));
 sky130_fd_sc_hd__and2_1 _3603_ (.A(\disp_song.mi6.in[2] ),
    .B(_0926_),
    .X(_0964_));
 sky130_fd_sc_hd__a21o_1 _3604_ (.A1(\disp_song.mi6.in[3] ),
    .A2(_0964_),
    .B1(_0929_),
    .X(_0965_));
 sky130_fd_sc_hd__buf_6 _3605_ (.A(_2654_),
    .X(_0966_));
 sky130_fd_sc_hd__a221o_1 _3606_ (.A1(_0949_),
    .A2(_0961_),
    .B1(_0965_),
    .B2(_0966_),
    .C1(_0953_),
    .X(_0967_));
 sky130_fd_sc_hd__o21a_1 _3607_ (.A1(_0963_),
    .A2(_0967_),
    .B1(_0935_),
    .X(net25));
 sky130_fd_sc_hd__a211o_1 _3608_ (.A1(_0849_),
    .A2(_0855_),
    .B1(_0856_),
    .C1(_0861_),
    .X(_0968_));
 sky130_fd_sc_hd__or3_1 _3609_ (.A(_0617_),
    .B(_0609_),
    .C(_0614_),
    .X(_0969_));
 sky130_fd_sc_hd__and2b_1 _3610_ (.A_N(_0914_),
    .B(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__o21a_1 _3611_ (.A1(_0936_),
    .A2(_0970_),
    .B1(_0919_),
    .X(_0971_));
 sky130_fd_sc_hd__o21ai_1 _3612_ (.A1(_0916_),
    .A2(_0971_),
    .B1(_0261_),
    .Y(_0972_));
 sky130_fd_sc_hd__or2_1 _3613_ (.A(_0887_),
    .B(_0939_),
    .X(_0973_));
 sky130_fd_sc_hd__a21o_1 _3614_ (.A1(_0894_),
    .A2(_0973_),
    .B1(_0896_),
    .X(_0974_));
 sky130_fd_sc_hd__or2_1 _3615_ (.A(\highest_score.highest_score[4] ),
    .B(_0902_),
    .X(_0975_));
 sky130_fd_sc_hd__a21o_1 _3616_ (.A1(_0907_),
    .A2(_0975_),
    .B1(_0258_),
    .X(_0976_));
 sky130_fd_sc_hd__a31o_1 _3617_ (.A1(_0972_),
    .A2(_0974_),
    .A3(_0976_),
    .B1(_0921_),
    .X(_0977_));
 sky130_fd_sc_hd__nand2_1 _3618_ (.A(_0879_),
    .B(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__nor2_1 _3619_ (.A(_0259_),
    .B(_0977_),
    .Y(_0979_));
 sky130_fd_sc_hd__a31o_1 _3620_ (.A1(net39),
    .A2(_0968_),
    .A3(_0978_),
    .B1(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__o31a_1 _3621_ (.A1(_0931_),
    .A2(_0953_),
    .A3(_0980_),
    .B1(_0935_),
    .X(net26));
 sky130_fd_sc_hd__o21a_1 _3622_ (.A1(_0956_),
    .A2(_0971_),
    .B1(_0261_),
    .X(_0981_));
 sky130_fd_sc_hd__o2111a_1 _3623_ (.A1(\highest_score.highest_score[4] ),
    .A2(_0906_),
    .B1(_0975_),
    .C1(_0255_),
    .D1(_0904_),
    .X(_0982_));
 sky130_fd_sc_hd__nor2_1 _3624_ (.A(_0887_),
    .B(_0939_),
    .Y(_0983_));
 sky130_fd_sc_hd__or3_1 _3625_ (.A(_0893_),
    .B(_0959_),
    .C(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__a2bb2o_1 _3626_ (.A1_N(_0258_),
    .A2_N(_0982_),
    .B1(_0984_),
    .B2(_0941_),
    .X(_0985_));
 sky130_fd_sc_hd__o211a_1 _3627_ (.A1(_0849_),
    .A2(_0850_),
    .B1(_0855_),
    .C1(net39),
    .X(_0986_));
 sky130_fd_sc_hd__o221a_1 _3628_ (.A1(_0981_),
    .A2(_0985_),
    .B1(_0986_),
    .B2(_0949_),
    .C1(\modetrans.mode[3] ),
    .X(_0987_));
 sky130_fd_sc_hd__or2b_1 _3629_ (.A(_0928_),
    .B_N(_0965_),
    .X(_0988_));
 sky130_fd_sc_hd__a22o_1 _3630_ (.A1(_0214_),
    .A2(_0988_),
    .B1(_0986_),
    .B2(_0211_),
    .X(_0989_));
 sky130_fd_sc_hd__o31a_1 _3631_ (.A1(_0953_),
    .A2(_0987_),
    .A3(_0989_),
    .B1(_0935_),
    .X(net27));
 sky130_fd_sc_hd__nor2_1 _3632_ (.A(_0840_),
    .B(_0855_),
    .Y(_0990_));
 sky130_fd_sc_hd__o21ai_1 _3633_ (.A1(_0835_),
    .A2(_0990_),
    .B1(_0848_),
    .Y(_0991_));
 sky130_fd_sc_hd__o21bai_1 _3634_ (.A1(_0667_),
    .A2(_0969_),
    .B1_N(_0914_),
    .Y(_0992_));
 sky130_fd_sc_hd__a211o_1 _3635_ (.A1(_0919_),
    .A2(_0970_),
    .B1(_0992_),
    .C1(_0915_),
    .X(_0993_));
 sky130_fd_sc_hd__a31o_1 _3636_ (.A1(_0608_),
    .A2(_0675_),
    .A3(_0671_),
    .B1(_0886_),
    .X(_0994_));
 sky130_fd_sc_hd__o31a_1 _3637_ (.A1(_0891_),
    .A2(_0893_),
    .A3(_0994_),
    .B1(_0941_),
    .X(_0995_));
 sky130_fd_sc_hd__and3b_1 _3638_ (.A_N(_0943_),
    .B(_0255_),
    .C(_0901_),
    .X(_0996_));
 sky130_fd_sc_hd__a21oi_1 _3639_ (.A1(_0904_),
    .A2(_0996_),
    .B1(_0258_),
    .Y(_0997_));
 sky130_fd_sc_hd__a211o_1 _3640_ (.A1(_0261_),
    .A2(_0993_),
    .B1(_0995_),
    .C1(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__nand2_1 _3641_ (.A(\modetrans.mode[3] ),
    .B(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__inv_2 _3642_ (.A(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__o221a_1 _3643_ (.A1(_0856_),
    .A2(_0991_),
    .B1(_1000_),
    .B2(_0211_),
    .C1(net39),
    .X(_1001_));
 sky130_fd_sc_hd__a22o_1 _3644_ (.A1(_0214_),
    .A2(_0928_),
    .B1(_1000_),
    .B2(_0949_),
    .X(_1002_));
 sky130_fd_sc_hd__o21a_1 _3645_ (.A1(_1001_),
    .A2(_1002_),
    .B1(_0935_),
    .X(net28));
 sky130_fd_sc_hd__nor2_1 _3646_ (.A(_0840_),
    .B(_0859_),
    .Y(_1003_));
 sky130_fd_sc_hd__o21ai_1 _3647_ (.A1(_0892_),
    .A2(_0994_),
    .B1(_0941_),
    .Y(_1004_));
 sky130_fd_sc_hd__o21ai_1 _3648_ (.A1(_0918_),
    .A2(_0992_),
    .B1(_0261_),
    .Y(_1005_));
 sky130_fd_sc_hd__a21o_1 _3649_ (.A1(_0906_),
    .A2(_0996_),
    .B1(_0258_),
    .X(_1006_));
 sky130_fd_sc_hd__a31o_1 _3650_ (.A1(_1004_),
    .A2(_1005_),
    .A3(_1006_),
    .B1(_0921_),
    .X(_1007_));
 sky130_fd_sc_hd__inv_2 _3651_ (.A(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__o221a_1 _3652_ (.A1(_1003_),
    .A2(_0991_),
    .B1(_1008_),
    .B2(_0211_),
    .C1(net38),
    .X(_1009_));
 sky130_fd_sc_hd__nor2_1 _3653_ (.A(_0259_),
    .B(_1007_),
    .Y(_1010_));
 sky130_fd_sc_hd__o41a_2 _3654_ (.A1(_0930_),
    .A2(_0953_),
    .A3(_1009_),
    .A4(_1010_),
    .B1(_0935_),
    .X(net29));
 sky130_fd_sc_hd__inv_2 _3655_ (.A(_0789_),
    .Y(_1011_));
 sky130_fd_sc_hd__inv_2 _3656_ (.A(_0806_),
    .Y(_1012_));
 sky130_fd_sc_hd__and2_1 _3657_ (.A(_0661_),
    .B(_0665_),
    .X(_1013_));
 sky130_fd_sc_hd__or2b_1 _3658_ (.A(_0662_),
    .B_N(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__nand2_1 _3659_ (.A(_0788_),
    .B(_1014_),
    .Y(_1015_));
 sky130_fd_sc_hd__or2_1 _3660_ (.A(_0787_),
    .B(_1013_),
    .X(_1016_));
 sky130_fd_sc_hd__and3_1 _3661_ (.A(_0786_),
    .B(_0806_),
    .C(_1016_),
    .X(_1017_));
 sky130_fd_sc_hd__a22o_1 _3662_ (.A1(_1012_),
    .A2(_0807_),
    .B1(_1015_),
    .B2(_1017_),
    .X(_1018_));
 sky130_fd_sc_hd__and4bb_1 _3663_ (.A_N(_0775_),
    .B_N(_1018_),
    .C(_0776_),
    .D(net43),
    .X(_1019_));
 sky130_fd_sc_hd__or3b_1 _3664_ (.A(_0806_),
    .B(_1015_),
    .C_N(_1016_),
    .X(_1020_));
 sky130_fd_sc_hd__a41o_1 _3665_ (.A1(_0786_),
    .A2(_1011_),
    .A3(_1019_),
    .A4(_1020_),
    .B1(_0830_),
    .X(_1021_));
 sky130_fd_sc_hd__o21ai_2 _3666_ (.A1(_0834_),
    .A2(_1015_),
    .B1(_0830_),
    .Y(_1022_));
 sky130_fd_sc_hd__o311a_1 _3667_ (.A1(_0762_),
    .A2(_0824_),
    .A3(_0825_),
    .B1(_0826_),
    .C1(_0786_),
    .X(_1023_));
 sky130_fd_sc_hd__o2bb2a_2 _3668_ (.A1_N(_0830_),
    .A2_N(_0834_),
    .B1(_1019_),
    .B2(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__and3_1 _3669_ (.A(_1021_),
    .B(_1022_),
    .C(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__a21oi_1 _3670_ (.A1(_1021_),
    .A2(_1022_),
    .B1(_1024_),
    .Y(_1026_));
 sky130_fd_sc_hd__or4_1 _3671_ (.A(_0775_),
    .B(_0831_),
    .C(_0790_),
    .D(_0844_),
    .X(_1027_));
 sky130_fd_sc_hd__mux2_2 _3672_ (.A0(_0834_),
    .A1(_1027_),
    .S(net42),
    .X(_1028_));
 sky130_fd_sc_hd__a21oi_2 _3673_ (.A1(net42),
    .A2(_0806_),
    .B1(_1016_),
    .Y(_1029_));
 sky130_fd_sc_hd__o21a_1 _3674_ (.A1(_0807_),
    .A2(_1017_),
    .B1(net42),
    .X(_1030_));
 sky130_fd_sc_hd__or3_4 _3675_ (.A(_1028_),
    .B(_1029_),
    .C(_1030_),
    .X(_1031_));
 sky130_fd_sc_hd__mux2_2 _3676_ (.A0(_1025_),
    .A1(_1026_),
    .S(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__a21boi_2 _3677_ (.A1(_1021_),
    .A2(_1022_),
    .B1_N(_1024_),
    .Y(_1033_));
 sky130_fd_sc_hd__or2_2 _3678_ (.A(_1012_),
    .B(_1028_),
    .X(_1034_));
 sky130_fd_sc_hd__nor3_2 _3679_ (.A(_1028_),
    .B(_1029_),
    .C(_1030_),
    .Y(_1035_));
 sky130_fd_sc_hd__mux2_1 _3680_ (.A0(_1025_),
    .A1(_1033_),
    .S(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__a311oi_4 _3681_ (.A1(_1031_),
    .A2(_1033_),
    .A3(_1034_),
    .B1(_1036_),
    .C1(_1032_),
    .Y(_1037_));
 sky130_fd_sc_hd__and3_1 _3682_ (.A(_1025_),
    .B(_1031_),
    .C(_1034_),
    .X(_1038_));
 sky130_fd_sc_hd__a21o_1 _3683_ (.A1(_1035_),
    .A2(_1033_),
    .B1(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__and3_1 _3684_ (.A(_0625_),
    .B(_0649_),
    .C(net44),
    .X(_1040_));
 sky130_fd_sc_hd__o21ai_1 _3685_ (.A1(_0625_),
    .A2(_0880_),
    .B1(net44),
    .Y(_1041_));
 sky130_fd_sc_hd__a21oi_1 _3686_ (.A1(_0642_),
    .A2(_1040_),
    .B1(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__or2b_1 _3687_ (.A(_0642_),
    .B_N(_1040_),
    .X(_1043_));
 sky130_fd_sc_hd__nand2_1 _3688_ (.A(_0625_),
    .B(net44),
    .Y(_1044_));
 sky130_fd_sc_hd__or3b_1 _3689_ (.A(_0649_),
    .B(_1044_),
    .C_N(_0642_),
    .X(_1045_));
 sky130_fd_sc_hd__nand2_1 _3690_ (.A(_1043_),
    .B(_1045_),
    .Y(_1046_));
 sky130_fd_sc_hd__or2_1 _3691_ (.A(_0649_),
    .B(_1044_),
    .X(_1047_));
 sky130_fd_sc_hd__o31ai_1 _3692_ (.A1(_0642_),
    .A2(_0638_),
    .A3(_1047_),
    .B1(_1042_),
    .Y(_1048_));
 sky130_fd_sc_hd__or2_1 _3693_ (.A(_1046_),
    .B(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__o211a_1 _3694_ (.A1(_0638_),
    .A2(_1043_),
    .B1(_1045_),
    .C1(_1049_),
    .X(_1050_));
 sky130_fd_sc_hd__a21o_1 _3695_ (.A1(_1042_),
    .A2(_1050_),
    .B1(_0896_),
    .X(_1051_));
 sky130_fd_sc_hd__inv_2 _3696_ (.A(\highest_score.highest_score[1] ),
    .Y(_1052_));
 sky130_fd_sc_hd__inv_2 _3697_ (.A(\highest_score.highest_score[2] ),
    .Y(_1053_));
 sky130_fd_sc_hd__or2_1 _3698_ (.A(\highest_score.highest_score[3] ),
    .B(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__or3b_1 _3699_ (.A(\highest_score.highest_score[2] ),
    .B(\highest_score.highest_score[1] ),
    .C_N(\highest_score.highest_score[3] ),
    .X(_1055_));
 sky130_fd_sc_hd__o21a_1 _3700_ (.A1(_1052_),
    .A2(_1054_),
    .B1(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__inv_2 _3701_ (.A(\highest_score.highest_score[0] ),
    .Y(_1057_));
 sky130_fd_sc_hd__a31o_1 _3702_ (.A1(_1053_),
    .A2(_1052_),
    .A3(_1057_),
    .B1(\highest_score.highest_score[3] ),
    .X(_1058_));
 sky130_fd_sc_hd__nand2_1 _3703_ (.A(_1055_),
    .B(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__and2_1 _3704_ (.A(_0255_),
    .B(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__or3_1 _3705_ (.A(\highest_score.highest_score[3] ),
    .B(\highest_score.highest_score[2] ),
    .C(_1052_),
    .X(_1061_));
 sky130_fd_sc_hd__o311a_1 _3706_ (.A1(\highest_score.highest_score[1] ),
    .A2(_1057_),
    .A3(_1054_),
    .B1(_1060_),
    .C1(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__a21o_1 _3707_ (.A1(_1056_),
    .A2(_1062_),
    .B1(_0258_),
    .X(_1063_));
 sky130_fd_sc_hd__nand2_1 _3708_ (.A(_0651_),
    .B(_0652_),
    .Y(_1064_));
 sky130_fd_sc_hd__or3b_1 _3709_ (.A(_0633_),
    .B(_0912_),
    .C_N(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__or2_1 _3710_ (.A(_0629_),
    .B(_1065_),
    .X(_1066_));
 sky130_fd_sc_hd__or3_1 _3711_ (.A(_0633_),
    .B(_1064_),
    .C(_0912_),
    .X(_1067_));
 sky130_fd_sc_hd__or2_1 _3712_ (.A(_0641_),
    .B(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__o21ai_1 _3713_ (.A1(_0636_),
    .A2(_1066_),
    .B1(_1068_),
    .Y(_1069_));
 sky130_fd_sc_hd__or2_1 _3714_ (.A(_0629_),
    .B(_0636_),
    .X(_1070_));
 sky130_fd_sc_hd__o211a_1 _3715_ (.A1(_1067_),
    .A2(_1070_),
    .B1(_1066_),
    .C1(_1068_),
    .X(_1071_));
 sky130_fd_sc_hd__o21ai_1 _3716_ (.A1(_1069_),
    .A2(_1071_),
    .B1(_0261_),
    .Y(_1072_));
 sky130_fd_sc_hd__a31o_1 _3717_ (.A1(_1051_),
    .A2(_1063_),
    .A3(_1072_),
    .B1(_0921_),
    .X(_1073_));
 sky130_fd_sc_hd__nand2_1 _3718_ (.A(_0879_),
    .B(_1073_),
    .Y(_1074_));
 sky130_fd_sc_hd__o311a_1 _3719_ (.A1(_1032_),
    .A2(_1037_),
    .A3(_1039_),
    .B1(_1074_),
    .C1(net38),
    .X(_1075_));
 sky130_fd_sc_hd__o21a_1 _3720_ (.A1(\lvls.level[2] ),
    .A2(\lvls.level[1] ),
    .B1(\modetrans.mode[5] ),
    .X(_1076_));
 sky130_fd_sc_hd__clkbuf_4 _3721_ (.A(\disp_song.mi6.in[0] ),
    .X(_1077_));
 sky130_fd_sc_hd__nand2_1 _3722_ (.A(\disp_song.mi6.in[3] ),
    .B(_0926_),
    .Y(_1078_));
 sky130_fd_sc_hd__or2_1 _3723_ (.A(\disp_song.mi6.in[3] ),
    .B(_0926_),
    .X(_1079_));
 sky130_fd_sc_hd__and2_1 _3724_ (.A(_1078_),
    .B(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__inv_2 _3725_ (.A(\disp_song.mi6.in[2] ),
    .Y(_1081_));
 sky130_fd_sc_hd__nand2_2 _3726_ (.A(\disp_song.mi6.in[3] ),
    .B(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__nor2_1 _3727_ (.A(_1077_),
    .B(_1082_),
    .Y(_1083_));
 sky130_fd_sc_hd__nor2_1 _3728_ (.A(_1081_),
    .B(_1080_),
    .Y(_1084_));
 sky130_fd_sc_hd__o221a_1 _3729_ (.A1(_1077_),
    .A2(_1080_),
    .B1(_1083_),
    .B2(_1084_),
    .C1(_0925_),
    .X(_1085_));
 sky130_fd_sc_hd__nor2_1 _3730_ (.A(\disp_song.mi6.in[2] ),
    .B(_1077_),
    .Y(_1086_));
 sky130_fd_sc_hd__a2111o_1 _3731_ (.A1(_1077_),
    .A2(_1084_),
    .B1(_1086_),
    .C1(_0925_),
    .D1(_1080_),
    .X(_1087_));
 sky130_fd_sc_hd__or3b_1 _3732_ (.A(_0352_),
    .B(_1085_),
    .C_N(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__o21ai_1 _3733_ (.A1(_0259_),
    .A2(_1073_),
    .B1(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__o31a_2 _3734_ (.A1(_1075_),
    .A2(_1076_),
    .A3(_1089_),
    .B1(_0935_),
    .X(net16));
 sky130_fd_sc_hd__inv_2 _3735_ (.A(net38),
    .Y(_1090_));
 sky130_fd_sc_hd__and3_1 _3736_ (.A(_0806_),
    .B(_1025_),
    .C(_1035_),
    .X(_1091_));
 sky130_fd_sc_hd__and2b_1 _3737_ (.A_N(_0912_),
    .B(_0636_),
    .X(_1092_));
 sky130_fd_sc_hd__nand2_1 _3738_ (.A(_0629_),
    .B(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__a21o_1 _3739_ (.A1(_1070_),
    .A2(_1093_),
    .B1(_1065_),
    .X(_1094_));
 sky130_fd_sc_hd__nor2_1 _3740_ (.A(_0642_),
    .B(_0638_),
    .Y(_1095_));
 sky130_fd_sc_hd__and3_1 _3741_ (.A(_0642_),
    .B(_0638_),
    .C(net44),
    .X(_1096_));
 sky130_fd_sc_hd__o21ai_1 _3742_ (.A1(_1095_),
    .A2(_1096_),
    .B1(_1040_),
    .Y(_1097_));
 sky130_fd_sc_hd__a21o_1 _3743_ (.A1(\highest_score.highest_score[1] ),
    .A2(\highest_score.highest_score[0] ),
    .B1(_1054_),
    .X(_1098_));
 sky130_fd_sc_hd__o21ai_1 _3744_ (.A1(\highest_score.highest_score[1] ),
    .A2(\highest_score.highest_score[0] ),
    .B1(_0255_),
    .Y(_1099_));
 sky130_fd_sc_hd__o21a_1 _3745_ (.A1(_1098_),
    .A2(_1099_),
    .B1(_0895_),
    .X(_1100_));
 sky130_fd_sc_hd__a221o_1 _3746_ (.A1(_0261_),
    .A2(_1094_),
    .B1(_1097_),
    .B2(_0941_),
    .C1(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__a21oi_1 _3747_ (.A1(\modetrans.mode[3] ),
    .A2(_1101_),
    .B1(_0211_),
    .Y(_1102_));
 sky130_fd_sc_hd__nor4_1 _3748_ (.A(_1090_),
    .B(_1038_),
    .C(_1091_),
    .D(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__nor2_1 _3749_ (.A(_1077_),
    .B(_0926_),
    .Y(_1104_));
 sky130_fd_sc_hd__nand2_1 _3750_ (.A(_1077_),
    .B(_0926_),
    .Y(_1105_));
 sky130_fd_sc_hd__or3b_1 _3751_ (.A(_1104_),
    .B(_1082_),
    .C_N(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__or2_1 _3752_ (.A(_1077_),
    .B(_0926_),
    .X(_1107_));
 sky130_fd_sc_hd__or3_1 _3753_ (.A(\disp_song.mi6.in[3] ),
    .B(\disp_song.mi6.in[2] ),
    .C(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__a21bo_1 _3754_ (.A1(_1106_),
    .A2(_1108_),
    .B1_N(_0925_),
    .X(_1109_));
 sky130_fd_sc_hd__a21oi_1 _3755_ (.A1(_1105_),
    .A2(_1107_),
    .B1(\disp_song.mi6.in[3] ),
    .Y(_1110_));
 sky130_fd_sc_hd__a2111o_1 _3756_ (.A1(\disp_song.mi6.in[3] ),
    .A2(_1105_),
    .B1(_1110_),
    .C1(_1081_),
    .D1(_0925_),
    .X(_1111_));
 sky130_fd_sc_hd__a31o_1 _3757_ (.A1(_0966_),
    .A2(_1109_),
    .A3(_1111_),
    .B1(_0953_),
    .X(_1112_));
 sky130_fd_sc_hd__a31o_1 _3758_ (.A1(\modetrans.mode[3] ),
    .A2(_0949_),
    .A3(_1101_),
    .B1(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__o21a_1 _3759_ (.A1(_1103_),
    .A2(_1113_),
    .B1(_0935_),
    .X(net17));
 sky130_fd_sc_hd__inv_2 _3760_ (.A(_1077_),
    .Y(_1114_));
 sky130_fd_sc_hd__nor2_1 _3761_ (.A(_0925_),
    .B(_0964_),
    .Y(_1115_));
 sky130_fd_sc_hd__nand2_1 _3762_ (.A(\disp_song.mi6.in[2] ),
    .B(_0926_),
    .Y(_1116_));
 sky130_fd_sc_hd__nor2_1 _3763_ (.A(\disp_song.mi6.in[3] ),
    .B(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__a32o_1 _3764_ (.A1(_1079_),
    .A2(_1082_),
    .A3(_1115_),
    .B1(_1117_),
    .B2(_0925_),
    .X(_1118_));
 sky130_fd_sc_hd__a21oi_1 _3765_ (.A1(_1114_),
    .A2(_1118_),
    .B1(_0352_),
    .Y(_1119_));
 sky130_fd_sc_hd__and3_1 _3766_ (.A(_0806_),
    .B(_1035_),
    .C(_1033_),
    .X(_1120_));
 sky130_fd_sc_hd__nor2_1 _3767_ (.A(_1090_),
    .B(_1120_),
    .Y(_1121_));
 sky130_fd_sc_hd__or2_1 _3768_ (.A(_1067_),
    .B(_1093_),
    .X(_1122_));
 sky130_fd_sc_hd__or2_1 _3769_ (.A(\highest_score.highest_score[0] ),
    .B(_1061_),
    .X(_1123_));
 sky130_fd_sc_hd__a21bo_1 _3770_ (.A1(_0895_),
    .A2(_1123_),
    .B1_N(_0255_),
    .X(_1124_));
 sky130_fd_sc_hd__and2b_1 _3771_ (.A_N(_1047_),
    .B(_1096_),
    .X(_1125_));
 sky130_fd_sc_hd__nand2_1 _3772_ (.A(_0258_),
    .B(_1125_),
    .Y(_1126_));
 sky130_fd_sc_hd__a22o_1 _3773_ (.A1(_0261_),
    .A2(_1122_),
    .B1(_1124_),
    .B2(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__o211a_1 _3774_ (.A1(_0949_),
    .A2(_1121_),
    .B1(_1127_),
    .C1(\modetrans.mode[3] ),
    .X(_1128_));
 sky130_fd_sc_hd__a22o_1 _3775_ (.A1(\modetrans.mode[5] ),
    .A2(_0952_),
    .B1(_1121_),
    .B2(_0211_),
    .X(_1129_));
 sky130_fd_sc_hd__o31a_2 _3776_ (.A1(_1119_),
    .A2(_1128_),
    .A3(_1129_),
    .B1(_0935_),
    .X(net18));
 sky130_fd_sc_hd__and2b_1 _3777_ (.A_N(_1034_),
    .B(_1032_),
    .X(_1130_));
 sky130_fd_sc_hd__a21oi_1 _3778_ (.A1(_0633_),
    .A2(_0630_),
    .B1(_0912_),
    .Y(_1131_));
 sky130_fd_sc_hd__o21a_1 _3779_ (.A1(_0633_),
    .A2(_0653_),
    .B1(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__o21ai_1 _3780_ (.A1(_1092_),
    .A2(_1132_),
    .B1(_1071_),
    .Y(_1133_));
 sky130_fd_sc_hd__and2b_1 _3781_ (.A_N(_1069_),
    .B(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__or2_1 _3782_ (.A(\highest_score.highest_score[0] ),
    .B(_1056_),
    .X(_1135_));
 sky130_fd_sc_hd__a21o_1 _3783_ (.A1(_1062_),
    .A2(_1135_),
    .B1(_0258_),
    .X(_1136_));
 sky130_fd_sc_hd__or3b_1 _3784_ (.A(_0639_),
    .B(_1042_),
    .C_N(net44),
    .X(_1137_));
 sky130_fd_sc_hd__a21o_1 _3785_ (.A1(_1050_),
    .A2(_1137_),
    .B1(_0896_),
    .X(_1138_));
 sky130_fd_sc_hd__o211a_1 _3786_ (.A1(_0955_),
    .A2(_1134_),
    .B1(_1136_),
    .C1(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__nor2_1 _3787_ (.A(_0921_),
    .B(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__or2_1 _3788_ (.A(_0210_),
    .B(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__o311a_1 _3789_ (.A1(_1037_),
    .A2(_1039_),
    .A3(_1130_),
    .B1(_1141_),
    .C1(net38),
    .X(_1142_));
 sky130_fd_sc_hd__o221a_1 _3790_ (.A1(\disp_song.mi6.in[3] ),
    .A2(_1116_),
    .B1(_1082_),
    .B2(_0926_),
    .C1(_1077_),
    .X(_1143_));
 sky130_fd_sc_hd__o31ai_1 _3791_ (.A1(_1077_),
    .A2(_0926_),
    .A3(_1082_),
    .B1(_0925_),
    .Y(_1144_));
 sky130_fd_sc_hd__o21bai_1 _3792_ (.A1(_1077_),
    .A2(_1078_),
    .B1_N(_1110_),
    .Y(_1145_));
 sky130_fd_sc_hd__o21ai_1 _3793_ (.A1(\disp_song.mi6.in[2] ),
    .A2(_0926_),
    .B1(_1082_),
    .Y(_1146_));
 sky130_fd_sc_hd__a221o_1 _3794_ (.A1(\disp_song.mi6.in[2] ),
    .A2(_1145_),
    .B1(_1146_),
    .B2(_1077_),
    .C1(_0925_),
    .X(_1147_));
 sky130_fd_sc_hd__o21ai_1 _3795_ (.A1(_1143_),
    .A2(_1144_),
    .B1(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__a221o_1 _3796_ (.A1(_0949_),
    .A2(_1140_),
    .B1(_1148_),
    .B2(_0966_),
    .C1(_1076_),
    .X(_1149_));
 sky130_fd_sc_hd__o21a_1 _3797_ (.A1(_1142_),
    .A2(_1149_),
    .B1(_0935_),
    .X(net19));
 sky130_fd_sc_hd__inv_2 _3798_ (.A(_1125_),
    .Y(_1150_));
 sky130_fd_sc_hd__a31o_1 _3799_ (.A1(_1049_),
    .A2(_1150_),
    .A3(_1137_),
    .B1(_0896_),
    .X(_1151_));
 sky130_fd_sc_hd__a31o_1 _3800_ (.A1(_1060_),
    .A2(_1123_),
    .A3(_1135_),
    .B1(_0258_),
    .X(_1152_));
 sky130_fd_sc_hd__a21o_1 _3801_ (.A1(_1122_),
    .A2(_1133_),
    .B1(_0955_),
    .X(_1153_));
 sky130_fd_sc_hd__a31o_1 _3802_ (.A1(_1151_),
    .A2(_1152_),
    .A3(_1153_),
    .B1(_0921_),
    .X(_1154_));
 sky130_fd_sc_hd__nand2_1 _3803_ (.A(_0879_),
    .B(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__o311a_1 _3804_ (.A1(_1037_),
    .A2(_1120_),
    .A3(_1130_),
    .B1(_1155_),
    .C1(net38),
    .X(_1156_));
 sky130_fd_sc_hd__nor2_1 _3805_ (.A(_0259_),
    .B(_1154_),
    .Y(_1157_));
 sky130_fd_sc_hd__o21ai_1 _3806_ (.A1(_0926_),
    .A2(_1082_),
    .B1(_0925_),
    .Y(_1158_));
 sky130_fd_sc_hd__o21ai_1 _3807_ (.A1(_0925_),
    .A2(_1084_),
    .B1(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__a32o_1 _3808_ (.A1(_0966_),
    .A2(_1114_),
    .A3(_1159_),
    .B1(\modetrans.mode[5] ),
    .B2(\lvls.level[1] ),
    .X(_1160_));
 sky130_fd_sc_hd__o31a_2 _3809_ (.A1(_1156_),
    .A2(_1157_),
    .A3(_1160_),
    .B1(_0935_),
    .X(net20));
 sky130_fd_sc_hd__and2_1 _3810_ (.A(_1025_),
    .B(_1031_),
    .X(_1161_));
 sky130_fd_sc_hd__a21o_1 _3811_ (.A1(_1031_),
    .A2(_1026_),
    .B1(_1091_),
    .X(_1162_));
 sky130_fd_sc_hd__nand2_1 _3812_ (.A(_1071_),
    .B(_1132_),
    .Y(_1163_));
 sky130_fd_sc_hd__or3b_1 _3813_ (.A(_0633_),
    .B(_0653_),
    .C_N(_0636_),
    .X(_1164_));
 sky130_fd_sc_hd__a41o_1 _3814_ (.A1(_1066_),
    .A2(_1131_),
    .A3(_1163_),
    .A4(_1164_),
    .B1(_0955_),
    .X(_1165_));
 sky130_fd_sc_hd__a31o_1 _3815_ (.A1(_0642_),
    .A2(_0638_),
    .A3(_1040_),
    .B1(_1041_),
    .X(_1166_));
 sky130_fd_sc_hd__inv_2 _3816_ (.A(_1166_),
    .Y(_1167_));
 sky130_fd_sc_hd__a31o_1 _3817_ (.A1(_1043_),
    .A2(_1049_),
    .A3(_1167_),
    .B1(_0896_),
    .X(_1168_));
 sky130_fd_sc_hd__and2_1 _3818_ (.A(_0255_),
    .B(_1055_),
    .X(_1169_));
 sky130_fd_sc_hd__a31o_1 _3819_ (.A1(_1059_),
    .A2(_1098_),
    .A3(_1169_),
    .B1(_0258_),
    .X(_1170_));
 sky130_fd_sc_hd__a31o_1 _3820_ (.A1(_1165_),
    .A2(_1168_),
    .A3(_1170_),
    .B1(_0921_),
    .X(_1171_));
 sky130_fd_sc_hd__nand2_1 _3821_ (.A(_0879_),
    .B(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__o311a_1 _3822_ (.A1(_1161_),
    .A2(_1037_),
    .A3(_1162_),
    .B1(_1172_),
    .C1(net38),
    .X(_1173_));
 sky130_fd_sc_hd__o221a_1 _3823_ (.A1(\disp_song.mi6.in[3] ),
    .A2(_1116_),
    .B1(_1080_),
    .B2(_1114_),
    .C1(_0925_),
    .X(_1174_));
 sky130_fd_sc_hd__and3b_1 _3824_ (.A_N(_1086_),
    .B(_0927_),
    .C(_1116_),
    .X(_1175_));
 sky130_fd_sc_hd__a211o_1 _3825_ (.A1(\disp_song.mi6.in[2] ),
    .A2(_1105_),
    .B1(_1104_),
    .C1(\disp_song.mi6.in[3] ),
    .X(_1176_));
 sky130_fd_sc_hd__or3b_1 _3826_ (.A(_0925_),
    .B(_1175_),
    .C_N(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__or2b_1 _3827_ (.A(_1174_),
    .B_N(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__a2bb2o_1 _3828_ (.A1_N(_0259_),
    .A2_N(_1171_),
    .B1(_1178_),
    .B2(_0214_),
    .X(_1179_));
 sky130_fd_sc_hd__o21a_1 _3829_ (.A1(_1173_),
    .A2(_1179_),
    .B1(_0935_),
    .X(net21));
 sky130_fd_sc_hd__o21ai_1 _3830_ (.A1(_1046_),
    .A2(_1166_),
    .B1(_0941_),
    .Y(_1180_));
 sky130_fd_sc_hd__a41o_1 _3831_ (.A1(_1068_),
    .A2(_1066_),
    .A3(_1131_),
    .A4(_1164_),
    .B1(_0955_),
    .X(_1181_));
 sky130_fd_sc_hd__a31o_1 _3832_ (.A1(_1061_),
    .A2(_1098_),
    .A3(_1169_),
    .B1(_0258_),
    .X(_1182_));
 sky130_fd_sc_hd__a31o_1 _3833_ (.A1(_1180_),
    .A2(_1181_),
    .A3(_1182_),
    .B1(_0921_),
    .X(_1183_));
 sky130_fd_sc_hd__nand2_1 _3834_ (.A(_0879_),
    .B(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__o211a_1 _3835_ (.A1(_1036_),
    .A2(_1162_),
    .B1(_1184_),
    .C1(net38),
    .X(_1185_));
 sky130_fd_sc_hd__o2bb2a_1 _3836_ (.A1_N(_1077_),
    .A2_N(_1117_),
    .B1(_1080_),
    .B2(\disp_song.mi6.in[2] ),
    .X(_1186_));
 sky130_fd_sc_hd__or3b_1 _3837_ (.A(_1080_),
    .B(_1086_),
    .C_N(_0925_),
    .X(_1187_));
 sky130_fd_sc_hd__o211a_1 _3838_ (.A1(_0925_),
    .A2(_1186_),
    .B1(_1187_),
    .C1(_0966_),
    .X(_1188_));
 sky130_fd_sc_hd__nor2_1 _3839_ (.A(_0259_),
    .B(_1183_),
    .Y(_1189_));
 sky130_fd_sc_hd__o41a_2 _3840_ (.A1(_1076_),
    .A2(_1185_),
    .A3(_1188_),
    .A4(_1189_),
    .B1(_0935_),
    .X(net22));
 sky130_fd_sc_hd__o21a_1 _3841_ (.A1(\game.hit_1 ),
    .A2(\game.hit_2 ),
    .B1(_0210_),
    .X(_1190_));
 sky130_fd_sc_hd__a221o_2 _3842_ (.A1(_0966_),
    .A2(\disp_song.toggle_green ),
    .B1(_0262_),
    .B2(\modetrans.mode[3] ),
    .C1(_1190_),
    .X(_1191_));
 sky130_fd_sc_hd__and2_1 _3843_ (.A(_0933_),
    .B(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__clkbuf_1 _3844_ (.A(_1192_),
    .X(net14));
 sky130_fd_sc_hd__o21a_1 _3845_ (.A1(\game.missed_1 ),
    .A2(\game.missed_2 ),
    .B1(_0211_),
    .X(_1193_));
 sky130_fd_sc_hd__a22o_1 _3846_ (.A1(\modetrans.mode[3] ),
    .A2(_0255_),
    .B1(\disp_song.toggle_red ),
    .B2(_0214_),
    .X(_1194_));
 sky130_fd_sc_hd__o21a_1 _3847_ (.A1(_1193_),
    .A2(_1194_),
    .B1(_0933_),
    .X(net15));
 sky130_fd_sc_hd__a221o_2 _3848_ (.A1(_0966_),
    .A2(\disp_song.display_note1[0] ),
    .B1(_0211_),
    .B2(\game.out[7] ),
    .C1(_0208_),
    .X(_1195_));
 sky130_fd_sc_hd__and2_1 _3849_ (.A(_0933_),
    .B(_1195_),
    .X(_1196_));
 sky130_fd_sc_hd__clkbuf_1 _3850_ (.A(_1196_),
    .X(net7));
 sky130_fd_sc_hd__a221o_2 _3851_ (.A1(_0966_),
    .A2(\disp_song.display_note1[1] ),
    .B1(_0211_),
    .B2(\game.out[8] ),
    .C1(_0208_),
    .X(_1197_));
 sky130_fd_sc_hd__and2_1 _3852_ (.A(_0933_),
    .B(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__clkbuf_1 _3853_ (.A(_1198_),
    .X(net8));
 sky130_fd_sc_hd__a221o_2 _3854_ (.A1(_0966_),
    .A2(\disp_song.display_note1[2] ),
    .B1(_0211_),
    .B2(\game.out[9] ),
    .C1(_0208_),
    .X(_1199_));
 sky130_fd_sc_hd__and2_1 _3855_ (.A(_0933_),
    .B(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__clkbuf_1 _3856_ (.A(_1200_),
    .X(net9));
 sky130_fd_sc_hd__a221o_2 _3857_ (.A1(_0966_),
    .A2(\disp_song.display_note1[3] ),
    .B1(_0211_),
    .B2(\game.out[10] ),
    .C1(_0208_),
    .X(_1201_));
 sky130_fd_sc_hd__and2_1 _3858_ (.A(_0933_),
    .B(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__clkbuf_1 _3859_ (.A(_1202_),
    .X(net10));
 sky130_fd_sc_hd__a221o_2 _3860_ (.A1(_0966_),
    .A2(\disp_song.display_note1[4] ),
    .B1(_0211_),
    .B2(\game.out[11] ),
    .C1(_0208_),
    .X(_1203_));
 sky130_fd_sc_hd__and2_1 _3861_ (.A(_0933_),
    .B(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__clkbuf_1 _3862_ (.A(_1204_),
    .X(net11));
 sky130_fd_sc_hd__a221o_1 _3863_ (.A1(_0966_),
    .A2(\disp_song.display_note1[5] ),
    .B1(_0211_),
    .B2(\game.out[12] ),
    .C1(_0208_),
    .X(_1205_));
 sky130_fd_sc_hd__and2_1 _3864_ (.A(_0933_),
    .B(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__clkbuf_1 _3865_ (.A(_1206_),
    .X(net12));
 sky130_fd_sc_hd__a221o_2 _3866_ (.A1(_0966_),
    .A2(\disp_song.display_note1[6] ),
    .B1(_0211_),
    .B2(\game.out[13] ),
    .C1(_0208_),
    .X(_1207_));
 sky130_fd_sc_hd__and2_1 _3867_ (.A(_0933_),
    .B(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__clkbuf_1 _3868_ (.A(_1208_),
    .X(net13));
 sky130_fd_sc_hd__a221o_2 _3869_ (.A1(_0966_),
    .A2(\disp_song.display_note2[0] ),
    .B1(_0211_),
    .B2(\game.out[0] ),
    .C1(_0208_),
    .X(_1209_));
 sky130_fd_sc_hd__and2_1 _3870_ (.A(_0933_),
    .B(_1209_),
    .X(_1210_));
 sky130_fd_sc_hd__clkbuf_1 _3871_ (.A(_1210_),
    .X(net30));
 sky130_fd_sc_hd__a221o_1 _3872_ (.A1(_0966_),
    .A2(\disp_song.display_note2[1] ),
    .B1(_0211_),
    .B2(\game.out[1] ),
    .C1(_0208_),
    .X(_1211_));
 sky130_fd_sc_hd__and2_1 _3873_ (.A(_0933_),
    .B(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__clkbuf_1 _3874_ (.A(_1212_),
    .X(net31));
 sky130_fd_sc_hd__a221o_1 _3875_ (.A1(_0966_),
    .A2(\disp_song.display_note2[2] ),
    .B1(_0211_),
    .B2(\game.out[2] ),
    .C1(_0208_),
    .X(_1213_));
 sky130_fd_sc_hd__and2_1 _3876_ (.A(_0933_),
    .B(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__clkbuf_1 _3877_ (.A(_1214_),
    .X(net32));
 sky130_fd_sc_hd__a221o_2 _3878_ (.A1(_0966_),
    .A2(\disp_song.display_note2[3] ),
    .B1(_0211_),
    .B2(\game.out[3] ),
    .C1(_0208_),
    .X(_1215_));
 sky130_fd_sc_hd__and2_1 _3879_ (.A(_0933_),
    .B(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__clkbuf_1 _3880_ (.A(_1216_),
    .X(net33));
 sky130_fd_sc_hd__a221o_1 _3881_ (.A1(_0966_),
    .A2(\disp_song.display_note2[4] ),
    .B1(_0210_),
    .B2(\game.out[4] ),
    .C1(_0208_),
    .X(_1217_));
 sky130_fd_sc_hd__and2_1 _3882_ (.A(_0933_),
    .B(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__clkbuf_1 _3883_ (.A(_1218_),
    .X(net34));
 sky130_fd_sc_hd__a221o_2 _3884_ (.A1(_0966_),
    .A2(\disp_song.display_note2[5] ),
    .B1(_0210_),
    .B2(\game.out[5] ),
    .C1(_0208_),
    .X(_1219_));
 sky130_fd_sc_hd__and2_1 _3885_ (.A(_0933_),
    .B(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__clkbuf_1 _3886_ (.A(_1220_),
    .X(net35));
 sky130_fd_sc_hd__a221o_2 _3887_ (.A1(_0966_),
    .A2(\disp_song.display_note2[6] ),
    .B1(_0210_),
    .B2(\game.out[6] ),
    .C1(_0208_),
    .X(_1221_));
 sky130_fd_sc_hd__and2_1 _3888_ (.A(_0933_),
    .B(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__clkbuf_1 _3889_ (.A(_1222_),
    .X(net36));
 sky130_fd_sc_hd__and2_1 _3890_ (.A(_0933_),
    .B(net4),
    .X(_1223_));
 sky130_fd_sc_hd__clkbuf_1 _3891_ (.A(_1223_),
    .X(\modetrans.pushed_4 ));
 sky130_fd_sc_hd__and2_1 _3892_ (.A(_0933_),
    .B(net3),
    .X(_1224_));
 sky130_fd_sc_hd__clkbuf_1 _3893_ (.A(_1224_),
    .X(\modetrans.pushed_3 ));
 sky130_fd_sc_hd__and3b_1 _3894_ (.A_N(\game.scoring_button_2.check_hit.edge_1 ),
    .B(\game.scoring_button_2.check_hit.edge_2 ),
    .C(\game.scoring_button_2.hit ),
    .X(_1225_));
 sky130_fd_sc_hd__buf_6 _3895_ (.A(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__nor2_8 _3896_ (.A(_0208_),
    .B(_1226_),
    .Y(_1227_));
 sky130_fd_sc_hd__mux2_1 _3897_ (.A0(_1226_),
    .A1(_1227_),
    .S(\game.addhits.add1.b[0] ),
    .X(_1228_));
 sky130_fd_sc_hd__clkbuf_1 _3898_ (.A(_1228_),
    .X(\game.scoring_button_2.next_num_hits[0] ));
 sky130_fd_sc_hd__nor2_1 _3899_ (.A(\game.addhits.add1.b[2] ),
    .B(\game.scoring_button_2.acc[2] ),
    .Y(_1229_));
 sky130_fd_sc_hd__or2_1 _3900_ (.A(\game.addhits.add1.b[1] ),
    .B(\game.scoring_button_2.acc[1] ),
    .X(_1230_));
 sky130_fd_sc_hd__nand2_1 _3901_ (.A(\game.addhits.add1.b[1] ),
    .B(\game.scoring_button_2.acc[1] ),
    .Y(_1231_));
 sky130_fd_sc_hd__a21boi_1 _3902_ (.A1(\game.addhits.add1.b[0] ),
    .A2(_1230_),
    .B1_N(_1231_),
    .Y(_1232_));
 sky130_fd_sc_hd__nand2_1 _3903_ (.A(\game.addhits.add1.b[2] ),
    .B(\game.scoring_button_2.acc[2] ),
    .Y(_1233_));
 sky130_fd_sc_hd__o21ai_1 _3904_ (.A1(_1229_),
    .A2(_1232_),
    .B1(_1233_),
    .Y(_1234_));
 sky130_fd_sc_hd__nor2_1 _3905_ (.A(\game.addhits.add1.b[3] ),
    .B(_1234_),
    .Y(_1235_));
 sky130_fd_sc_hd__nand2_1 _3906_ (.A(_1231_),
    .B(_1230_),
    .Y(_1236_));
 sky130_fd_sc_hd__xor2_1 _3907_ (.A(\game.addhits.add1.b[0] ),
    .B(_1236_),
    .X(_1237_));
 sky130_fd_sc_hd__or2_1 _3908_ (.A(\game.addhits.add1.b[2] ),
    .B(\game.scoring_button_2.acc[2] ),
    .X(_1238_));
 sky130_fd_sc_hd__nand2_1 _3909_ (.A(_1233_),
    .B(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__xnor2_1 _3910_ (.A(_1232_),
    .B(_1239_),
    .Y(_1240_));
 sky130_fd_sc_hd__nand2_1 _3911_ (.A(_1237_),
    .B(_1240_),
    .Y(_1241_));
 sky130_fd_sc_hd__inv_2 _3912_ (.A(_1241_),
    .Y(_1242_));
 sky130_fd_sc_hd__nand2_1 _3913_ (.A(\game.addhits.add1.b[3] ),
    .B(_1234_),
    .Y(_1243_));
 sky130_fd_sc_hd__o21ai_2 _3914_ (.A1(_1235_),
    .A2(_1242_),
    .B1(_1243_),
    .Y(_1244_));
 sky130_fd_sc_hd__mux2_1 _3915_ (.A0(_1235_),
    .A1(_1244_),
    .S(_1237_),
    .X(_1245_));
 sky130_fd_sc_hd__a22o_1 _3916_ (.A1(\game.addhits.add1.b[1] ),
    .A2(_1227_),
    .B1(_1245_),
    .B2(_1226_),
    .X(\game.scoring_button_2.next_num_hits[1] ));
 sky130_fd_sc_hd__or2_1 _3917_ (.A(_1243_),
    .B(_1241_),
    .X(_1246_));
 sky130_fd_sc_hd__a21o_1 _3918_ (.A1(_1237_),
    .A2(_1244_),
    .B1(_1240_),
    .X(_1247_));
 sky130_fd_sc_hd__nand2_1 _3919_ (.A(_1246_),
    .B(_1247_),
    .Y(_1248_));
 sky130_fd_sc_hd__a22o_1 _3920_ (.A1(net167),
    .A2(_1227_),
    .B1(_1248_),
    .B2(_1226_),
    .X(\game.scoring_button_2.next_num_hits[2] ));
 sky130_fd_sc_hd__o21ai_1 _3921_ (.A1(_1235_),
    .A2(_1241_),
    .B1(_1243_),
    .Y(_1249_));
 sky130_fd_sc_hd__a32o_1 _3922_ (.A1(_1226_),
    .A2(_1246_),
    .A3(_1249_),
    .B1(_1227_),
    .B2(net178),
    .X(\game.scoring_button_2.next_num_hits[3] ));
 sky130_fd_sc_hd__or2_1 _3923_ (.A(\game.addhits.add2.b[0] ),
    .B(_1244_),
    .X(_1250_));
 sky130_fd_sc_hd__and2_1 _3924_ (.A(\game.addhits.add2.b[0] ),
    .B(_1244_),
    .X(_1251_));
 sky130_fd_sc_hd__inv_2 _3925_ (.A(_1251_),
    .Y(_1252_));
 sky130_fd_sc_hd__a32o_1 _3926_ (.A1(_1226_),
    .A2(_1250_),
    .A3(_1252_),
    .B1(_1227_),
    .B2(net188),
    .X(\game.scoring_button_2.next_num_hits[4] ));
 sky130_fd_sc_hd__o31a_2 _3927_ (.A1(\game.addhits.add2.b[2] ),
    .A2(\game.addhits.add2.b[1] ),
    .A3(_1251_),
    .B1(\game.addhits.add2.b[3] ),
    .X(_1253_));
 sky130_fd_sc_hd__xnor2_1 _3928_ (.A(\game.addhits.add2.b[1] ),
    .B(_1251_),
    .Y(_1254_));
 sky130_fd_sc_hd__xnor2_1 _3929_ (.A(_1253_),
    .B(_1254_),
    .Y(_1255_));
 sky130_fd_sc_hd__a22o_1 _3930_ (.A1(\game.addhits.add2.b[1] ),
    .A2(_1227_),
    .B1(_1255_),
    .B2(_1226_),
    .X(\game.scoring_button_2.next_num_hits[5] ));
 sky130_fd_sc_hd__inv_2 _3931_ (.A(\game.addhits.add2.b[2] ),
    .Y(_1256_));
 sky130_fd_sc_hd__inv_2 _3932_ (.A(\game.addhits.add2.b[1] ),
    .Y(_1257_));
 sky130_fd_sc_hd__or3_1 _3933_ (.A(_1256_),
    .B(_1257_),
    .C(_1252_),
    .X(_1258_));
 sky130_fd_sc_hd__nor2_1 _3934_ (.A(\game.addhits.add2.b[3] ),
    .B(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__a31o_1 _3935_ (.A1(\game.addhits.add2.b[1] ),
    .A2(\game.addhits.add2.b[0] ),
    .A3(_1244_),
    .B1(\game.addhits.add2.b[2] ),
    .X(_1260_));
 sky130_fd_sc_hd__nand2_1 _3936_ (.A(_1226_),
    .B(_1260_),
    .Y(_1261_));
 sky130_fd_sc_hd__a31o_1 _3937_ (.A1(_1253_),
    .A2(_1254_),
    .A3(_1258_),
    .B1(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__a2bb2o_1 _3938_ (.A1_N(_1259_),
    .A2_N(_1262_),
    .B1(net253),
    .B2(_1227_),
    .X(\game.scoring_button_2.next_num_hits[6] ));
 sky130_fd_sc_hd__a41o_1 _3939_ (.A1(_1256_),
    .A2(_1257_),
    .A3(_1226_),
    .A4(_1252_),
    .B1(_1227_),
    .X(_1263_));
 sky130_fd_sc_hd__a22o_1 _3940_ (.A1(_1226_),
    .A2(_1259_),
    .B1(_1263_),
    .B2(net153),
    .X(\game.scoring_button_2.next_num_hits[7] ));
 sky130_fd_sc_hd__and2_1 _3941_ (.A(\game.addhits.add3.b[0] ),
    .B(_1253_),
    .X(_1264_));
 sky130_fd_sc_hd__o21ai_1 _3942_ (.A1(\game.addhits.add3.b[0] ),
    .A2(_1253_),
    .B1(_1226_),
    .Y(_1265_));
 sky130_fd_sc_hd__a2bb2o_1 _3943_ (.A1_N(_1264_),
    .A2_N(_1265_),
    .B1(net249),
    .B2(_1227_),
    .X(\game.scoring_button_2.next_num_hits[8] ));
 sky130_fd_sc_hd__nor2_1 _3944_ (.A(\game.addhits.add3.b[1] ),
    .B(_1264_),
    .Y(_1266_));
 sky130_fd_sc_hd__and3_1 _3945_ (.A(\game.addhits.add3.b[1] ),
    .B(\game.addhits.add3.b[0] ),
    .C(_1253_),
    .X(_1267_));
 sky130_fd_sc_hd__o31a_1 _3946_ (.A1(\game.addhits.add3.b[2] ),
    .A2(\game.addhits.add3.b[1] ),
    .A3(_1264_),
    .B1(\game.addhits.add3.b[3] ),
    .X(_1268_));
 sky130_fd_sc_hd__o21ai_1 _3947_ (.A1(_1266_),
    .A2(_1267_),
    .B1(_1268_),
    .Y(_1269_));
 sky130_fd_sc_hd__o31ai_1 _3948_ (.A1(\game.addhits.add3.b[3] ),
    .A2(_1266_),
    .A3(_1267_),
    .B1(_1269_),
    .Y(_1270_));
 sky130_fd_sc_hd__a22o_1 _3949_ (.A1(net258),
    .A2(_1227_),
    .B1(_1270_),
    .B2(_1226_),
    .X(\game.scoring_button_2.next_num_hits[9] ));
 sky130_fd_sc_hd__or2_1 _3950_ (.A(\game.addhits.add3.b[2] ),
    .B(_1267_),
    .X(_1271_));
 sky130_fd_sc_hd__and2_1 _3951_ (.A(\game.addhits.add3.b[2] ),
    .B(_1267_),
    .X(_1272_));
 sky130_fd_sc_hd__mux2_1 _3952_ (.A0(_1269_),
    .A1(\game.addhits.add3.b[3] ),
    .S(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__a32o_1 _3953_ (.A1(_1226_),
    .A2(_1271_),
    .A3(_1273_),
    .B1(_1227_),
    .B2(net198),
    .X(\game.scoring_button_2.next_num_hits[10] ));
 sky130_fd_sc_hd__o21ba_1 _3954_ (.A1(\game.addhits.add3.b[3] ),
    .A2(_1272_),
    .B1_N(_1268_),
    .X(_1274_));
 sky130_fd_sc_hd__a22o_1 _3955_ (.A1(net219),
    .A2(_1227_),
    .B1(_1274_),
    .B2(_1226_),
    .X(\game.scoring_button_2.next_num_hits[11] ));
 sky130_fd_sc_hd__and2_1 _3956_ (.A(\game.addhits.add4.b[0] ),
    .B(_1268_),
    .X(_1275_));
 sky130_fd_sc_hd__o21ai_1 _3957_ (.A1(\game.addhits.add4.b[0] ),
    .A2(_1268_),
    .B1(_1226_),
    .Y(_1276_));
 sky130_fd_sc_hd__a2bb2o_1 _3958_ (.A1_N(_1275_),
    .A2_N(_1276_),
    .B1(net182),
    .B2(_1227_),
    .X(\game.scoring_button_2.next_num_hits[12] ));
 sky130_fd_sc_hd__a21oi_1 _3959_ (.A1(\game.addhits.add4.b[1] ),
    .A2(_1275_),
    .B1(\game.addhits.add4.b[2] ),
    .Y(_1277_));
 sky130_fd_sc_hd__xnor2_1 _3960_ (.A(\game.addhits.add4.b[1] ),
    .B(_1275_),
    .Y(_1278_));
 sky130_fd_sc_hd__nand2_1 _3961_ (.A(\game.addhits.add4.b[3] ),
    .B(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__or2_1 _3962_ (.A(\game.addhits.add4.b[3] ),
    .B(_1278_),
    .X(_1280_));
 sky130_fd_sc_hd__o21ai_1 _3963_ (.A1(_1277_),
    .A2(_1279_),
    .B1(_1280_),
    .Y(_1281_));
 sky130_fd_sc_hd__a22o_1 _3964_ (.A1(net190),
    .A2(_1227_),
    .B1(_1281_),
    .B2(_1226_),
    .X(\game.scoring_button_2.next_num_hits[13] ));
 sky130_fd_sc_hd__and3_1 _3965_ (.A(\game.addhits.add4.b[1] ),
    .B(\game.addhits.add4.b[2] ),
    .C(_1275_),
    .X(_1282_));
 sky130_fd_sc_hd__a21oi_1 _3966_ (.A1(_0742_),
    .A2(_1282_),
    .B1(_1277_),
    .Y(_1283_));
 sky130_fd_sc_hd__or2_1 _3967_ (.A(_1279_),
    .B(_1282_),
    .X(_1284_));
 sky130_fd_sc_hd__a32o_1 _3968_ (.A1(_1226_),
    .A2(_1283_),
    .A3(_1284_),
    .B1(_1227_),
    .B2(net213),
    .X(\game.scoring_button_2.next_num_hits[14] ));
 sky130_fd_sc_hd__a21oi_1 _3969_ (.A1(\game.addhits.add4.b[3] ),
    .A2(_1278_),
    .B1(_1282_),
    .Y(_1285_));
 sky130_fd_sc_hd__nor2_1 _3970_ (.A(_1283_),
    .B(_1285_),
    .Y(_1286_));
 sky130_fd_sc_hd__a22o_1 _3971_ (.A1(\game.addhits.add4.b[3] ),
    .A2(_1227_),
    .B1(_1286_),
    .B2(_1226_),
    .X(\game.scoring_button_2.next_num_hits[15] ));
 sky130_fd_sc_hd__inv_2 _3972_ (.A(\game.scoring_button_2.check_hit.edge_2 ),
    .Y(_1287_));
 sky130_fd_sc_hd__or3_1 _3973_ (.A(\game.scoring_button_2.check_hit.edge_1 ),
    .B(_1287_),
    .C(\game.scoring_button_2.hit ),
    .X(_1288_));
 sky130_fd_sc_hd__clkbuf_8 _3974_ (.A(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__or3_1 _3975_ (.A(\game.scoring_button_2.counts[14] ),
    .B(\game.scoring_button_2.counts[13] ),
    .C(\game.scoring_button_2.counts[12] ),
    .X(_1290_));
 sky130_fd_sc_hd__or4_1 _3976_ (.A(\game.scoring_button_2.counts[16] ),
    .B(\game.scoring_button_2.counts[15] ),
    .C(\game.scoring_button_2.counts[11] ),
    .D(\game.scoring_button_2.counts[10] ),
    .X(_1291_));
 sky130_fd_sc_hd__or4_1 _3977_ (.A(\game.scoring_button_2.counts[9] ),
    .B(\game.scoring_button_2.counts[8] ),
    .C(\game.scoring_button_2.counts[7] ),
    .D(_1291_),
    .X(_1292_));
 sky130_fd_sc_hd__or4_1 _3978_ (.A(\game.scoring_button_2.counts[6] ),
    .B(\game.scoring_button_2.counts[5] ),
    .C(\game.scoring_button_2.counts[3] ),
    .D(\game.scoring_button_2.counts[4] ),
    .X(_1293_));
 sky130_fd_sc_hd__or4_2 _3979_ (.A(\game.scoring_button_2.counts[2] ),
    .B(\game.scoring_button_2.counts[1] ),
    .C(\game.scoring_button_2.counts[0] ),
    .D(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__or4_1 _3980_ (.A(\game.scoring_button_2.counts[20] ),
    .B(\game.scoring_button_2.counts[19] ),
    .C(\game.scoring_button_2.counts[18] ),
    .D(\game.scoring_button_2.counts[17] ),
    .X(_1295_));
 sky130_fd_sc_hd__or4_1 _3981_ (.A(\game.scoring_button_2.counts[21] ),
    .B(\game.scoring_button_2.counts[22] ),
    .C(_1294_),
    .D(_1295_),
    .X(_1296_));
 sky130_fd_sc_hd__a31o_1 _3982_ (.A1(\game.scoring_button_2.counts[8] ),
    .A2(\game.scoring_button_2.counts[7] ),
    .A3(_1294_),
    .B1(\game.scoring_button_2.counts[9] ),
    .X(_1297_));
 sky130_fd_sc_hd__a31o_1 _3983_ (.A1(\game.scoring_button_2.counts[11] ),
    .A2(\game.scoring_button_2.counts[10] ),
    .A3(_1297_),
    .B1(_1290_),
    .X(_1298_));
 sky130_fd_sc_hd__a41o_1 _3984_ (.A1(\game.scoring_button_2.counts[17] ),
    .A2(\game.scoring_button_2.counts[16] ),
    .A3(\game.scoring_button_2.counts[15] ),
    .A4(_1298_),
    .B1(\game.scoring_button_2.counts[18] ),
    .X(_1299_));
 sky130_fd_sc_hd__a31o_1 _3985_ (.A1(\game.scoring_button_2.counts[20] ),
    .A2(\game.scoring_button_2.counts[19] ),
    .A3(_1299_),
    .B1(\game.scoring_button_2.counts[21] ),
    .X(_1300_));
 sky130_fd_sc_hd__nand2_1 _3986_ (.A(\game.scoring_button_2.counts[22] ),
    .B(_1300_),
    .Y(_1301_));
 sky130_fd_sc_hd__o31a_1 _3987_ (.A1(_1290_),
    .A2(_1292_),
    .A3(_1296_),
    .B1(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__nand2_2 _3988_ (.A(_0209_),
    .B(_2658_),
    .Y(_1303_));
 sky130_fd_sc_hd__or2_1 _3989_ (.A(_1302_),
    .B(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__clkbuf_4 _3990_ (.A(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__inv_2 _3991_ (.A(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hd__nor2_2 _3992_ (.A(_0208_),
    .B(_1306_),
    .Y(_1307_));
 sky130_fd_sc_hd__a21oi_1 _3993_ (.A1(_1305_),
    .A2(_1289_),
    .B1(\game.addmisses.add1.b[0] ),
    .Y(_1308_));
 sky130_fd_sc_hd__a31o_1 _3994_ (.A1(\game.addmisses.add1.b[0] ),
    .A2(_1289_),
    .A3(_1307_),
    .B1(_1308_),
    .X(\game.scoring_button_2.next_num_misses[0] ));
 sky130_fd_sc_hd__xnor2_1 _3995_ (.A(\game.addmisses.add1.b[1] ),
    .B(\game.addmisses.add1.b[0] ),
    .Y(_1309_));
 sky130_fd_sc_hd__o2bb2a_1 _3996_ (.A1_N(\game.addmisses.add1.b[1] ),
    .A2_N(_1307_),
    .B1(_1309_),
    .B2(_1305_),
    .X(_1310_));
 sky130_fd_sc_hd__o31a_1 _3997_ (.A1(\game.addmisses.add1.b[2] ),
    .A2(\game.addmisses.add1.b[1] ),
    .A3(\game.addmisses.add1.b[0] ),
    .B1(\game.addmisses.add1.b[3] ),
    .X(_1311_));
 sky130_fd_sc_hd__and2_1 _3998_ (.A(_1309_),
    .B(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__nor3_1 _3999_ (.A(\game.scoring_button_2.check_hit.edge_1 ),
    .B(_1287_),
    .C(\game.scoring_button_2.hit ),
    .Y(_1313_));
 sky130_fd_sc_hd__o21ai_1 _4000_ (.A1(\game.addmisses.add1.b[3] ),
    .A2(_1309_),
    .B1(_1313_),
    .Y(_1314_));
 sky130_fd_sc_hd__o2bb2a_1 _4001_ (.A1_N(_1289_),
    .A2_N(_1310_),
    .B1(_1312_),
    .B2(_1314_),
    .X(\game.scoring_button_2.next_num_misses[1] ));
 sky130_fd_sc_hd__and3_1 _4002_ (.A(\game.addmisses.add1.b[2] ),
    .B(\game.addmisses.add1.b[1] ),
    .C(\game.addmisses.add1.b[0] ),
    .X(_1315_));
 sky130_fd_sc_hd__a21oi_1 _4003_ (.A1(\game.addmisses.add1.b[1] ),
    .A2(\game.addmisses.add1.b[0] ),
    .B1(\game.addmisses.add1.b[2] ),
    .Y(_1316_));
 sky130_fd_sc_hd__or2_1 _4004_ (.A(_1315_),
    .B(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__nor2_1 _4005_ (.A(_1312_),
    .B(_1317_),
    .Y(_1318_));
 sky130_fd_sc_hd__and2_2 _4006_ (.A(\game.addmisses.add1.b[3] ),
    .B(_1315_),
    .X(_1319_));
 sky130_fd_sc_hd__nor2_1 _4007_ (.A(_1305_),
    .B(_1317_),
    .Y(_1320_));
 sky130_fd_sc_hd__a211o_1 _4008_ (.A1(\game.addmisses.add1.b[2] ),
    .A2(_1307_),
    .B1(_1320_),
    .C1(net45),
    .X(_1321_));
 sky130_fd_sc_hd__o31a_1 _4009_ (.A1(_1289_),
    .A2(_1318_),
    .A3(_1319_),
    .B1(_1321_),
    .X(\game.scoring_button_2.next_num_misses[2] ));
 sky130_fd_sc_hd__nor2_1 _4010_ (.A(\game.addmisses.add1.b[3] ),
    .B(_1315_),
    .Y(_1322_));
 sky130_fd_sc_hd__nor2_1 _4011_ (.A(_1319_),
    .B(_1322_),
    .Y(_1323_));
 sky130_fd_sc_hd__nor2_1 _4012_ (.A(_1289_),
    .B(_1311_),
    .Y(_1324_));
 sky130_fd_sc_hd__a22o_1 _4013_ (.A1(\game.addmisses.add1.b[3] ),
    .A2(_1307_),
    .B1(_1323_),
    .B2(_1306_),
    .X(_1325_));
 sky130_fd_sc_hd__a22o_1 _4014_ (.A1(_1323_),
    .A2(_1324_),
    .B1(_1325_),
    .B2(_1289_),
    .X(\game.scoring_button_2.next_num_misses[3] ));
 sky130_fd_sc_hd__or2_1 _4015_ (.A(\game.addmisses.add2.b[0] ),
    .B(_1311_),
    .X(_1326_));
 sky130_fd_sc_hd__and2_1 _4016_ (.A(\game.addmisses.add2.b[0] ),
    .B(_1311_),
    .X(_1327_));
 sky130_fd_sc_hd__nor2_1 _4017_ (.A(_1289_),
    .B(_1327_),
    .Y(_1328_));
 sky130_fd_sc_hd__nand2_1 _4018_ (.A(\game.addmisses.add2.b[0] ),
    .B(_1319_),
    .Y(_1329_));
 sky130_fd_sc_hd__nand2_1 _4019_ (.A(\modetrans.mode[0] ),
    .B(_1305_),
    .Y(_1330_));
 sky130_fd_sc_hd__o21a_1 _4020_ (.A1(_1305_),
    .A2(_1329_),
    .B1(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__or3b_1 _4021_ (.A(\game.addmisses.add2.b[0] ),
    .B(_1305_),
    .C_N(_1319_),
    .X(_1332_));
 sky130_fd_sc_hd__a21bo_1 _4022_ (.A1(\game.addmisses.add2.b[0] ),
    .A2(_1331_),
    .B1_N(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__a22o_1 _4023_ (.A1(_1326_),
    .A2(_1328_),
    .B1(_1333_),
    .B2(_1289_),
    .X(\game.scoring_button_2.next_num_misses[4] ));
 sky130_fd_sc_hd__or2_1 _4024_ (.A(\game.addmisses.add2.b[1] ),
    .B(_1327_),
    .X(_1334_));
 sky130_fd_sc_hd__o21a_2 _4025_ (.A1(\game.addmisses.add2.b[2] ),
    .A2(_1334_),
    .B1(\game.addmisses.add2.b[3] ),
    .X(_1335_));
 sky130_fd_sc_hd__nand2_1 _4026_ (.A(\game.addmisses.add2.b[1] ),
    .B(_1327_),
    .Y(_1336_));
 sky130_fd_sc_hd__nand2_1 _4027_ (.A(_1334_),
    .B(_1336_),
    .Y(_1337_));
 sky130_fd_sc_hd__xor2_1 _4028_ (.A(_1335_),
    .B(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__nand2_1 _4029_ (.A(\game.addmisses.add2.b[1] ),
    .B(_1331_),
    .Y(_1339_));
 sky130_fd_sc_hd__o311a_1 _4030_ (.A1(\game.addmisses.add2.b[1] ),
    .A2(_1305_),
    .A3(_1329_),
    .B1(_1339_),
    .C1(_1289_),
    .X(_1340_));
 sky130_fd_sc_hd__a21oi_1 _4031_ (.A1(net45),
    .A2(_1338_),
    .B1(_1340_),
    .Y(\game.scoring_button_2.next_num_misses[5] ));
 sky130_fd_sc_hd__inv_2 _4032_ (.A(_1335_),
    .Y(_1341_));
 sky130_fd_sc_hd__a22o_1 _4033_ (.A1(\game.addmisses.add2.b[3] ),
    .A2(_1334_),
    .B1(_1341_),
    .B2(_1336_),
    .X(_1342_));
 sky130_fd_sc_hd__xnor2_1 _4034_ (.A(\game.addmisses.add2.b[2] ),
    .B(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__and4_1 _4035_ (.A(\game.addmisses.add2.b[2] ),
    .B(\game.addmisses.add2.b[1] ),
    .C(\game.addmisses.add2.b[0] ),
    .D(_1319_),
    .X(_1344_));
 sky130_fd_sc_hd__a31o_1 _4036_ (.A1(\game.addmisses.add2.b[1] ),
    .A2(\game.addmisses.add2.b[0] ),
    .A3(_1319_),
    .B1(\game.addmisses.add2.b[2] ),
    .X(_1345_));
 sky130_fd_sc_hd__or3b_1 _4037_ (.A(_1305_),
    .B(_1344_),
    .C_N(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__a21bo_1 _4038_ (.A1(\game.addmisses.add2.b[2] ),
    .A2(_1307_),
    .B1_N(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__mux2_1 _4039_ (.A0(_1343_),
    .A1(_1347_),
    .S(_1289_),
    .X(_1348_));
 sky130_fd_sc_hd__clkbuf_1 _4040_ (.A(_1348_),
    .X(\game.scoring_button_2.next_num_misses[6] ));
 sky130_fd_sc_hd__a31o_1 _4041_ (.A1(\game.addmisses.add2.b[2] ),
    .A2(\game.addmisses.add2.b[1] ),
    .A3(_1327_),
    .B1(\game.addmisses.add2.b[3] ),
    .X(_1349_));
 sky130_fd_sc_hd__nor2_1 _4042_ (.A(_1289_),
    .B(_1335_),
    .Y(_1350_));
 sky130_fd_sc_hd__nand2_1 _4043_ (.A(\game.addmisses.add2.b[3] ),
    .B(_1344_),
    .Y(_1351_));
 sky130_fd_sc_hd__or2_1 _4044_ (.A(\game.addmisses.add2.b[3] ),
    .B(_1344_),
    .X(_1352_));
 sky130_fd_sc_hd__a32o_1 _4045_ (.A1(_1306_),
    .A2(_1351_),
    .A3(_1352_),
    .B1(_1307_),
    .B2(\game.addmisses.add2.b[3] ),
    .X(_1353_));
 sky130_fd_sc_hd__a22o_1 _4046_ (.A1(_1349_),
    .A2(_1350_),
    .B1(_1353_),
    .B2(_1289_),
    .X(\game.scoring_button_2.next_num_misses[7] ));
 sky130_fd_sc_hd__or2_1 _4047_ (.A(\game.addmisses.add3.b[0] ),
    .B(_1335_),
    .X(_1354_));
 sky130_fd_sc_hd__and2_1 _4048_ (.A(\game.addmisses.add3.b[0] ),
    .B(_1335_),
    .X(_1355_));
 sky130_fd_sc_hd__inv_2 _4049_ (.A(_1355_),
    .Y(_1356_));
 sky130_fd_sc_hd__nor2_2 _4050_ (.A(_1305_),
    .B(_1351_),
    .Y(_1357_));
 sky130_fd_sc_hd__and2_1 _4051_ (.A(\modetrans.mode[0] ),
    .B(_1305_),
    .X(_1358_));
 sky130_fd_sc_hd__o21ai_1 _4052_ (.A1(_1358_),
    .A2(_1357_),
    .B1(\game.addmisses.add3.b[0] ),
    .Y(_1359_));
 sky130_fd_sc_hd__o211a_1 _4053_ (.A1(\game.addmisses.add3.b[0] ),
    .A2(_1357_),
    .B1(_1359_),
    .C1(_1289_),
    .X(_1360_));
 sky130_fd_sc_hd__a31o_1 _4054_ (.A1(net45),
    .A2(_1354_),
    .A3(_1356_),
    .B1(_1360_),
    .X(\game.scoring_button_2.next_num_misses[8] ));
 sky130_fd_sc_hd__nand2_1 _4055_ (.A(\game.addmisses.add3.b[1] ),
    .B(_1355_),
    .Y(_1361_));
 sky130_fd_sc_hd__or2_1 _4056_ (.A(\game.addmisses.add3.b[1] ),
    .B(_1355_),
    .X(_1362_));
 sky130_fd_sc_hd__o21a_1 _4057_ (.A1(\game.addmisses.add3.b[2] ),
    .A2(_1362_),
    .B1(\game.addmisses.add3.b[3] ),
    .X(_1363_));
 sky130_fd_sc_hd__a21boi_1 _4058_ (.A1(_1361_),
    .A2(_1362_),
    .B1_N(_1363_),
    .Y(_1364_));
 sky130_fd_sc_hd__and3b_1 _4059_ (.A_N(\game.addmisses.add3.b[3] ),
    .B(_1361_),
    .C(_1362_),
    .X(_1365_));
 sky130_fd_sc_hd__nand2_1 _4060_ (.A(\game.addmisses.add3.b[0] ),
    .B(_1357_),
    .Y(_1366_));
 sky130_fd_sc_hd__o21ai_1 _4061_ (.A1(\game.addmisses.add3.b[1] ),
    .A2(_1366_),
    .B1(_1289_),
    .Y(_1367_));
 sky130_fd_sc_hd__a31o_1 _4062_ (.A1(\game.addmisses.add3.b[1] ),
    .A2(_1330_),
    .A3(_1366_),
    .B1(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__o31a_1 _4063_ (.A1(_1289_),
    .A2(_1364_),
    .A3(_1365_),
    .B1(_1368_),
    .X(\game.scoring_button_2.next_num_misses[9] ));
 sky130_fd_sc_hd__and3_1 _4064_ (.A(\game.addmisses.add3.b[2] ),
    .B(\game.addmisses.add3.b[1] ),
    .C(_1355_),
    .X(_1369_));
 sky130_fd_sc_hd__a21oi_1 _4065_ (.A1(\game.addmisses.add3.b[1] ),
    .A2(_1355_),
    .B1(\game.addmisses.add3.b[2] ),
    .Y(_1370_));
 sky130_fd_sc_hd__or2_1 _4066_ (.A(_1369_),
    .B(_1370_),
    .X(_1371_));
 sky130_fd_sc_hd__a2bb2o_1 _4067_ (.A1_N(_1364_),
    .A2_N(_1371_),
    .B1(_1369_),
    .B2(\game.addmisses.add3.b[3] ),
    .X(_1372_));
 sky130_fd_sc_hd__a32o_1 _4068_ (.A1(\game.addmisses.add3.b[1] ),
    .A2(\game.addmisses.add3.b[0] ),
    .A3(_1357_),
    .B1(_1330_),
    .B2(\game.addmisses.add3.b[2] ),
    .X(_1373_));
 sky130_fd_sc_hd__and4_1 _4069_ (.A(\game.addmisses.add3.b[2] ),
    .B(\game.addmisses.add3.b[1] ),
    .C(\game.addmisses.add3.b[0] ),
    .D(_1357_),
    .X(_1374_));
 sky130_fd_sc_hd__nor2_1 _4070_ (.A(net45),
    .B(_1374_),
    .Y(_1375_));
 sky130_fd_sc_hd__a22o_1 _4071_ (.A1(net45),
    .A2(_1372_),
    .B1(_1373_),
    .B2(_1375_),
    .X(\game.scoring_button_2.next_num_misses[10] ));
 sky130_fd_sc_hd__nor2_1 _4072_ (.A(\game.addmisses.add3.b[2] ),
    .B(_1362_),
    .Y(_1376_));
 sky130_fd_sc_hd__nor2_1 _4073_ (.A(_1358_),
    .B(_1374_),
    .Y(_1377_));
 sky130_fd_sc_hd__mux4_1 _4074_ (.A0(_1369_),
    .A1(_1374_),
    .A2(_1376_),
    .A3(_1377_),
    .S0(_1289_),
    .S1(\game.addmisses.add3.b[3] ),
    .X(_1378_));
 sky130_fd_sc_hd__clkbuf_1 _4075_ (.A(_1378_),
    .X(\game.scoring_button_2.next_num_misses[11] ));
 sky130_fd_sc_hd__and2_1 _4076_ (.A(\game.addmisses.add4.b[0] ),
    .B(_1363_),
    .X(_1379_));
 sky130_fd_sc_hd__nor2_1 _4077_ (.A(\game.addmisses.add4.b[0] ),
    .B(_1363_),
    .Y(_1380_));
 sky130_fd_sc_hd__and3_1 _4078_ (.A(\game.addmisses.add3.b[3] ),
    .B(_1357_),
    .C(_1369_),
    .X(_1381_));
 sky130_fd_sc_hd__nor2_1 _4079_ (.A(\game.addmisses.add4.b[0] ),
    .B(_1381_),
    .Y(_1382_));
 sky130_fd_sc_hd__nand2_1 _4080_ (.A(\game.addmisses.add4.b[0] ),
    .B(_1381_),
    .Y(_1383_));
 sky130_fd_sc_hd__or4b_1 _4081_ (.A(net45),
    .B(_1358_),
    .C(_1382_),
    .D_N(_1383_),
    .X(_1384_));
 sky130_fd_sc_hd__o31ai_1 _4082_ (.A1(_1289_),
    .A2(_1379_),
    .A3(_1380_),
    .B1(_1384_),
    .Y(\game.scoring_button_2.next_num_misses[12] ));
 sky130_fd_sc_hd__and3_2 _4083_ (.A(\game.addmisses.add4.b[0] ),
    .B(\game.addmisses.add4.b[1] ),
    .C(_1363_),
    .X(_1385_));
 sky130_fd_sc_hd__nor2_1 _4084_ (.A(\game.addmisses.add4.b[1] ),
    .B(_1379_),
    .Y(_1386_));
 sky130_fd_sc_hd__or2_1 _4085_ (.A(_1385_),
    .B(_1386_),
    .X(_1387_));
 sky130_fd_sc_hd__nand2_1 _4086_ (.A(\game.addmisses.add4.b[3] ),
    .B(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__o21bai_1 _4087_ (.A1(\game.addmisses.add4.b[2] ),
    .A2(_1385_),
    .B1_N(_1388_),
    .Y(_1389_));
 sky130_fd_sc_hd__o21ai_1 _4088_ (.A1(\game.addmisses.add4.b[3] ),
    .A2(_1387_),
    .B1(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__and3_1 _4089_ (.A(\game.addmisses.add4.b[1] ),
    .B(_1330_),
    .C(_1383_),
    .X(_1391_));
 sky130_fd_sc_hd__o21ai_1 _4090_ (.A1(\game.addmisses.add4.b[1] ),
    .A2(_1383_),
    .B1(_1289_),
    .Y(_1392_));
 sky130_fd_sc_hd__o22a_1 _4091_ (.A1(_1289_),
    .A2(_1390_),
    .B1(_1391_),
    .B2(_1392_),
    .X(\game.scoring_button_2.next_num_misses[13] ));
 sky130_fd_sc_hd__and2_1 _4092_ (.A(_1381_),
    .B(_1385_),
    .X(_1393_));
 sky130_fd_sc_hd__and3_1 _4093_ (.A(\game.addmisses.add4.b[2] ),
    .B(_1381_),
    .C(_1385_),
    .X(_1394_));
 sky130_fd_sc_hd__or2_1 _4094_ (.A(_1358_),
    .B(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__o21ba_1 _4095_ (.A1(\game.addmisses.add4.b[2] ),
    .A2(_1393_),
    .B1_N(_1395_),
    .X(_1396_));
 sky130_fd_sc_hd__o21a_1 _4096_ (.A1(\game.addmisses.add4.b[2] ),
    .A2(_1385_),
    .B1(_1388_),
    .X(_1397_));
 sky130_fd_sc_hd__nand2_1 _4097_ (.A(\game.addmisses.add4.b[2] ),
    .B(_1385_),
    .Y(_1398_));
 sky130_fd_sc_hd__mux2_1 _4098_ (.A0(\game.addmisses.add4.b[3] ),
    .A1(_1397_),
    .S(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__mux2_1 _4099_ (.A0(_1396_),
    .A1(_1399_),
    .S(net45),
    .X(_1400_));
 sky130_fd_sc_hd__clkbuf_1 _4100_ (.A(_1400_),
    .X(\game.scoring_button_2.next_num_misses[14] ));
 sky130_fd_sc_hd__or3_1 _4101_ (.A(\game.addmisses.add4.b[2] ),
    .B(\game.addmisses.add4.b[1] ),
    .C(_1379_),
    .X(_1401_));
 sky130_fd_sc_hd__mux2_1 _4102_ (.A0(_1398_),
    .A1(_1401_),
    .S(\game.addmisses.add4.b[3] ),
    .X(_1402_));
 sky130_fd_sc_hd__nor2_1 _4103_ (.A(\game.addmisses.add4.b[3] ),
    .B(_1394_),
    .Y(_1403_));
 sky130_fd_sc_hd__a211o_1 _4104_ (.A1(\game.addmisses.add4.b[3] ),
    .A2(_1395_),
    .B1(_1403_),
    .C1(net45),
    .X(_1404_));
 sky130_fd_sc_hd__o21ai_1 _4105_ (.A1(_1289_),
    .A2(_1402_),
    .B1(_1404_),
    .Y(\game.scoring_button_2.next_num_misses[15] ));
 sky130_fd_sc_hd__clkbuf_8 _4106_ (.A(\game.scoring_button_2.check_hit.in ),
    .X(_1405_));
 sky130_fd_sc_hd__or4b_1 _4107_ (.A(\game.scoring_button_2.flash_counter_1[5] ),
    .B(\game.scoring_button_2.flash_counter_1[4] ),
    .C(\game.scoring_button_2.flash_counter_1[7] ),
    .D_N(\game.scoring_button_2.flash_counter_1[6] ),
    .X(_1406_));
 sky130_fd_sc_hd__or4_1 _4108_ (.A(\game.scoring_button_2.flash_counter_1[1] ),
    .B(\game.scoring_button_2.flash_counter_1[0] ),
    .C(\game.scoring_button_2.flash_counter_1[3] ),
    .D(\game.scoring_button_2.flash_counter_1[2] ),
    .X(_1407_));
 sky130_fd_sc_hd__or4b_1 _4109_ (.A(\game.scoring_button_2.flash_counter_1[13] ),
    .B(\game.scoring_button_2.flash_counter_1[12] ),
    .C(\game.scoring_button_2.flash_counter_1[15] ),
    .D_N(\game.scoring_button_2.flash_counter_1[14] ),
    .X(_1408_));
 sky130_fd_sc_hd__or4b_1 _4110_ (.A(\game.scoring_button_2.flash_counter_1[8] ),
    .B(\game.scoring_button_2.flash_counter_1[11] ),
    .C(\game.scoring_button_2.flash_counter_1[10] ),
    .D_N(\game.scoring_button_2.flash_counter_1[9] ),
    .X(_1409_));
 sky130_fd_sc_hd__or3_1 _4111_ (.A(\game.scoring_button_2.flash_counter_1[21] ),
    .B(\game.scoring_button_2.flash_counter_1[20] ),
    .C(\game.scoring_button_2.flash_counter_1[22] ),
    .X(_1410_));
 sky130_fd_sc_hd__and4_1 _4112_ (.A(\game.scoring_button_2.flash_counter_1[17] ),
    .B(\game.scoring_button_2.flash_counter_1[16] ),
    .C(\game.scoring_button_2.flash_counter_1[19] ),
    .D(\game.scoring_button_2.flash_counter_1[18] ),
    .X(_1411_));
 sky130_fd_sc_hd__or4b_1 _4113_ (.A(_1408_),
    .B(_1409_),
    .C(_1410_),
    .D_N(_1411_),
    .X(_1412_));
 sky130_fd_sc_hd__o31a_4 _4114_ (.A1(_1406_),
    .A2(_1407_),
    .A3(_1412_),
    .B1(\game.hit_2 ),
    .X(_1413_));
 sky130_fd_sc_hd__a31o_1 _4115_ (.A1(_0219_),
    .A2(_1405_),
    .A3(_2658_),
    .B1(_1413_),
    .X(\game.scoring_button_2.next_good ));
 sky130_fd_sc_hd__and2b_1 _4116_ (.A_N(\game.counter[0] ),
    .B(\game.scoring_button_2.check_hit.in ),
    .X(_1414_));
 sky130_fd_sc_hd__clkbuf_1 _4117_ (.A(_1414_),
    .X(\game.scoring_button_2.next_count[0] ));
 sky130_fd_sc_hd__nand2_1 _4118_ (.A(\game.counter[1] ),
    .B(\game.counter[0] ),
    .Y(_1415_));
 sky130_fd_sc_hd__and3_1 _4119_ (.A(\game.scoring_button_2.check_hit.in ),
    .B(_0248_),
    .C(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__clkbuf_1 _4120_ (.A(_1416_),
    .X(\game.scoring_button_2.next_count[1] ));
 sky130_fd_sc_hd__xnor2_1 _4121_ (.A(net199),
    .B(_1415_),
    .Y(_0024_));
 sky130_fd_sc_hd__and2_1 _4122_ (.A(_1405_),
    .B(_0024_),
    .X(_1417_));
 sky130_fd_sc_hd__clkbuf_1 _4123_ (.A(_1417_),
    .X(\game.scoring_button_2.next_count[2] ));
 sky130_fd_sc_hd__and4_1 _4124_ (.A(\game.counter[1] ),
    .B(\game.counter[0] ),
    .C(\game.counter[3] ),
    .D(\game.counter[2] ),
    .X(_1418_));
 sky130_fd_sc_hd__a31o_1 _4125_ (.A1(\game.counter[1] ),
    .A2(\game.counter[0] ),
    .A3(\game.counter[2] ),
    .B1(\game.counter[3] ),
    .X(_1419_));
 sky130_fd_sc_hd__and2b_1 _4126_ (.A_N(_1418_),
    .B(_1419_),
    .X(_1420_));
 sky130_fd_sc_hd__buf_1 _4127_ (.A(_1420_),
    .X(_0025_));
 sky130_fd_sc_hd__and2_1 _4128_ (.A(_1405_),
    .B(_0025_),
    .X(_1421_));
 sky130_fd_sc_hd__clkbuf_1 _4129_ (.A(_1421_),
    .X(\game.scoring_button_2.next_count[3] ));
 sky130_fd_sc_hd__xor2_1 _4130_ (.A(net168),
    .B(_1418_),
    .X(_0026_));
 sky130_fd_sc_hd__and2_1 _4131_ (.A(_1405_),
    .B(_0026_),
    .X(_1422_));
 sky130_fd_sc_hd__clkbuf_1 _4132_ (.A(_1422_),
    .X(\game.scoring_button_2.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _4133_ (.A(\game.counter[5] ),
    .B(\game.counter[4] ),
    .C(_1418_),
    .X(_1423_));
 sky130_fd_sc_hd__a21oi_1 _4134_ (.A1(\game.counter[4] ),
    .A2(_1418_),
    .B1(\game.counter[5] ),
    .Y(_1424_));
 sky130_fd_sc_hd__nor2_1 _4135_ (.A(_1423_),
    .B(_1424_),
    .Y(_0027_));
 sky130_fd_sc_hd__and2_1 _4136_ (.A(_1405_),
    .B(_0027_),
    .X(_1425_));
 sky130_fd_sc_hd__clkbuf_1 _4137_ (.A(_1425_),
    .X(\game.scoring_button_2.next_count[5] ));
 sky130_fd_sc_hd__xor2_1 _4138_ (.A(\game.counter[6] ),
    .B(_1423_),
    .X(_1426_));
 sky130_fd_sc_hd__and2_1 _4139_ (.A(_1405_),
    .B(_1426_),
    .X(_1427_));
 sky130_fd_sc_hd__clkbuf_1 _4140_ (.A(_1427_),
    .X(\game.scoring_button_2.next_count[6] ));
 sky130_fd_sc_hd__a21oi_1 _4141_ (.A1(\game.counter[6] ),
    .A2(_1423_),
    .B1(\game.counter[7] ),
    .Y(_1428_));
 sky130_fd_sc_hd__and3_1 _4142_ (.A(\game.counter[6] ),
    .B(\game.counter[7] ),
    .C(_1423_),
    .X(_1429_));
 sky130_fd_sc_hd__nor2_1 _4143_ (.A(_1428_),
    .B(_1429_),
    .Y(_1430_));
 sky130_fd_sc_hd__and2_1 _4144_ (.A(_1405_),
    .B(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__clkbuf_1 _4145_ (.A(_1431_),
    .X(\game.scoring_button_2.next_count[7] ));
 sky130_fd_sc_hd__xor2_1 _4146_ (.A(\game.counter[8] ),
    .B(_1429_),
    .X(_1432_));
 sky130_fd_sc_hd__and2_1 _4147_ (.A(_1405_),
    .B(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__clkbuf_1 _4148_ (.A(_1433_),
    .X(\game.scoring_button_2.next_count[8] ));
 sky130_fd_sc_hd__a21oi_1 _4149_ (.A1(\game.counter[8] ),
    .A2(_1429_),
    .B1(\game.counter[9] ),
    .Y(_1434_));
 sky130_fd_sc_hd__and3_1 _4150_ (.A(\game.counter[8] ),
    .B(\game.counter[9] ),
    .C(_1429_),
    .X(_1435_));
 sky130_fd_sc_hd__nor2_1 _4151_ (.A(_1434_),
    .B(_1435_),
    .Y(_1436_));
 sky130_fd_sc_hd__and2_1 _4152_ (.A(_1405_),
    .B(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__clkbuf_1 _4153_ (.A(_1437_),
    .X(\game.scoring_button_2.next_count[9] ));
 sky130_fd_sc_hd__nor2_1 _4154_ (.A(\game.counter[10] ),
    .B(_1435_),
    .Y(_1438_));
 sky130_fd_sc_hd__and2_1 _4155_ (.A(\game.counter[10] ),
    .B(_1435_),
    .X(_1439_));
 sky130_fd_sc_hd__nor2_1 _4156_ (.A(_1438_),
    .B(_1439_),
    .Y(_1440_));
 sky130_fd_sc_hd__and2_1 _4157_ (.A(_1405_),
    .B(_1440_),
    .X(_1441_));
 sky130_fd_sc_hd__clkbuf_1 _4158_ (.A(_1441_),
    .X(\game.scoring_button_2.next_count[10] ));
 sky130_fd_sc_hd__or2_1 _4159_ (.A(\game.counter[11] ),
    .B(_1439_),
    .X(_1442_));
 sky130_fd_sc_hd__nand2_2 _4160_ (.A(\game.counter[11] ),
    .B(_1439_),
    .Y(_1443_));
 sky130_fd_sc_hd__and3_1 _4161_ (.A(\game.scoring_button_2.check_hit.in ),
    .B(_1442_),
    .C(_1443_),
    .X(_1444_));
 sky130_fd_sc_hd__clkbuf_1 _4162_ (.A(_1444_),
    .X(\game.scoring_button_2.next_count[11] ));
 sky130_fd_sc_hd__xnor2_1 _4163_ (.A(net144),
    .B(_1443_),
    .Y(_0012_));
 sky130_fd_sc_hd__and2_1 _4164_ (.A(_1405_),
    .B(_0012_),
    .X(_1445_));
 sky130_fd_sc_hd__clkbuf_1 _4165_ (.A(_1445_),
    .X(\game.scoring_button_2.next_count[12] ));
 sky130_fd_sc_hd__nand2_1 _4166_ (.A(\game.counter[13] ),
    .B(\game.counter[12] ),
    .Y(_1446_));
 sky130_fd_sc_hd__a31o_1 _4167_ (.A1(\game.counter[11] ),
    .A2(\game.counter[12] ),
    .A3(_1439_),
    .B1(\game.counter[13] ),
    .X(_1447_));
 sky130_fd_sc_hd__o21a_1 _4168_ (.A1(_1443_),
    .A2(_1446_),
    .B1(_1447_),
    .X(_0013_));
 sky130_fd_sc_hd__and2_1 _4169_ (.A(_1405_),
    .B(_0013_),
    .X(_1448_));
 sky130_fd_sc_hd__clkbuf_1 _4170_ (.A(_1448_),
    .X(\game.scoring_button_2.next_count[13] ));
 sky130_fd_sc_hd__nor2_1 _4171_ (.A(_1443_),
    .B(_1446_),
    .Y(_1449_));
 sky130_fd_sc_hd__nor2_1 _4172_ (.A(\game.counter[14] ),
    .B(_1449_),
    .Y(_1450_));
 sky130_fd_sc_hd__and2_1 _4173_ (.A(\game.counter[14] ),
    .B(_1449_),
    .X(_1451_));
 sky130_fd_sc_hd__nor2_1 _4174_ (.A(_1450_),
    .B(_1451_),
    .Y(_1452_));
 sky130_fd_sc_hd__and2_1 _4175_ (.A(_1405_),
    .B(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__clkbuf_1 _4176_ (.A(_1453_),
    .X(\game.scoring_button_2.next_count[14] ));
 sky130_fd_sc_hd__xnor2_1 _4177_ (.A(_0240_),
    .B(_1451_),
    .Y(_1454_));
 sky130_fd_sc_hd__and2_1 _4178_ (.A(_1405_),
    .B(_1454_),
    .X(_1455_));
 sky130_fd_sc_hd__clkbuf_1 _4179_ (.A(_1455_),
    .X(\game.scoring_button_2.next_count[15] ));
 sky130_fd_sc_hd__a21oi_1 _4180_ (.A1(\game.counter[15] ),
    .A2(_1451_),
    .B1(\game.counter[16] ),
    .Y(_1456_));
 sky130_fd_sc_hd__and3_1 _4181_ (.A(\game.counter[15] ),
    .B(\game.counter[16] ),
    .C(_1451_),
    .X(_1457_));
 sky130_fd_sc_hd__nor2_1 _4182_ (.A(_1456_),
    .B(_1457_),
    .Y(_1458_));
 sky130_fd_sc_hd__and2_1 _4183_ (.A(_1405_),
    .B(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__clkbuf_1 _4184_ (.A(_1459_),
    .X(\game.scoring_button_2.next_count[16] ));
 sky130_fd_sc_hd__nor2_1 _4185_ (.A(\game.counter[17] ),
    .B(_1457_),
    .Y(_1460_));
 sky130_fd_sc_hd__and2_1 _4186_ (.A(\game.counter[17] ),
    .B(_1457_),
    .X(_1461_));
 sky130_fd_sc_hd__nor2_1 _4187_ (.A(_1460_),
    .B(_1461_),
    .Y(_0017_));
 sky130_fd_sc_hd__and2_1 _4188_ (.A(_1405_),
    .B(_0017_),
    .X(_1462_));
 sky130_fd_sc_hd__clkbuf_1 _4189_ (.A(_1462_),
    .X(\game.scoring_button_2.next_count[17] ));
 sky130_fd_sc_hd__xor2_1 _4190_ (.A(\game.counter[18] ),
    .B(_1461_),
    .X(_1463_));
 sky130_fd_sc_hd__and2_1 _4191_ (.A(_1405_),
    .B(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__clkbuf_1 _4192_ (.A(_1464_),
    .X(\game.scoring_button_2.next_count[18] ));
 sky130_fd_sc_hd__a21oi_1 _4193_ (.A1(\game.counter[18] ),
    .A2(_1461_),
    .B1(\game.counter[19] ),
    .Y(_1465_));
 sky130_fd_sc_hd__and3_1 _4194_ (.A(\game.counter[19] ),
    .B(\game.counter[18] ),
    .C(_1461_),
    .X(_1466_));
 sky130_fd_sc_hd__nor2_1 _4195_ (.A(_1465_),
    .B(_1466_),
    .Y(_1467_));
 sky130_fd_sc_hd__and2_1 _4196_ (.A(_1405_),
    .B(_1467_),
    .X(_1468_));
 sky130_fd_sc_hd__clkbuf_1 _4197_ (.A(_1468_),
    .X(\game.scoring_button_2.next_count[19] ));
 sky130_fd_sc_hd__nor2_1 _4198_ (.A(\game.counter[20] ),
    .B(_1466_),
    .Y(_1469_));
 sky130_fd_sc_hd__and2_1 _4199_ (.A(\game.counter[20] ),
    .B(_1466_),
    .X(_1470_));
 sky130_fd_sc_hd__nor2_1 _4200_ (.A(_1469_),
    .B(_1470_),
    .Y(_1471_));
 sky130_fd_sc_hd__and2_1 _4201_ (.A(\game.scoring_button_2.check_hit.in ),
    .B(_1471_),
    .X(_1472_));
 sky130_fd_sc_hd__clkbuf_1 _4202_ (.A(_1472_),
    .X(\game.scoring_button_2.next_count[20] ));
 sky130_fd_sc_hd__or2_1 _4203_ (.A(\game.counter[21] ),
    .B(_1470_),
    .X(_1473_));
 sky130_fd_sc_hd__nand2_1 _4204_ (.A(\game.counter[21] ),
    .B(_1470_),
    .Y(_1474_));
 sky130_fd_sc_hd__and2_1 _4205_ (.A(_1473_),
    .B(_1474_),
    .X(_1475_));
 sky130_fd_sc_hd__and2_1 _4206_ (.A(\game.scoring_button_2.check_hit.in ),
    .B(_1475_),
    .X(_1476_));
 sky130_fd_sc_hd__clkbuf_1 _4207_ (.A(_1476_),
    .X(\game.scoring_button_2.next_count[21] ));
 sky130_fd_sc_hd__xnor2_1 _4208_ (.A(\game.counter[22] ),
    .B(_1474_),
    .Y(_1477_));
 sky130_fd_sc_hd__and2_1 _4209_ (.A(\game.scoring_button_2.check_hit.in ),
    .B(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__clkbuf_1 _4210_ (.A(_1478_),
    .X(\game.scoring_button_2.next_count[22] ));
 sky130_fd_sc_hd__or4b_1 _4211_ (.A(\game.scoring_button_2.flash_counter_2[5] ),
    .B(\game.scoring_button_2.flash_counter_2[4] ),
    .C(\game.scoring_button_2.flash_counter_2[7] ),
    .D_N(\game.scoring_button_2.flash_counter_2[6] ),
    .X(_1479_));
 sky130_fd_sc_hd__or4_1 _4212_ (.A(\game.scoring_button_2.flash_counter_2[1] ),
    .B(\game.scoring_button_2.flash_counter_2[0] ),
    .C(\game.scoring_button_2.flash_counter_2[3] ),
    .D(\game.scoring_button_2.flash_counter_2[2] ),
    .X(_1480_));
 sky130_fd_sc_hd__or4b_1 _4213_ (.A(\game.scoring_button_2.flash_counter_2[13] ),
    .B(\game.scoring_button_2.flash_counter_2[12] ),
    .C(\game.scoring_button_2.flash_counter_2[15] ),
    .D_N(\game.scoring_button_2.flash_counter_2[14] ),
    .X(_1481_));
 sky130_fd_sc_hd__or4b_1 _4214_ (.A(\game.scoring_button_2.flash_counter_2[8] ),
    .B(\game.scoring_button_2.flash_counter_2[11] ),
    .C(\game.scoring_button_2.flash_counter_2[10] ),
    .D_N(\game.scoring_button_2.flash_counter_2[9] ),
    .X(_1482_));
 sky130_fd_sc_hd__or3_1 _4215_ (.A(\game.scoring_button_2.flash_counter_2[21] ),
    .B(\game.scoring_button_2.flash_counter_2[20] ),
    .C(\game.scoring_button_2.flash_counter_2[22] ),
    .X(_1483_));
 sky130_fd_sc_hd__and4_1 _4216_ (.A(\game.scoring_button_2.flash_counter_2[17] ),
    .B(\game.scoring_button_2.flash_counter_2[16] ),
    .C(\game.scoring_button_2.flash_counter_2[19] ),
    .D(\game.scoring_button_2.flash_counter_2[18] ),
    .X(_1484_));
 sky130_fd_sc_hd__or4b_1 _4217_ (.A(_1481_),
    .B(_1482_),
    .C(_1483_),
    .D_N(_1484_),
    .X(_1485_));
 sky130_fd_sc_hd__o31a_2 _4218_ (.A1(_1479_),
    .A2(_1480_),
    .A3(_1485_),
    .B1(\game.missed_2 ),
    .X(_1486_));
 sky130_fd_sc_hd__o21bai_1 _4219_ (.A1(_1405_),
    .A2(_1303_),
    .B1_N(_1486_),
    .Y(\game.scoring_button_2.next_missed ));
 sky130_fd_sc_hd__nand2_1 _4220_ (.A(\game.counter[6] ),
    .B(\game.counter[7] ),
    .Y(_1487_));
 sky130_fd_sc_hd__or4b_1 _4221_ (.A(\game.counter[4] ),
    .B(\game.counter[16] ),
    .C(\game.counter[17] ),
    .D_N(\game.counter[5] ),
    .X(_1488_));
 sky130_fd_sc_hd__or4_1 _4222_ (.A(\game.counter[13] ),
    .B(\game.counter[12] ),
    .C(_1487_),
    .D(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__or4_1 _4223_ (.A(_0237_),
    .B(_0240_),
    .C(\game.counter[19] ),
    .D(\game.counter[18] ),
    .X(_1490_));
 sky130_fd_sc_hd__or4b_1 _4224_ (.A(\game.counter[8] ),
    .B(\game.counter[9] ),
    .C(\game.counter[10] ),
    .D_N(\game.counter[11] ),
    .X(_1491_));
 sky130_fd_sc_hd__or3b_1 _4225_ (.A(\game.counter[21] ),
    .B(\game.counter[22] ),
    .C_N(\game.counter[20] ),
    .X(_1492_));
 sky130_fd_sc_hd__or4_1 _4226_ (.A(_0249_),
    .B(_1490_),
    .C(_1491_),
    .D(_1492_),
    .X(_1493_));
 sky130_fd_sc_hd__nor2_1 _4227_ (.A(_1489_),
    .B(_1493_),
    .Y(_1494_));
 sky130_fd_sc_hd__inv_2 _4228_ (.A(_1494_),
    .Y(_1495_));
 sky130_fd_sc_hd__a21o_1 _4229_ (.A1(\game.counter[9] ),
    .A2(_0243_),
    .B1(\game.counter[14] ),
    .X(_1496_));
 sky130_fd_sc_hd__o22a_1 _4230_ (.A1(\game.counter[16] ),
    .A2(\game.counter[17] ),
    .B1(\game.counter[18] ),
    .B2(_0245_),
    .X(_1497_));
 sky130_fd_sc_hd__inv_2 _4231_ (.A(\game.counter[21] ),
    .Y(_1498_));
 sky130_fd_sc_hd__o31a_1 _4232_ (.A1(\game.counter[13] ),
    .A2(\game.counter[12] ),
    .A3(_1498_),
    .B1(_0227_),
    .X(_1499_));
 sky130_fd_sc_hd__a211oi_1 _4233_ (.A1(_0241_),
    .A2(_1446_),
    .B1(_1497_),
    .C1(_1499_),
    .Y(_1500_));
 sky130_fd_sc_hd__and4bb_1 _4234_ (.A_N(\game.counter[4] ),
    .B_N(\game.counter[22] ),
    .C(\game.counter[19] ),
    .D(\game.counter[5] ),
    .X(_1501_));
 sky130_fd_sc_hd__o221a_1 _4235_ (.A1(\game.counter[17] ),
    .A2(\game.counter[18] ),
    .B1(\game.counter[20] ),
    .B2(_0240_),
    .C1(_1501_),
    .X(_1502_));
 sky130_fd_sc_hd__a22o_1 _4236_ (.A1(\game.counter[21] ),
    .A2(_0241_),
    .B1(_0243_),
    .B2(\game.counter[14] ),
    .X(_1503_));
 sky130_fd_sc_hd__a211oi_1 _4237_ (.A1(\game.counter[9] ),
    .A2(_0245_),
    .B1(_1503_),
    .C1(_0236_),
    .Y(_1504_));
 sky130_fd_sc_hd__and2b_1 _4238_ (.A_N(_0249_),
    .B(_0223_),
    .X(_1505_));
 sky130_fd_sc_hd__o2111a_1 _4239_ (.A1(\game.counter[15] ),
    .A2(_0222_),
    .B1(_0229_),
    .C1(_0230_),
    .D1(_1505_),
    .X(_1506_));
 sky130_fd_sc_hd__o2111a_1 _4240_ (.A1(\game.counter[16] ),
    .A2(_0245_),
    .B1(_1502_),
    .C1(_1504_),
    .D1(_1506_),
    .X(_1507_));
 sky130_fd_sc_hd__and4_1 _4241_ (.A(_0228_),
    .B(_1496_),
    .C(_1500_),
    .D(_1507_),
    .X(_1508_));
 sky130_fd_sc_hd__a22o_1 _4242_ (.A1(_1405_),
    .A2(_1495_),
    .B1(_1508_),
    .B2(net135),
    .X(\game.scoring_button_2.next_start_count ));
 sky130_fd_sc_hd__and2b_1 _4243_ (.A_N(\game.scoring_button_2.flash_counter_2[0] ),
    .B(_1486_),
    .X(_1509_));
 sky130_fd_sc_hd__clkbuf_1 _4244_ (.A(_1509_),
    .X(\game.scoring_button_2.next_flash_counter_2[0] ));
 sky130_fd_sc_hd__o21ai_1 _4245_ (.A1(net107),
    .A2(\game.scoring_button_2.flash_counter_2[0] ),
    .B1(\game.missed_2 ),
    .Y(_1510_));
 sky130_fd_sc_hd__a21oi_1 _4246_ (.A1(net107),
    .A2(\game.scoring_button_2.flash_counter_2[0] ),
    .B1(_1510_),
    .Y(\game.scoring_button_2.next_flash_counter_2[1] ));
 sky130_fd_sc_hd__and3_1 _4247_ (.A(\game.scoring_button_2.flash_counter_2[1] ),
    .B(\game.scoring_button_2.flash_counter_2[0] ),
    .C(\game.scoring_button_2.flash_counter_2[2] ),
    .X(_1511_));
 sky130_fd_sc_hd__a21o_1 _4248_ (.A1(\game.scoring_button_2.flash_counter_2[1] ),
    .A2(\game.scoring_button_2.flash_counter_2[0] ),
    .B1(\game.scoring_button_2.flash_counter_2[2] ),
    .X(_1512_));
 sky130_fd_sc_hd__and3b_1 _4249_ (.A_N(_1511_),
    .B(\game.missed_2 ),
    .C(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__clkbuf_1 _4250_ (.A(_1513_),
    .X(\game.scoring_button_2.next_flash_counter_2[2] ));
 sky130_fd_sc_hd__and2_1 _4251_ (.A(\game.scoring_button_2.flash_counter_2[3] ),
    .B(_1511_),
    .X(_1514_));
 sky130_fd_sc_hd__or2_1 _4252_ (.A(\game.scoring_button_2.flash_counter_2[3] ),
    .B(_1511_),
    .X(_1515_));
 sky130_fd_sc_hd__and3b_1 _4253_ (.A_N(_1514_),
    .B(\game.missed_2 ),
    .C(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__clkbuf_1 _4254_ (.A(_1516_),
    .X(\game.scoring_button_2.next_flash_counter_2[3] ));
 sky130_fd_sc_hd__a21boi_1 _4255_ (.A1(\game.scoring_button_2.flash_counter_2[4] ),
    .A2(_1514_),
    .B1_N(\game.missed_2 ),
    .Y(_1517_));
 sky130_fd_sc_hd__o21a_1 _4256_ (.A1(net201),
    .A2(_1514_),
    .B1(_1517_),
    .X(\game.scoring_button_2.next_flash_counter_2[4] ));
 sky130_fd_sc_hd__and3_1 _4257_ (.A(\game.scoring_button_2.flash_counter_2[5] ),
    .B(\game.scoring_button_2.flash_counter_2[4] ),
    .C(_1514_),
    .X(_1518_));
 sky130_fd_sc_hd__a31o_1 _4258_ (.A1(\game.scoring_button_2.flash_counter_2[3] ),
    .A2(\game.scoring_button_2.flash_counter_2[4] ),
    .A3(_1511_),
    .B1(\game.scoring_button_2.flash_counter_2[5] ),
    .X(_1519_));
 sky130_fd_sc_hd__and3b_1 _4259_ (.A_N(_1518_),
    .B(\game.missed_2 ),
    .C(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__clkbuf_1 _4260_ (.A(_1520_),
    .X(\game.scoring_button_2.next_flash_counter_2[5] ));
 sky130_fd_sc_hd__and2_1 _4261_ (.A(\game.scoring_button_2.flash_counter_2[6] ),
    .B(_1518_),
    .X(_1521_));
 sky130_fd_sc_hd__or2_1 _4262_ (.A(\game.scoring_button_2.flash_counter_2[6] ),
    .B(_1518_),
    .X(_1522_));
 sky130_fd_sc_hd__and3b_1 _4263_ (.A_N(_1521_),
    .B(_1486_),
    .C(_1522_),
    .X(_1523_));
 sky130_fd_sc_hd__clkbuf_1 _4264_ (.A(_1523_),
    .X(\game.scoring_button_2.next_flash_counter_2[6] ));
 sky130_fd_sc_hd__a21boi_1 _4265_ (.A1(net151),
    .A2(_1521_),
    .B1_N(\game.missed_2 ),
    .Y(_1524_));
 sky130_fd_sc_hd__o21a_1 _4266_ (.A1(net151),
    .A2(_1521_),
    .B1(_1524_),
    .X(\game.scoring_button_2.next_flash_counter_2[7] ));
 sky130_fd_sc_hd__and3_1 _4267_ (.A(\game.scoring_button_2.flash_counter_2[7] ),
    .B(\game.scoring_button_2.flash_counter_2[8] ),
    .C(_1521_),
    .X(_1525_));
 sky130_fd_sc_hd__a31o_1 _4268_ (.A1(\game.scoring_button_2.flash_counter_2[7] ),
    .A2(\game.scoring_button_2.flash_counter_2[6] ),
    .A3(_1518_),
    .B1(\game.scoring_button_2.flash_counter_2[8] ),
    .X(_1526_));
 sky130_fd_sc_hd__and3b_1 _4269_ (.A_N(_1525_),
    .B(\game.missed_2 ),
    .C(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__clkbuf_1 _4270_ (.A(_1527_),
    .X(\game.scoring_button_2.next_flash_counter_2[8] ));
 sky130_fd_sc_hd__and2_1 _4271_ (.A(\game.scoring_button_2.flash_counter_2[9] ),
    .B(_1525_),
    .X(_1528_));
 sky130_fd_sc_hd__or2_1 _4272_ (.A(\game.scoring_button_2.flash_counter_2[9] ),
    .B(_1525_),
    .X(_1529_));
 sky130_fd_sc_hd__and3b_1 _4273_ (.A_N(_1528_),
    .B(_1486_),
    .C(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__clkbuf_1 _4274_ (.A(_1530_),
    .X(\game.scoring_button_2.next_flash_counter_2[9] ));
 sky130_fd_sc_hd__a21boi_1 _4275_ (.A1(net166),
    .A2(_1528_),
    .B1_N(\game.missed_2 ),
    .Y(_1531_));
 sky130_fd_sc_hd__o21a_1 _4276_ (.A1(net166),
    .A2(_1528_),
    .B1(_1531_),
    .X(\game.scoring_button_2.next_flash_counter_2[10] ));
 sky130_fd_sc_hd__and3_1 _4277_ (.A(\game.scoring_button_2.flash_counter_2[11] ),
    .B(\game.scoring_button_2.flash_counter_2[10] ),
    .C(_1528_),
    .X(_1532_));
 sky130_fd_sc_hd__a31o_1 _4278_ (.A1(\game.scoring_button_2.flash_counter_2[9] ),
    .A2(\game.scoring_button_2.flash_counter_2[10] ),
    .A3(_1525_),
    .B1(\game.scoring_button_2.flash_counter_2[11] ),
    .X(_1533_));
 sky130_fd_sc_hd__and3b_1 _4279_ (.A_N(_1532_),
    .B(\game.missed_2 ),
    .C(_1533_),
    .X(_1534_));
 sky130_fd_sc_hd__clkbuf_1 _4280_ (.A(_1534_),
    .X(\game.scoring_button_2.next_flash_counter_2[11] ));
 sky130_fd_sc_hd__and2_1 _4281_ (.A(\game.scoring_button_2.flash_counter_2[12] ),
    .B(_1532_),
    .X(_1535_));
 sky130_fd_sc_hd__or2_1 _4282_ (.A(\game.scoring_button_2.flash_counter_2[12] ),
    .B(_1532_),
    .X(_1536_));
 sky130_fd_sc_hd__and3b_1 _4283_ (.A_N(_1535_),
    .B(\game.missed_2 ),
    .C(_1536_),
    .X(_1537_));
 sky130_fd_sc_hd__clkbuf_1 _4284_ (.A(_1537_),
    .X(\game.scoring_button_2.next_flash_counter_2[12] ));
 sky130_fd_sc_hd__a21boi_1 _4285_ (.A1(net159),
    .A2(_1535_),
    .B1_N(\game.missed_2 ),
    .Y(_1538_));
 sky130_fd_sc_hd__o21a_1 _4286_ (.A1(net159),
    .A2(_1535_),
    .B1(_1538_),
    .X(\game.scoring_button_2.next_flash_counter_2[13] ));
 sky130_fd_sc_hd__and3_1 _4287_ (.A(\game.scoring_button_2.flash_counter_2[13] ),
    .B(\game.scoring_button_2.flash_counter_2[14] ),
    .C(_1535_),
    .X(_1539_));
 sky130_fd_sc_hd__a31o_1 _4288_ (.A1(\game.scoring_button_2.flash_counter_2[13] ),
    .A2(\game.scoring_button_2.flash_counter_2[12] ),
    .A3(_1532_),
    .B1(\game.scoring_button_2.flash_counter_2[14] ),
    .X(_1540_));
 sky130_fd_sc_hd__and3b_1 _4289_ (.A_N(_1539_),
    .B(_1486_),
    .C(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__clkbuf_1 _4290_ (.A(_1541_),
    .X(\game.scoring_button_2.next_flash_counter_2[14] ));
 sky130_fd_sc_hd__and2_1 _4291_ (.A(\game.scoring_button_2.flash_counter_2[15] ),
    .B(_1539_),
    .X(_1542_));
 sky130_fd_sc_hd__or2_1 _4292_ (.A(\game.scoring_button_2.flash_counter_2[15] ),
    .B(_1539_),
    .X(_1543_));
 sky130_fd_sc_hd__and3b_1 _4293_ (.A_N(_1542_),
    .B(\game.missed_2 ),
    .C(_1543_),
    .X(_1544_));
 sky130_fd_sc_hd__clkbuf_1 _4294_ (.A(_1544_),
    .X(\game.scoring_button_2.next_flash_counter_2[15] ));
 sky130_fd_sc_hd__a21boi_1 _4295_ (.A1(\game.scoring_button_2.flash_counter_2[16] ),
    .A2(_1542_),
    .B1_N(_1486_),
    .Y(_1545_));
 sky130_fd_sc_hd__o21a_1 _4296_ (.A1(net185),
    .A2(_1542_),
    .B1(_1545_),
    .X(\game.scoring_button_2.next_flash_counter_2[16] ));
 sky130_fd_sc_hd__and3_1 _4297_ (.A(\game.scoring_button_2.flash_counter_2[17] ),
    .B(\game.scoring_button_2.flash_counter_2[16] ),
    .C(_1542_),
    .X(_1546_));
 sky130_fd_sc_hd__a31o_1 _4298_ (.A1(\game.scoring_button_2.flash_counter_2[15] ),
    .A2(\game.scoring_button_2.flash_counter_2[16] ),
    .A3(_1539_),
    .B1(\game.scoring_button_2.flash_counter_2[17] ),
    .X(_1547_));
 sky130_fd_sc_hd__and3b_1 _4299_ (.A_N(_1546_),
    .B(_1486_),
    .C(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__clkbuf_1 _4300_ (.A(_1548_),
    .X(\game.scoring_button_2.next_flash_counter_2[17] ));
 sky130_fd_sc_hd__and2_1 _4301_ (.A(\game.scoring_button_2.flash_counter_2[18] ),
    .B(_1546_),
    .X(_1549_));
 sky130_fd_sc_hd__or2_1 _4302_ (.A(\game.scoring_button_2.flash_counter_2[18] ),
    .B(_1546_),
    .X(_1550_));
 sky130_fd_sc_hd__and3b_1 _4303_ (.A_N(_1549_),
    .B(_1486_),
    .C(_1550_),
    .X(_1551_));
 sky130_fd_sc_hd__clkbuf_1 _4304_ (.A(_1551_),
    .X(\game.scoring_button_2.next_flash_counter_2[18] ));
 sky130_fd_sc_hd__a21boi_1 _4305_ (.A1(net169),
    .A2(_1549_),
    .B1_N(_1486_),
    .Y(_1552_));
 sky130_fd_sc_hd__o21a_1 _4306_ (.A1(net169),
    .A2(_1549_),
    .B1(_1552_),
    .X(\game.scoring_button_2.next_flash_counter_2[19] ));
 sky130_fd_sc_hd__and3_1 _4307_ (.A(\game.scoring_button_2.flash_counter_2[19] ),
    .B(\game.scoring_button_2.flash_counter_2[20] ),
    .C(_1549_),
    .X(_1553_));
 sky130_fd_sc_hd__a31o_1 _4308_ (.A1(\game.scoring_button_2.flash_counter_2[19] ),
    .A2(\game.scoring_button_2.flash_counter_2[18] ),
    .A3(_1546_),
    .B1(\game.scoring_button_2.flash_counter_2[20] ),
    .X(_1554_));
 sky130_fd_sc_hd__and3b_1 _4309_ (.A_N(_1553_),
    .B(\game.missed_2 ),
    .C(_1554_),
    .X(_1555_));
 sky130_fd_sc_hd__clkbuf_1 _4310_ (.A(_1555_),
    .X(\game.scoring_button_2.next_flash_counter_2[20] ));
 sky130_fd_sc_hd__and2_1 _4311_ (.A(\game.scoring_button_2.flash_counter_2[21] ),
    .B(_1553_),
    .X(_1556_));
 sky130_fd_sc_hd__or2_1 _4312_ (.A(\game.scoring_button_2.flash_counter_2[21] ),
    .B(_1553_),
    .X(_1557_));
 sky130_fd_sc_hd__and3b_1 _4313_ (.A_N(_1556_),
    .B(\game.missed_2 ),
    .C(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__clkbuf_1 _4314_ (.A(_1558_),
    .X(\game.scoring_button_2.next_flash_counter_2[21] ));
 sky130_fd_sc_hd__o21ai_1 _4315_ (.A1(net87),
    .A2(_1556_),
    .B1(\game.missed_2 ),
    .Y(_1559_));
 sky130_fd_sc_hd__a21oi_1 _4316_ (.A1(net87),
    .A2(_1556_),
    .B1(_1559_),
    .Y(\game.scoring_button_2.next_flash_counter_2[22] ));
 sky130_fd_sc_hd__and2b_1 _4317_ (.A_N(\game.scoring_button_2.flash_counter_1[0] ),
    .B(_1413_),
    .X(_1560_));
 sky130_fd_sc_hd__clkbuf_1 _4318_ (.A(_1560_),
    .X(\game.scoring_button_2.next_flash_counter_1[0] ));
 sky130_fd_sc_hd__o21ai_1 _4319_ (.A1(net103),
    .A2(\game.scoring_button_2.flash_counter_1[0] ),
    .B1(\game.hit_2 ),
    .Y(_1561_));
 sky130_fd_sc_hd__a21oi_1 _4320_ (.A1(net103),
    .A2(\game.scoring_button_2.flash_counter_1[0] ),
    .B1(_1561_),
    .Y(\game.scoring_button_2.next_flash_counter_1[1] ));
 sky130_fd_sc_hd__and3_1 _4321_ (.A(\game.scoring_button_2.flash_counter_1[1] ),
    .B(\game.scoring_button_2.flash_counter_1[0] ),
    .C(\game.scoring_button_2.flash_counter_1[2] ),
    .X(_1562_));
 sky130_fd_sc_hd__a21o_1 _4322_ (.A1(\game.scoring_button_2.flash_counter_1[1] ),
    .A2(\game.scoring_button_2.flash_counter_1[0] ),
    .B1(\game.scoring_button_2.flash_counter_1[2] ),
    .X(_1563_));
 sky130_fd_sc_hd__and3b_1 _4323_ (.A_N(_1562_),
    .B(\game.hit_2 ),
    .C(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__clkbuf_1 _4324_ (.A(_1564_),
    .X(\game.scoring_button_2.next_flash_counter_1[2] ));
 sky130_fd_sc_hd__and2_1 _4325_ (.A(\game.scoring_button_2.flash_counter_1[3] ),
    .B(_1562_),
    .X(_1565_));
 sky130_fd_sc_hd__or2_1 _4326_ (.A(\game.scoring_button_2.flash_counter_1[3] ),
    .B(_1562_),
    .X(_1566_));
 sky130_fd_sc_hd__and3b_1 _4327_ (.A_N(_1565_),
    .B(\game.hit_2 ),
    .C(_1566_),
    .X(_1567_));
 sky130_fd_sc_hd__clkbuf_1 _4328_ (.A(_1567_),
    .X(\game.scoring_button_2.next_flash_counter_1[3] ));
 sky130_fd_sc_hd__a21boi_1 _4329_ (.A1(net176),
    .A2(_1565_),
    .B1_N(\game.hit_2 ),
    .Y(_1568_));
 sky130_fd_sc_hd__o21a_1 _4330_ (.A1(net176),
    .A2(_1565_),
    .B1(_1568_),
    .X(\game.scoring_button_2.next_flash_counter_1[4] ));
 sky130_fd_sc_hd__and3_1 _4331_ (.A(\game.scoring_button_2.flash_counter_1[5] ),
    .B(\game.scoring_button_2.flash_counter_1[4] ),
    .C(_1565_),
    .X(_1569_));
 sky130_fd_sc_hd__a31o_1 _4332_ (.A1(\game.scoring_button_2.flash_counter_1[3] ),
    .A2(\game.scoring_button_2.flash_counter_1[4] ),
    .A3(_1562_),
    .B1(\game.scoring_button_2.flash_counter_1[5] ),
    .X(_1570_));
 sky130_fd_sc_hd__and3b_1 _4333_ (.A_N(_1569_),
    .B(\game.hit_2 ),
    .C(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__clkbuf_1 _4334_ (.A(_1571_),
    .X(\game.scoring_button_2.next_flash_counter_1[5] ));
 sky130_fd_sc_hd__and2_1 _4335_ (.A(\game.scoring_button_2.flash_counter_1[6] ),
    .B(_1569_),
    .X(_1572_));
 sky130_fd_sc_hd__or2_1 _4336_ (.A(\game.scoring_button_2.flash_counter_1[6] ),
    .B(_1569_),
    .X(_1573_));
 sky130_fd_sc_hd__and3b_1 _4337_ (.A_N(_1572_),
    .B(_1413_),
    .C(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__clkbuf_1 _4338_ (.A(_1574_),
    .X(\game.scoring_button_2.next_flash_counter_1[6] ));
 sky130_fd_sc_hd__a21boi_1 _4339_ (.A1(\game.scoring_button_2.flash_counter_1[7] ),
    .A2(_1572_),
    .B1_N(\game.hit_2 ),
    .Y(_1575_));
 sky130_fd_sc_hd__o21a_1 _4340_ (.A1(net192),
    .A2(_1572_),
    .B1(_1575_),
    .X(\game.scoring_button_2.next_flash_counter_1[7] ));
 sky130_fd_sc_hd__and3_1 _4341_ (.A(\game.scoring_button_2.flash_counter_1[7] ),
    .B(\game.scoring_button_2.flash_counter_1[8] ),
    .C(_1572_),
    .X(_1576_));
 sky130_fd_sc_hd__a31o_1 _4342_ (.A1(\game.scoring_button_2.flash_counter_1[7] ),
    .A2(\game.scoring_button_2.flash_counter_1[6] ),
    .A3(_1569_),
    .B1(\game.scoring_button_2.flash_counter_1[8] ),
    .X(_1577_));
 sky130_fd_sc_hd__and3b_1 _4343_ (.A_N(_1576_),
    .B(\game.hit_2 ),
    .C(_1577_),
    .X(_1578_));
 sky130_fd_sc_hd__clkbuf_1 _4344_ (.A(_1578_),
    .X(\game.scoring_button_2.next_flash_counter_1[8] ));
 sky130_fd_sc_hd__and2_1 _4345_ (.A(\game.scoring_button_2.flash_counter_1[9] ),
    .B(_1576_),
    .X(_1579_));
 sky130_fd_sc_hd__or2_1 _4346_ (.A(\game.scoring_button_2.flash_counter_1[9] ),
    .B(_1576_),
    .X(_1580_));
 sky130_fd_sc_hd__and3b_1 _4347_ (.A_N(_1579_),
    .B(_1413_),
    .C(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__clkbuf_1 _4348_ (.A(_1581_),
    .X(\game.scoring_button_2.next_flash_counter_1[9] ));
 sky130_fd_sc_hd__a21boi_1 _4349_ (.A1(net156),
    .A2(_1579_),
    .B1_N(\game.hit_2 ),
    .Y(_1582_));
 sky130_fd_sc_hd__o21a_1 _4350_ (.A1(net156),
    .A2(_1579_),
    .B1(_1582_),
    .X(\game.scoring_button_2.next_flash_counter_1[10] ));
 sky130_fd_sc_hd__and3_1 _4351_ (.A(\game.scoring_button_2.flash_counter_1[11] ),
    .B(\game.scoring_button_2.flash_counter_1[10] ),
    .C(_1579_),
    .X(_1583_));
 sky130_fd_sc_hd__a31o_1 _4352_ (.A1(\game.scoring_button_2.flash_counter_1[9] ),
    .A2(\game.scoring_button_2.flash_counter_1[10] ),
    .A3(_1576_),
    .B1(\game.scoring_button_2.flash_counter_1[11] ),
    .X(_1584_));
 sky130_fd_sc_hd__and3b_1 _4353_ (.A_N(_1583_),
    .B(\game.hit_2 ),
    .C(_1584_),
    .X(_1585_));
 sky130_fd_sc_hd__clkbuf_1 _4354_ (.A(_1585_),
    .X(\game.scoring_button_2.next_flash_counter_1[11] ));
 sky130_fd_sc_hd__and2_1 _4355_ (.A(\game.scoring_button_2.flash_counter_1[12] ),
    .B(_1583_),
    .X(_1586_));
 sky130_fd_sc_hd__or2_1 _4356_ (.A(\game.scoring_button_2.flash_counter_1[12] ),
    .B(_1583_),
    .X(_1587_));
 sky130_fd_sc_hd__and3b_1 _4357_ (.A_N(_1586_),
    .B(\game.hit_2 ),
    .C(_1587_),
    .X(_1588_));
 sky130_fd_sc_hd__clkbuf_1 _4358_ (.A(_1588_),
    .X(\game.scoring_button_2.next_flash_counter_1[12] ));
 sky130_fd_sc_hd__a21boi_1 _4359_ (.A1(net173),
    .A2(_1586_),
    .B1_N(\game.hit_2 ),
    .Y(_1589_));
 sky130_fd_sc_hd__o21a_1 _4360_ (.A1(net173),
    .A2(_1586_),
    .B1(_1589_),
    .X(\game.scoring_button_2.next_flash_counter_1[13] ));
 sky130_fd_sc_hd__and3_1 _4361_ (.A(\game.scoring_button_2.flash_counter_1[13] ),
    .B(\game.scoring_button_2.flash_counter_1[14] ),
    .C(_1586_),
    .X(_1590_));
 sky130_fd_sc_hd__a31o_1 _4362_ (.A1(\game.scoring_button_2.flash_counter_1[13] ),
    .A2(\game.scoring_button_2.flash_counter_1[12] ),
    .A3(_1583_),
    .B1(\game.scoring_button_2.flash_counter_1[14] ),
    .X(_1591_));
 sky130_fd_sc_hd__and3b_1 _4363_ (.A_N(_1590_),
    .B(_1413_),
    .C(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__clkbuf_1 _4364_ (.A(_1592_),
    .X(\game.scoring_button_2.next_flash_counter_1[14] ));
 sky130_fd_sc_hd__and2_1 _4365_ (.A(\game.scoring_button_2.flash_counter_1[15] ),
    .B(_1590_),
    .X(_1593_));
 sky130_fd_sc_hd__or2_1 _4366_ (.A(\game.scoring_button_2.flash_counter_1[15] ),
    .B(_1590_),
    .X(_1594_));
 sky130_fd_sc_hd__and3b_1 _4367_ (.A_N(_1593_),
    .B(\game.hit_2 ),
    .C(_1594_),
    .X(_1595_));
 sky130_fd_sc_hd__clkbuf_1 _4368_ (.A(_1595_),
    .X(\game.scoring_button_2.next_flash_counter_1[15] ));
 sky130_fd_sc_hd__a21boi_1 _4369_ (.A1(net174),
    .A2(_1593_),
    .B1_N(_1413_),
    .Y(_1596_));
 sky130_fd_sc_hd__o21a_1 _4370_ (.A1(net174),
    .A2(_1593_),
    .B1(_1596_),
    .X(\game.scoring_button_2.next_flash_counter_1[16] ));
 sky130_fd_sc_hd__and3_1 _4371_ (.A(\game.scoring_button_2.flash_counter_1[17] ),
    .B(\game.scoring_button_2.flash_counter_1[16] ),
    .C(_1593_),
    .X(_1597_));
 sky130_fd_sc_hd__a31o_1 _4372_ (.A1(\game.scoring_button_2.flash_counter_1[15] ),
    .A2(\game.scoring_button_2.flash_counter_1[16] ),
    .A3(_1590_),
    .B1(\game.scoring_button_2.flash_counter_1[17] ),
    .X(_1598_));
 sky130_fd_sc_hd__and3b_1 _4373_ (.A_N(_1597_),
    .B(_1413_),
    .C(_1598_),
    .X(_1599_));
 sky130_fd_sc_hd__clkbuf_1 _4374_ (.A(_1599_),
    .X(\game.scoring_button_2.next_flash_counter_1[17] ));
 sky130_fd_sc_hd__and2_1 _4375_ (.A(\game.scoring_button_2.flash_counter_1[18] ),
    .B(_1597_),
    .X(_1600_));
 sky130_fd_sc_hd__or2_1 _4376_ (.A(\game.scoring_button_2.flash_counter_1[18] ),
    .B(_1597_),
    .X(_1601_));
 sky130_fd_sc_hd__and3b_1 _4377_ (.A_N(_1600_),
    .B(_1413_),
    .C(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__clkbuf_1 _4378_ (.A(_1602_),
    .X(\game.scoring_button_2.next_flash_counter_1[18] ));
 sky130_fd_sc_hd__a21boi_1 _4379_ (.A1(net171),
    .A2(_1600_),
    .B1_N(_1413_),
    .Y(_1603_));
 sky130_fd_sc_hd__o21a_1 _4380_ (.A1(net171),
    .A2(_1600_),
    .B1(_1603_),
    .X(\game.scoring_button_2.next_flash_counter_1[19] ));
 sky130_fd_sc_hd__and3_1 _4381_ (.A(\game.scoring_button_2.flash_counter_1[19] ),
    .B(\game.scoring_button_2.flash_counter_1[20] ),
    .C(_1600_),
    .X(_1604_));
 sky130_fd_sc_hd__a31o_1 _4382_ (.A1(\game.scoring_button_2.flash_counter_1[19] ),
    .A2(\game.scoring_button_2.flash_counter_1[18] ),
    .A3(_1597_),
    .B1(\game.scoring_button_2.flash_counter_1[20] ),
    .X(_1605_));
 sky130_fd_sc_hd__and3b_1 _4383_ (.A_N(_1604_),
    .B(\game.hit_2 ),
    .C(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__clkbuf_1 _4384_ (.A(_1606_),
    .X(\game.scoring_button_2.next_flash_counter_1[20] ));
 sky130_fd_sc_hd__and2_1 _4385_ (.A(\game.scoring_button_2.flash_counter_1[21] ),
    .B(_1604_),
    .X(_1607_));
 sky130_fd_sc_hd__or2_1 _4386_ (.A(\game.scoring_button_2.flash_counter_1[21] ),
    .B(_1604_),
    .X(_1608_));
 sky130_fd_sc_hd__and3b_1 _4387_ (.A_N(_1607_),
    .B(\game.hit_2 ),
    .C(_1608_),
    .X(_1609_));
 sky130_fd_sc_hd__clkbuf_1 _4388_ (.A(_1609_),
    .X(\game.scoring_button_2.next_flash_counter_1[21] ));
 sky130_fd_sc_hd__o21ai_1 _4389_ (.A1(net89),
    .A2(_1607_),
    .B1(\game.hit_2 ),
    .Y(_1610_));
 sky130_fd_sc_hd__a21oi_1 _4390_ (.A1(net89),
    .A2(_1607_),
    .B1(_1610_),
    .Y(\game.scoring_button_2.next_flash_counter_1[22] ));
 sky130_fd_sc_hd__and3b_1 _4391_ (.A_N(\game.scoring_button_1.check_hit.edge_1 ),
    .B(\game.scoring_button_1.check_hit.edge_2 ),
    .C(\game.scoring_button_1.hit ),
    .X(_1611_));
 sky130_fd_sc_hd__buf_6 _4392_ (.A(_1611_),
    .X(_1612_));
 sky130_fd_sc_hd__nor2_8 _4393_ (.A(_0208_),
    .B(_1612_),
    .Y(_1613_));
 sky130_fd_sc_hd__mux2_1 _4394_ (.A0(_1612_),
    .A1(_1613_),
    .S(\game.addhits.a[0] ),
    .X(_1614_));
 sky130_fd_sc_hd__clkbuf_1 _4395_ (.A(_1614_),
    .X(\game.scoring_button_1.next_num_hits[0] ));
 sky130_fd_sc_hd__nor2_1 _4396_ (.A(\game.addhits.a[2] ),
    .B(\game.scoring_button_1.acc[2] ),
    .Y(_1615_));
 sky130_fd_sc_hd__or2_1 _4397_ (.A(\game.addhits.a[1] ),
    .B(\game.scoring_button_1.acc[1] ),
    .X(_1616_));
 sky130_fd_sc_hd__nand2_1 _4398_ (.A(\game.addhits.a[1] ),
    .B(\game.scoring_button_1.acc[1] ),
    .Y(_1617_));
 sky130_fd_sc_hd__a21boi_1 _4399_ (.A1(\game.addhits.a[0] ),
    .A2(_1616_),
    .B1_N(_1617_),
    .Y(_1618_));
 sky130_fd_sc_hd__nand2_1 _4400_ (.A(\game.addhits.a[2] ),
    .B(\game.scoring_button_1.acc[2] ),
    .Y(_1619_));
 sky130_fd_sc_hd__o21ai_1 _4401_ (.A1(_1615_),
    .A2(_1618_),
    .B1(_1619_),
    .Y(_1620_));
 sky130_fd_sc_hd__nor2_1 _4402_ (.A(\game.addhits.a[3] ),
    .B(_1620_),
    .Y(_1621_));
 sky130_fd_sc_hd__nand2_1 _4403_ (.A(_1617_),
    .B(_1616_),
    .Y(_1622_));
 sky130_fd_sc_hd__xor2_1 _4404_ (.A(\game.addhits.a[0] ),
    .B(_1622_),
    .X(_1623_));
 sky130_fd_sc_hd__or2_1 _4405_ (.A(\game.addhits.a[2] ),
    .B(\game.scoring_button_1.acc[2] ),
    .X(_1624_));
 sky130_fd_sc_hd__nand2_1 _4406_ (.A(_1619_),
    .B(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__xnor2_1 _4407_ (.A(_1618_),
    .B(_1625_),
    .Y(_1626_));
 sky130_fd_sc_hd__nand2_1 _4408_ (.A(_1623_),
    .B(_1626_),
    .Y(_1627_));
 sky130_fd_sc_hd__inv_2 _4409_ (.A(_1627_),
    .Y(_1628_));
 sky130_fd_sc_hd__nand2_1 _4410_ (.A(\game.addhits.a[3] ),
    .B(_1620_),
    .Y(_1629_));
 sky130_fd_sc_hd__o21ai_2 _4411_ (.A1(_1621_),
    .A2(_1628_),
    .B1(_1629_),
    .Y(_1630_));
 sky130_fd_sc_hd__mux2_1 _4412_ (.A0(_1621_),
    .A1(_1630_),
    .S(_1623_),
    .X(_1631_));
 sky130_fd_sc_hd__a22o_1 _4413_ (.A1(\game.addhits.a[1] ),
    .A2(_1613_),
    .B1(_1631_),
    .B2(_1612_),
    .X(\game.scoring_button_1.next_num_hits[1] ));
 sky130_fd_sc_hd__or2_1 _4414_ (.A(_1629_),
    .B(_1627_),
    .X(_1632_));
 sky130_fd_sc_hd__a21o_1 _4415_ (.A1(_1623_),
    .A2(_1630_),
    .B1(_1626_),
    .X(_1633_));
 sky130_fd_sc_hd__nand2_1 _4416_ (.A(_1632_),
    .B(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__a22o_1 _4417_ (.A1(net208),
    .A2(_1613_),
    .B1(_1634_),
    .B2(_1612_),
    .X(\game.scoring_button_1.next_num_hits[2] ));
 sky130_fd_sc_hd__o21ai_1 _4418_ (.A1(_1621_),
    .A2(_1627_),
    .B1(_1629_),
    .Y(_1635_));
 sky130_fd_sc_hd__a32o_1 _4419_ (.A1(_1612_),
    .A2(_1632_),
    .A3(_1635_),
    .B1(_1613_),
    .B2(net202),
    .X(\game.scoring_button_1.next_num_hits[3] ));
 sky130_fd_sc_hd__or2_1 _4420_ (.A(\game.addhits.a[4] ),
    .B(_1630_),
    .X(_1636_));
 sky130_fd_sc_hd__and2_1 _4421_ (.A(\game.addhits.a[4] ),
    .B(_1630_),
    .X(_1637_));
 sky130_fd_sc_hd__inv_2 _4422_ (.A(_1637_),
    .Y(_1638_));
 sky130_fd_sc_hd__a32o_1 _4423_ (.A1(_1612_),
    .A2(_1636_),
    .A3(_1638_),
    .B1(_1613_),
    .B2(net267),
    .X(\game.scoring_button_1.next_num_hits[4] ));
 sky130_fd_sc_hd__o31a_2 _4424_ (.A1(\game.addhits.a[6] ),
    .A2(\game.addhits.a[5] ),
    .A3(_1637_),
    .B1(\game.addhits.a[7] ),
    .X(_1639_));
 sky130_fd_sc_hd__xnor2_1 _4425_ (.A(\game.addhits.a[5] ),
    .B(_1637_),
    .Y(_1640_));
 sky130_fd_sc_hd__xnor2_1 _4426_ (.A(_1639_),
    .B(_1640_),
    .Y(_1641_));
 sky130_fd_sc_hd__a22o_1 _4427_ (.A1(\game.addhits.a[5] ),
    .A2(_1613_),
    .B1(_1641_),
    .B2(_1612_),
    .X(\game.scoring_button_1.next_num_hits[5] ));
 sky130_fd_sc_hd__inv_2 _4428_ (.A(\game.addhits.a[6] ),
    .Y(_1642_));
 sky130_fd_sc_hd__inv_2 _4429_ (.A(\game.addhits.a[5] ),
    .Y(_1643_));
 sky130_fd_sc_hd__or3_1 _4430_ (.A(_1642_),
    .B(_1643_),
    .C(_1638_),
    .X(_1644_));
 sky130_fd_sc_hd__nor2_1 _4431_ (.A(\game.addhits.a[7] ),
    .B(_1644_),
    .Y(_1645_));
 sky130_fd_sc_hd__a31o_1 _4432_ (.A1(\game.addhits.a[5] ),
    .A2(\game.addhits.a[4] ),
    .A3(_1630_),
    .B1(\game.addhits.a[6] ),
    .X(_1646_));
 sky130_fd_sc_hd__nand2_1 _4433_ (.A(_1612_),
    .B(_1646_),
    .Y(_1647_));
 sky130_fd_sc_hd__a31o_1 _4434_ (.A1(_1639_),
    .A2(_1640_),
    .A3(_1644_),
    .B1(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__a2bb2o_1 _4435_ (.A1_N(_1645_),
    .A2_N(_1648_),
    .B1(net257),
    .B2(_1613_),
    .X(\game.scoring_button_1.next_num_hits[6] ));
 sky130_fd_sc_hd__a41o_1 _4436_ (.A1(_1642_),
    .A2(_1643_),
    .A3(_1612_),
    .A4(_1638_),
    .B1(_1613_),
    .X(_1649_));
 sky130_fd_sc_hd__a22o_1 _4437_ (.A1(_1612_),
    .A2(_1645_),
    .B1(_1649_),
    .B2(net220),
    .X(\game.scoring_button_1.next_num_hits[7] ));
 sky130_fd_sc_hd__and2_1 _4438_ (.A(\game.addhits.a[8] ),
    .B(_1639_),
    .X(_1650_));
 sky130_fd_sc_hd__o21ai_1 _4439_ (.A1(\game.addhits.a[8] ),
    .A2(_1639_),
    .B1(_1612_),
    .Y(_1651_));
 sky130_fd_sc_hd__a2bb2o_1 _4440_ (.A1_N(_1650_),
    .A2_N(_1651_),
    .B1(net216),
    .B2(_1613_),
    .X(\game.scoring_button_1.next_num_hits[8] ));
 sky130_fd_sc_hd__nor2_1 _4441_ (.A(\game.addhits.a[9] ),
    .B(_1650_),
    .Y(_1652_));
 sky130_fd_sc_hd__and3_1 _4442_ (.A(\game.addhits.a[9] ),
    .B(\game.addhits.a[8] ),
    .C(_1639_),
    .X(_1653_));
 sky130_fd_sc_hd__o31a_1 _4443_ (.A1(\game.addhits.a[10] ),
    .A2(\game.addhits.a[9] ),
    .A3(_1650_),
    .B1(\game.addhits.a[11] ),
    .X(_1654_));
 sky130_fd_sc_hd__o21ai_1 _4444_ (.A1(_1652_),
    .A2(_1653_),
    .B1(_1654_),
    .Y(_1655_));
 sky130_fd_sc_hd__o31ai_1 _4445_ (.A1(\game.addhits.a[11] ),
    .A2(_1652_),
    .A3(_1653_),
    .B1(_1655_),
    .Y(_1656_));
 sky130_fd_sc_hd__a22o_1 _4446_ (.A1(net260),
    .A2(_1613_),
    .B1(_1656_),
    .B2(_1612_),
    .X(\game.scoring_button_1.next_num_hits[9] ));
 sky130_fd_sc_hd__or2_1 _4447_ (.A(\game.addhits.a[10] ),
    .B(_1653_),
    .X(_1657_));
 sky130_fd_sc_hd__and2_1 _4448_ (.A(\game.addhits.a[10] ),
    .B(_1653_),
    .X(_1658_));
 sky130_fd_sc_hd__mux2_1 _4449_ (.A0(_1655_),
    .A1(\game.addhits.a[11] ),
    .S(_1658_),
    .X(_1659_));
 sky130_fd_sc_hd__a32o_1 _4450_ (.A1(_1612_),
    .A2(_1657_),
    .A3(_1659_),
    .B1(_1613_),
    .B2(net196),
    .X(\game.scoring_button_1.next_num_hits[10] ));
 sky130_fd_sc_hd__o21ba_1 _4451_ (.A1(\game.addhits.a[11] ),
    .A2(_1658_),
    .B1_N(_1654_),
    .X(_1660_));
 sky130_fd_sc_hd__a22o_1 _4452_ (.A1(net228),
    .A2(_1613_),
    .B1(_1660_),
    .B2(_1612_),
    .X(\game.scoring_button_1.next_num_hits[11] ));
 sky130_fd_sc_hd__and2_1 _4453_ (.A(\game.addhits.a[12] ),
    .B(_1654_),
    .X(_1661_));
 sky130_fd_sc_hd__o21ai_1 _4454_ (.A1(\game.addhits.a[12] ),
    .A2(_1654_),
    .B1(_1612_),
    .Y(_1662_));
 sky130_fd_sc_hd__a2bb2o_1 _4455_ (.A1_N(_1661_),
    .A2_N(_1662_),
    .B1(net189),
    .B2(_1613_),
    .X(\game.scoring_button_1.next_num_hits[12] ));
 sky130_fd_sc_hd__a21oi_1 _4456_ (.A1(\game.addhits.a[13] ),
    .A2(_1661_),
    .B1(\game.addhits.a[14] ),
    .Y(_1663_));
 sky130_fd_sc_hd__xnor2_1 _4457_ (.A(\game.addhits.a[13] ),
    .B(_1661_),
    .Y(_1664_));
 sky130_fd_sc_hd__nand2_1 _4458_ (.A(\game.addhits.a[15] ),
    .B(_1664_),
    .Y(_1665_));
 sky130_fd_sc_hd__or2_1 _4459_ (.A(\game.addhits.a[15] ),
    .B(_1664_),
    .X(_1666_));
 sky130_fd_sc_hd__o21ai_1 _4460_ (.A1(_1663_),
    .A2(_1665_),
    .B1(_1666_),
    .Y(_1667_));
 sky130_fd_sc_hd__a22o_1 _4461_ (.A1(net215),
    .A2(_1613_),
    .B1(_1667_),
    .B2(_1612_),
    .X(\game.scoring_button_1.next_num_hits[13] ));
 sky130_fd_sc_hd__and3_1 _4462_ (.A(\game.addhits.a[13] ),
    .B(\game.addhits.a[14] ),
    .C(_1661_),
    .X(_1668_));
 sky130_fd_sc_hd__a21oi_1 _4463_ (.A1(_0741_),
    .A2(_1668_),
    .B1(_1663_),
    .Y(_1669_));
 sky130_fd_sc_hd__or2_1 _4464_ (.A(_1665_),
    .B(_1668_),
    .X(_1670_));
 sky130_fd_sc_hd__a32o_1 _4465_ (.A1(_1612_),
    .A2(_1669_),
    .A3(_1670_),
    .B1(_1613_),
    .B2(net206),
    .X(\game.scoring_button_1.next_num_hits[14] ));
 sky130_fd_sc_hd__a21oi_1 _4466_ (.A1(\game.addhits.a[15] ),
    .A2(_1664_),
    .B1(_1668_),
    .Y(_1671_));
 sky130_fd_sc_hd__nor2_1 _4467_ (.A(_1669_),
    .B(_1671_),
    .Y(_1672_));
 sky130_fd_sc_hd__a22o_1 _4468_ (.A1(\game.addhits.a[15] ),
    .A2(_1613_),
    .B1(_1672_),
    .B2(_1612_),
    .X(\game.scoring_button_1.next_num_hits[15] ));
 sky130_fd_sc_hd__or2b_2 _4469_ (.A(\game.scoring_button_1.check_hit.edge_1 ),
    .B_N(\game.scoring_button_1.check_hit.edge_2 ),
    .X(_1673_));
 sky130_fd_sc_hd__or2_1 _4470_ (.A(\game.scoring_button_1.hit ),
    .B(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__clkbuf_8 _4471_ (.A(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__or3_1 _4472_ (.A(\game.scoring_button_1.counts[13] ),
    .B(\game.scoring_button_1.counts[12] ),
    .C(\game.scoring_button_1.counts[14] ),
    .X(_1676_));
 sky130_fd_sc_hd__or4_1 _4473_ (.A(\game.scoring_button_1.counts[19] ),
    .B(\game.scoring_button_1.counts[18] ),
    .C(\game.scoring_button_1.counts[17] ),
    .D(\game.scoring_button_1.counts[16] ),
    .X(_1677_));
 sky130_fd_sc_hd__or4_1 _4474_ (.A(\game.scoring_button_1.counts[22] ),
    .B(\game.scoring_button_1.counts[21] ),
    .C(\game.scoring_button_1.counts[20] ),
    .D(_1677_),
    .X(_1678_));
 sky130_fd_sc_hd__or4_1 _4475_ (.A(\game.scoring_button_1.counts[1] ),
    .B(\game.scoring_button_1.counts[3] ),
    .C(\game.scoring_button_1.counts[2] ),
    .D(\game.scoring_button_1.counts[4] ),
    .X(_1679_));
 sky130_fd_sc_hd__or4_1 _4476_ (.A(\game.scoring_button_1.counts[0] ),
    .B(\game.scoring_button_1.counts[6] ),
    .C(\game.scoring_button_1.counts[5] ),
    .D(_1679_),
    .X(_1680_));
 sky130_fd_sc_hd__or4_1 _4477_ (.A(\game.scoring_button_1.counts[10] ),
    .B(\game.scoring_button_1.counts[9] ),
    .C(\game.scoring_button_1.counts[8] ),
    .D(\game.scoring_button_1.counts[15] ),
    .X(_1681_));
 sky130_fd_sc_hd__or4_1 _4478_ (.A(\game.scoring_button_1.counts[7] ),
    .B(\game.scoring_button_1.counts[11] ),
    .C(_1680_),
    .D(_1681_),
    .X(_1682_));
 sky130_fd_sc_hd__a31o_1 _4479_ (.A1(\game.scoring_button_1.counts[7] ),
    .A2(\game.scoring_button_1.counts[8] ),
    .A3(_1680_),
    .B1(\game.scoring_button_1.counts[9] ),
    .X(_1683_));
 sky130_fd_sc_hd__a31o_1 _4480_ (.A1(\game.scoring_button_1.counts[11] ),
    .A2(\game.scoring_button_1.counts[10] ),
    .A3(_1683_),
    .B1(_1676_),
    .X(_1684_));
 sky130_fd_sc_hd__a41o_1 _4481_ (.A1(\game.scoring_button_1.counts[15] ),
    .A2(\game.scoring_button_1.counts[17] ),
    .A3(\game.scoring_button_1.counts[16] ),
    .A4(_1684_),
    .B1(\game.scoring_button_1.counts[18] ),
    .X(_1685_));
 sky130_fd_sc_hd__a31o_1 _4482_ (.A1(\game.scoring_button_1.counts[19] ),
    .A2(\game.scoring_button_1.counts[20] ),
    .A3(_1685_),
    .B1(\game.scoring_button_1.counts[21] ),
    .X(_1686_));
 sky130_fd_sc_hd__nand2_1 _4483_ (.A(\game.scoring_button_1.counts[22] ),
    .B(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hd__o31a_1 _4484_ (.A1(_1676_),
    .A2(_1678_),
    .A3(_1682_),
    .B1(_1687_),
    .X(_1688_));
 sky130_fd_sc_hd__nand2_2 _4485_ (.A(_0209_),
    .B(_2656_),
    .Y(_1689_));
 sky130_fd_sc_hd__or2_1 _4486_ (.A(_1688_),
    .B(_1689_),
    .X(_1690_));
 sky130_fd_sc_hd__clkbuf_4 _4487_ (.A(_1690_),
    .X(_1691_));
 sky130_fd_sc_hd__inv_2 _4488_ (.A(_1691_),
    .Y(_1692_));
 sky130_fd_sc_hd__nor2_2 _4489_ (.A(\modetrans.mode[0] ),
    .B(_1692_),
    .Y(_1693_));
 sky130_fd_sc_hd__a21oi_1 _4490_ (.A1(_1691_),
    .A2(_1675_),
    .B1(\game.addmisses.a[0] ),
    .Y(_1694_));
 sky130_fd_sc_hd__a31o_1 _4491_ (.A1(\game.addmisses.a[0] ),
    .A2(_1675_),
    .A3(_1693_),
    .B1(_1694_),
    .X(\game.scoring_button_1.next_num_misses[0] ));
 sky130_fd_sc_hd__xnor2_1 _4492_ (.A(\game.addmisses.a[1] ),
    .B(\game.addmisses.a[0] ),
    .Y(_1695_));
 sky130_fd_sc_hd__o2bb2a_1 _4493_ (.A1_N(\game.addmisses.a[1] ),
    .A2_N(_1693_),
    .B1(_1695_),
    .B2(_1691_),
    .X(_1696_));
 sky130_fd_sc_hd__o31a_1 _4494_ (.A1(\game.addmisses.a[2] ),
    .A2(\game.addmisses.a[1] ),
    .A3(\game.addmisses.a[0] ),
    .B1(\game.addmisses.a[3] ),
    .X(_1697_));
 sky130_fd_sc_hd__and2_1 _4495_ (.A(_1695_),
    .B(_1697_),
    .X(_1698_));
 sky130_fd_sc_hd__nor2_4 _4496_ (.A(\game.scoring_button_1.hit ),
    .B(_1673_),
    .Y(_1699_));
 sky130_fd_sc_hd__o21ai_1 _4497_ (.A1(\game.addmisses.a[3] ),
    .A2(_1695_),
    .B1(_1699_),
    .Y(_1700_));
 sky130_fd_sc_hd__o2bb2a_1 _4498_ (.A1_N(_1675_),
    .A2_N(_1696_),
    .B1(_1698_),
    .B2(_1700_),
    .X(\game.scoring_button_1.next_num_misses[1] ));
 sky130_fd_sc_hd__and3_1 _4499_ (.A(\game.addmisses.a[2] ),
    .B(\game.addmisses.a[1] ),
    .C(\game.addmisses.a[0] ),
    .X(_1701_));
 sky130_fd_sc_hd__a21oi_1 _4500_ (.A1(\game.addmisses.a[1] ),
    .A2(\game.addmisses.a[0] ),
    .B1(\game.addmisses.a[2] ),
    .Y(_1702_));
 sky130_fd_sc_hd__or2_1 _4501_ (.A(_1701_),
    .B(_1702_),
    .X(_1703_));
 sky130_fd_sc_hd__nor2_1 _4502_ (.A(_1698_),
    .B(_1703_),
    .Y(_1704_));
 sky130_fd_sc_hd__and2_1 _4503_ (.A(\game.addmisses.a[3] ),
    .B(_1701_),
    .X(_1705_));
 sky130_fd_sc_hd__nor2_1 _4504_ (.A(_1691_),
    .B(_1703_),
    .Y(_1706_));
 sky130_fd_sc_hd__a211o_1 _4505_ (.A1(\game.addmisses.a[2] ),
    .A2(_1693_),
    .B1(_1706_),
    .C1(_1699_),
    .X(_1707_));
 sky130_fd_sc_hd__o31a_1 _4506_ (.A1(_1675_),
    .A2(_1704_),
    .A3(_1705_),
    .B1(_1707_),
    .X(\game.scoring_button_1.next_num_misses[2] ));
 sky130_fd_sc_hd__nor2_1 _4507_ (.A(\game.addmisses.a[3] ),
    .B(_1701_),
    .Y(_1708_));
 sky130_fd_sc_hd__nor2_1 _4508_ (.A(_1705_),
    .B(_1708_),
    .Y(_1709_));
 sky130_fd_sc_hd__nor2_1 _4509_ (.A(_1675_),
    .B(_1697_),
    .Y(_1710_));
 sky130_fd_sc_hd__a22o_1 _4510_ (.A1(\game.addmisses.a[3] ),
    .A2(_1693_),
    .B1(_1709_),
    .B2(_1692_),
    .X(_1711_));
 sky130_fd_sc_hd__a22o_1 _4511_ (.A1(_1709_),
    .A2(_1710_),
    .B1(_1711_),
    .B2(_1675_),
    .X(\game.scoring_button_1.next_num_misses[3] ));
 sky130_fd_sc_hd__or2_1 _4512_ (.A(\game.addmisses.a[4] ),
    .B(_1697_),
    .X(_1712_));
 sky130_fd_sc_hd__and2_1 _4513_ (.A(\game.addmisses.a[4] ),
    .B(_1697_),
    .X(_1713_));
 sky130_fd_sc_hd__nor2_1 _4514_ (.A(_1675_),
    .B(_1713_),
    .Y(_1714_));
 sky130_fd_sc_hd__nand2_1 _4515_ (.A(\game.addmisses.a[4] ),
    .B(_1705_),
    .Y(_1715_));
 sky130_fd_sc_hd__nand2_1 _4516_ (.A(\modetrans.mode[0] ),
    .B(_1691_),
    .Y(_1716_));
 sky130_fd_sc_hd__o21a_1 _4517_ (.A1(_1691_),
    .A2(_1715_),
    .B1(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__or3b_1 _4518_ (.A(\game.addmisses.a[4] ),
    .B(_1691_),
    .C_N(_1705_),
    .X(_1718_));
 sky130_fd_sc_hd__a21bo_1 _4519_ (.A1(\game.addmisses.a[4] ),
    .A2(_1717_),
    .B1_N(_1718_),
    .X(_1719_));
 sky130_fd_sc_hd__a22o_1 _4520_ (.A1(_1712_),
    .A2(_1714_),
    .B1(_1719_),
    .B2(_1675_),
    .X(\game.scoring_button_1.next_num_misses[4] ));
 sky130_fd_sc_hd__or2_1 _4521_ (.A(\game.addmisses.a[5] ),
    .B(_1713_),
    .X(_1720_));
 sky130_fd_sc_hd__o21a_2 _4522_ (.A1(\game.addmisses.a[6] ),
    .A2(_1720_),
    .B1(\game.addmisses.a[7] ),
    .X(_1721_));
 sky130_fd_sc_hd__nand2_1 _4523_ (.A(\game.addmisses.a[5] ),
    .B(_1713_),
    .Y(_1722_));
 sky130_fd_sc_hd__nand2_1 _4524_ (.A(_1720_),
    .B(_1722_),
    .Y(_1723_));
 sky130_fd_sc_hd__xor2_1 _4525_ (.A(_1721_),
    .B(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__nand2_1 _4526_ (.A(\game.addmisses.a[5] ),
    .B(_1717_),
    .Y(_1725_));
 sky130_fd_sc_hd__o311a_1 _4527_ (.A1(\game.addmisses.a[5] ),
    .A2(_1691_),
    .A3(_1715_),
    .B1(_1725_),
    .C1(_1675_),
    .X(_1726_));
 sky130_fd_sc_hd__a21oi_1 _4528_ (.A1(_1699_),
    .A2(_1724_),
    .B1(_1726_),
    .Y(\game.scoring_button_1.next_num_misses[5] ));
 sky130_fd_sc_hd__inv_2 _4529_ (.A(_1721_),
    .Y(_1727_));
 sky130_fd_sc_hd__a22o_1 _4530_ (.A1(\game.addmisses.a[7] ),
    .A2(_1720_),
    .B1(_1727_),
    .B2(_1722_),
    .X(_1728_));
 sky130_fd_sc_hd__xnor2_1 _4531_ (.A(\game.addmisses.a[6] ),
    .B(_1728_),
    .Y(_1729_));
 sky130_fd_sc_hd__and4_1 _4532_ (.A(\game.addmisses.a[6] ),
    .B(\game.addmisses.a[5] ),
    .C(\game.addmisses.a[4] ),
    .D(_1705_),
    .X(_1730_));
 sky130_fd_sc_hd__a31o_1 _4533_ (.A1(\game.addmisses.a[5] ),
    .A2(\game.addmisses.a[4] ),
    .A3(_1705_),
    .B1(\game.addmisses.a[6] ),
    .X(_1731_));
 sky130_fd_sc_hd__or3b_1 _4534_ (.A(_1691_),
    .B(_1730_),
    .C_N(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__a21bo_1 _4535_ (.A1(\game.addmisses.a[6] ),
    .A2(_1693_),
    .B1_N(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__mux2_1 _4536_ (.A0(_1729_),
    .A1(_1733_),
    .S(_1675_),
    .X(_1734_));
 sky130_fd_sc_hd__clkbuf_1 _4537_ (.A(_1734_),
    .X(\game.scoring_button_1.next_num_misses[6] ));
 sky130_fd_sc_hd__a31o_1 _4538_ (.A1(\game.addmisses.a[6] ),
    .A2(\game.addmisses.a[5] ),
    .A3(_1713_),
    .B1(\game.addmisses.a[7] ),
    .X(_1735_));
 sky130_fd_sc_hd__nor2_1 _4539_ (.A(_1675_),
    .B(_1721_),
    .Y(_1736_));
 sky130_fd_sc_hd__nand2_1 _4540_ (.A(\game.addmisses.a[7] ),
    .B(_1730_),
    .Y(_1737_));
 sky130_fd_sc_hd__or2_1 _4541_ (.A(\game.addmisses.a[7] ),
    .B(_1730_),
    .X(_1738_));
 sky130_fd_sc_hd__a32o_1 _4542_ (.A1(_1692_),
    .A2(_1737_),
    .A3(_1738_),
    .B1(_1693_),
    .B2(\game.addmisses.a[7] ),
    .X(_1739_));
 sky130_fd_sc_hd__a22o_1 _4543_ (.A1(_1735_),
    .A2(_1736_),
    .B1(_1739_),
    .B2(_1675_),
    .X(\game.scoring_button_1.next_num_misses[7] ));
 sky130_fd_sc_hd__or2_1 _4544_ (.A(\game.addmisses.a[8] ),
    .B(_1721_),
    .X(_1740_));
 sky130_fd_sc_hd__and2_1 _4545_ (.A(\game.addmisses.a[8] ),
    .B(_1721_),
    .X(_1741_));
 sky130_fd_sc_hd__inv_2 _4546_ (.A(_1741_),
    .Y(_1742_));
 sky130_fd_sc_hd__nor2_2 _4547_ (.A(_1691_),
    .B(_1737_),
    .Y(_1743_));
 sky130_fd_sc_hd__and2_1 _4548_ (.A(\modetrans.mode[0] ),
    .B(_1691_),
    .X(_1744_));
 sky130_fd_sc_hd__o21ai_1 _4549_ (.A1(_1744_),
    .A2(_1743_),
    .B1(\game.addmisses.a[8] ),
    .Y(_1745_));
 sky130_fd_sc_hd__o211a_1 _4550_ (.A1(\game.addmisses.a[8] ),
    .A2(_1743_),
    .B1(_1745_),
    .C1(_1675_),
    .X(_1746_));
 sky130_fd_sc_hd__a31o_1 _4551_ (.A1(_1699_),
    .A2(_1740_),
    .A3(_1742_),
    .B1(_1746_),
    .X(\game.scoring_button_1.next_num_misses[8] ));
 sky130_fd_sc_hd__nand2_1 _4552_ (.A(\game.addmisses.a[9] ),
    .B(_1741_),
    .Y(_1747_));
 sky130_fd_sc_hd__or2_1 _4553_ (.A(\game.addmisses.a[9] ),
    .B(_1741_),
    .X(_1748_));
 sky130_fd_sc_hd__o21a_1 _4554_ (.A1(\game.addmisses.a[10] ),
    .A2(_1748_),
    .B1(\game.addmisses.a[11] ),
    .X(_1749_));
 sky130_fd_sc_hd__a21boi_1 _4555_ (.A1(_1747_),
    .A2(_1748_),
    .B1_N(_1749_),
    .Y(_1750_));
 sky130_fd_sc_hd__and3b_1 _4556_ (.A_N(\game.addmisses.a[11] ),
    .B(_1747_),
    .C(_1748_),
    .X(_1751_));
 sky130_fd_sc_hd__nand2_1 _4557_ (.A(\game.addmisses.a[8] ),
    .B(_1743_),
    .Y(_1752_));
 sky130_fd_sc_hd__o21ai_1 _4558_ (.A1(\game.addmisses.a[9] ),
    .A2(_1752_),
    .B1(_1675_),
    .Y(_1753_));
 sky130_fd_sc_hd__a31o_1 _4559_ (.A1(\game.addmisses.a[9] ),
    .A2(_1716_),
    .A3(_1752_),
    .B1(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__o31a_1 _4560_ (.A1(_1675_),
    .A2(_1750_),
    .A3(_1751_),
    .B1(_1754_),
    .X(\game.scoring_button_1.next_num_misses[9] ));
 sky130_fd_sc_hd__and3_1 _4561_ (.A(\game.addmisses.a[10] ),
    .B(\game.addmisses.a[9] ),
    .C(_1741_),
    .X(_1755_));
 sky130_fd_sc_hd__a21oi_1 _4562_ (.A1(\game.addmisses.a[9] ),
    .A2(_1741_),
    .B1(\game.addmisses.a[10] ),
    .Y(_1756_));
 sky130_fd_sc_hd__or2_1 _4563_ (.A(_1755_),
    .B(_1756_),
    .X(_1757_));
 sky130_fd_sc_hd__a2bb2o_1 _4564_ (.A1_N(_1750_),
    .A2_N(_1757_),
    .B1(_1755_),
    .B2(\game.addmisses.a[11] ),
    .X(_1758_));
 sky130_fd_sc_hd__a32o_1 _4565_ (.A1(\game.addmisses.a[9] ),
    .A2(\game.addmisses.a[8] ),
    .A3(_1743_),
    .B1(_1716_),
    .B2(\game.addmisses.a[10] ),
    .X(_1759_));
 sky130_fd_sc_hd__and4_1 _4566_ (.A(\game.addmisses.a[10] ),
    .B(\game.addmisses.a[9] ),
    .C(\game.addmisses.a[8] ),
    .D(_1743_),
    .X(_1760_));
 sky130_fd_sc_hd__nor2_1 _4567_ (.A(_1699_),
    .B(_1760_),
    .Y(_1761_));
 sky130_fd_sc_hd__a22o_1 _4568_ (.A1(_1699_),
    .A2(_1758_),
    .B1(_1759_),
    .B2(_1761_),
    .X(\game.scoring_button_1.next_num_misses[10] ));
 sky130_fd_sc_hd__nor2_1 _4569_ (.A(\game.addmisses.a[10] ),
    .B(_1748_),
    .Y(_1762_));
 sky130_fd_sc_hd__nor2_1 _4570_ (.A(_1744_),
    .B(_1760_),
    .Y(_1763_));
 sky130_fd_sc_hd__mux4_1 _4571_ (.A0(_1755_),
    .A1(_1760_),
    .A2(_1762_),
    .A3(_1763_),
    .S0(_1675_),
    .S1(\game.addmisses.a[11] ),
    .X(_1764_));
 sky130_fd_sc_hd__clkbuf_1 _4572_ (.A(_1764_),
    .X(\game.scoring_button_1.next_num_misses[11] ));
 sky130_fd_sc_hd__and2_1 _4573_ (.A(\game.addmisses.a[12] ),
    .B(_1749_),
    .X(_1765_));
 sky130_fd_sc_hd__nor2_1 _4574_ (.A(\game.addmisses.a[12] ),
    .B(_1749_),
    .Y(_1766_));
 sky130_fd_sc_hd__and3_1 _4575_ (.A(\game.addmisses.a[11] ),
    .B(_1743_),
    .C(_1755_),
    .X(_1767_));
 sky130_fd_sc_hd__nor2_1 _4576_ (.A(\game.addmisses.a[12] ),
    .B(_1767_),
    .Y(_1768_));
 sky130_fd_sc_hd__nand2_1 _4577_ (.A(net248),
    .B(_1767_),
    .Y(_1769_));
 sky130_fd_sc_hd__or4b_1 _4578_ (.A(_1699_),
    .B(_1744_),
    .C(_1768_),
    .D_N(_1769_),
    .X(_1770_));
 sky130_fd_sc_hd__o31ai_1 _4579_ (.A1(_1675_),
    .A2(_1765_),
    .A3(_1766_),
    .B1(_1770_),
    .Y(\game.scoring_button_1.next_num_misses[12] ));
 sky130_fd_sc_hd__and3_1 _4580_ (.A(\game.addmisses.a[12] ),
    .B(\game.addmisses.a[13] ),
    .C(_1749_),
    .X(_1771_));
 sky130_fd_sc_hd__nor2_1 _4581_ (.A(\game.addmisses.a[13] ),
    .B(_1765_),
    .Y(_1772_));
 sky130_fd_sc_hd__or2_1 _4582_ (.A(_1771_),
    .B(_1772_),
    .X(_1773_));
 sky130_fd_sc_hd__nand2_1 _4583_ (.A(\game.addmisses.a[15] ),
    .B(_1773_),
    .Y(_1774_));
 sky130_fd_sc_hd__o21bai_1 _4584_ (.A1(\game.addmisses.a[14] ),
    .A2(_1771_),
    .B1_N(_1774_),
    .Y(_1775_));
 sky130_fd_sc_hd__o21ai_1 _4585_ (.A1(\game.addmisses.a[15] ),
    .A2(_1773_),
    .B1(_1775_),
    .Y(_1776_));
 sky130_fd_sc_hd__and3_1 _4586_ (.A(\game.addmisses.a[13] ),
    .B(_1716_),
    .C(_1769_),
    .X(_1777_));
 sky130_fd_sc_hd__o21ai_1 _4587_ (.A1(\game.addmisses.a[13] ),
    .A2(_1769_),
    .B1(_1675_),
    .Y(_1778_));
 sky130_fd_sc_hd__o22a_1 _4588_ (.A1(_1675_),
    .A2(_1776_),
    .B1(_1777_),
    .B2(_1778_),
    .X(\game.scoring_button_1.next_num_misses[13] ));
 sky130_fd_sc_hd__and2_1 _4589_ (.A(_1767_),
    .B(_1771_),
    .X(_1779_));
 sky130_fd_sc_hd__and3_1 _4590_ (.A(\game.addmisses.a[14] ),
    .B(_1767_),
    .C(_1771_),
    .X(_1780_));
 sky130_fd_sc_hd__or2_1 _4591_ (.A(_1744_),
    .B(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__o21ba_1 _4592_ (.A1(\game.addmisses.a[14] ),
    .A2(_1779_),
    .B1_N(_1781_),
    .X(_1782_));
 sky130_fd_sc_hd__o21a_1 _4593_ (.A1(\game.addmisses.a[14] ),
    .A2(_1771_),
    .B1(_1774_),
    .X(_1783_));
 sky130_fd_sc_hd__nand2_1 _4594_ (.A(\game.addmisses.a[14] ),
    .B(_1771_),
    .Y(_1784_));
 sky130_fd_sc_hd__mux2_1 _4595_ (.A0(\game.addmisses.a[15] ),
    .A1(_1783_),
    .S(_1784_),
    .X(_1785_));
 sky130_fd_sc_hd__mux2_1 _4596_ (.A0(_1782_),
    .A1(_1785_),
    .S(_1699_),
    .X(_1786_));
 sky130_fd_sc_hd__clkbuf_1 _4597_ (.A(_1786_),
    .X(\game.scoring_button_1.next_num_misses[14] ));
 sky130_fd_sc_hd__or3_1 _4598_ (.A(\game.addmisses.a[14] ),
    .B(\game.addmisses.a[13] ),
    .C(_1765_),
    .X(_1787_));
 sky130_fd_sc_hd__mux2_1 _4599_ (.A0(_1784_),
    .A1(_1787_),
    .S(\game.addmisses.a[15] ),
    .X(_1788_));
 sky130_fd_sc_hd__nor2_1 _4600_ (.A(\game.addmisses.a[15] ),
    .B(_1780_),
    .Y(_1789_));
 sky130_fd_sc_hd__a211o_1 _4601_ (.A1(\game.addmisses.a[15] ),
    .A2(_1781_),
    .B1(_1789_),
    .C1(_1699_),
    .X(_1790_));
 sky130_fd_sc_hd__o21ai_1 _4602_ (.A1(_1675_),
    .A2(_1788_),
    .B1(_1790_),
    .Y(\game.scoring_button_1.next_num_misses[15] ));
 sky130_fd_sc_hd__buf_6 _4603_ (.A(\game.scoring_button_1.check_hit.in ),
    .X(_1791_));
 sky130_fd_sc_hd__or4b_1 _4604_ (.A(\game.scoring_button_1.flash_counter_1[5] ),
    .B(\game.scoring_button_1.flash_counter_1[4] ),
    .C(\game.scoring_button_1.flash_counter_1[7] ),
    .D_N(\game.scoring_button_1.flash_counter_1[6] ),
    .X(_1792_));
 sky130_fd_sc_hd__or4_1 _4605_ (.A(\game.scoring_button_1.flash_counter_1[1] ),
    .B(\game.scoring_button_1.flash_counter_1[0] ),
    .C(\game.scoring_button_1.flash_counter_1[3] ),
    .D(\game.scoring_button_1.flash_counter_1[2] ),
    .X(_1793_));
 sky130_fd_sc_hd__or4b_1 _4606_ (.A(\game.scoring_button_1.flash_counter_1[13] ),
    .B(\game.scoring_button_1.flash_counter_1[12] ),
    .C(\game.scoring_button_1.flash_counter_1[15] ),
    .D_N(\game.scoring_button_1.flash_counter_1[14] ),
    .X(_1794_));
 sky130_fd_sc_hd__or4b_1 _4607_ (.A(\game.scoring_button_1.flash_counter_1[8] ),
    .B(\game.scoring_button_1.flash_counter_1[11] ),
    .C(\game.scoring_button_1.flash_counter_1[10] ),
    .D_N(\game.scoring_button_1.flash_counter_1[9] ),
    .X(_1795_));
 sky130_fd_sc_hd__or3_1 _4608_ (.A(\game.scoring_button_1.flash_counter_1[21] ),
    .B(\game.scoring_button_1.flash_counter_1[20] ),
    .C(\game.scoring_button_1.flash_counter_1[22] ),
    .X(_1796_));
 sky130_fd_sc_hd__and4_1 _4609_ (.A(\game.scoring_button_1.flash_counter_1[17] ),
    .B(\game.scoring_button_1.flash_counter_1[16] ),
    .C(\game.scoring_button_1.flash_counter_1[19] ),
    .D(\game.scoring_button_1.flash_counter_1[18] ),
    .X(_1797_));
 sky130_fd_sc_hd__or4b_1 _4610_ (.A(_1794_),
    .B(_1795_),
    .C(_1796_),
    .D_N(_1797_),
    .X(_1798_));
 sky130_fd_sc_hd__o31a_2 _4611_ (.A1(_1792_),
    .A2(_1793_),
    .A3(_1798_),
    .B1(\game.hit_1 ),
    .X(_1799_));
 sky130_fd_sc_hd__a31o_1 _4612_ (.A1(_0219_),
    .A2(_1791_),
    .A3(_2656_),
    .B1(_1799_),
    .X(\game.scoring_button_1.next_good ));
 sky130_fd_sc_hd__and2b_1 _4613_ (.A_N(\game.counter[0] ),
    .B(\game.scoring_button_1.check_hit.in ),
    .X(_1800_));
 sky130_fd_sc_hd__clkbuf_1 _4614_ (.A(_1800_),
    .X(\game.scoring_button_1.next_count[0] ));
 sky130_fd_sc_hd__and3_1 _4615_ (.A(\game.scoring_button_1.check_hit.in ),
    .B(_0248_),
    .C(_1415_),
    .X(_1801_));
 sky130_fd_sc_hd__clkbuf_1 _4616_ (.A(_1801_),
    .X(\game.scoring_button_1.next_count[1] ));
 sky130_fd_sc_hd__and2_1 _4617_ (.A(_1791_),
    .B(_0024_),
    .X(_1802_));
 sky130_fd_sc_hd__clkbuf_1 _4618_ (.A(_1802_),
    .X(\game.scoring_button_1.next_count[2] ));
 sky130_fd_sc_hd__and2_1 _4619_ (.A(_1791_),
    .B(_0025_),
    .X(_1803_));
 sky130_fd_sc_hd__clkbuf_1 _4620_ (.A(_1803_),
    .X(\game.scoring_button_1.next_count[3] ));
 sky130_fd_sc_hd__and2_1 _4621_ (.A(_1791_),
    .B(_0026_),
    .X(_1804_));
 sky130_fd_sc_hd__clkbuf_1 _4622_ (.A(_1804_),
    .X(\game.scoring_button_1.next_count[4] ));
 sky130_fd_sc_hd__and2_1 _4623_ (.A(_1791_),
    .B(_0027_),
    .X(_1805_));
 sky130_fd_sc_hd__clkbuf_1 _4624_ (.A(_1805_),
    .X(\game.scoring_button_1.next_count[5] ));
 sky130_fd_sc_hd__and2_1 _4625_ (.A(_1791_),
    .B(_1426_),
    .X(_1806_));
 sky130_fd_sc_hd__clkbuf_1 _4626_ (.A(_1806_),
    .X(\game.scoring_button_1.next_count[6] ));
 sky130_fd_sc_hd__and2_1 _4627_ (.A(_1791_),
    .B(_1430_),
    .X(_1807_));
 sky130_fd_sc_hd__clkbuf_1 _4628_ (.A(_1807_),
    .X(\game.scoring_button_1.next_count[7] ));
 sky130_fd_sc_hd__and2_1 _4629_ (.A(_1791_),
    .B(_1432_),
    .X(_1808_));
 sky130_fd_sc_hd__clkbuf_1 _4630_ (.A(_1808_),
    .X(\game.scoring_button_1.next_count[8] ));
 sky130_fd_sc_hd__and2_1 _4631_ (.A(_1791_),
    .B(_1436_),
    .X(_1809_));
 sky130_fd_sc_hd__clkbuf_1 _4632_ (.A(_1809_),
    .X(\game.scoring_button_1.next_count[9] ));
 sky130_fd_sc_hd__and2_1 _4633_ (.A(_1791_),
    .B(_1440_),
    .X(_1810_));
 sky130_fd_sc_hd__clkbuf_1 _4634_ (.A(_1810_),
    .X(\game.scoring_button_1.next_count[10] ));
 sky130_fd_sc_hd__and3_1 _4635_ (.A(\game.scoring_button_1.check_hit.in ),
    .B(_1442_),
    .C(_1443_),
    .X(_1811_));
 sky130_fd_sc_hd__clkbuf_1 _4636_ (.A(_1811_),
    .X(\game.scoring_button_1.next_count[11] ));
 sky130_fd_sc_hd__and2_1 _4637_ (.A(_1791_),
    .B(_0012_),
    .X(_1812_));
 sky130_fd_sc_hd__clkbuf_1 _4638_ (.A(_1812_),
    .X(\game.scoring_button_1.next_count[12] ));
 sky130_fd_sc_hd__and2_1 _4639_ (.A(_1791_),
    .B(_0013_),
    .X(_1813_));
 sky130_fd_sc_hd__clkbuf_1 _4640_ (.A(_1813_),
    .X(\game.scoring_button_1.next_count[13] ));
 sky130_fd_sc_hd__and2_1 _4641_ (.A(_1791_),
    .B(_1452_),
    .X(_1814_));
 sky130_fd_sc_hd__clkbuf_1 _4642_ (.A(_1814_),
    .X(\game.scoring_button_1.next_count[14] ));
 sky130_fd_sc_hd__and2_1 _4643_ (.A(_1791_),
    .B(_1454_),
    .X(_1815_));
 sky130_fd_sc_hd__clkbuf_1 _4644_ (.A(_1815_),
    .X(\game.scoring_button_1.next_count[15] ));
 sky130_fd_sc_hd__and2_1 _4645_ (.A(_1791_),
    .B(_1458_),
    .X(_1816_));
 sky130_fd_sc_hd__clkbuf_1 _4646_ (.A(_1816_),
    .X(\game.scoring_button_1.next_count[16] ));
 sky130_fd_sc_hd__and2_1 _4647_ (.A(_1791_),
    .B(_0017_),
    .X(_1817_));
 sky130_fd_sc_hd__clkbuf_1 _4648_ (.A(_1817_),
    .X(\game.scoring_button_1.next_count[17] ));
 sky130_fd_sc_hd__and2_1 _4649_ (.A(_1791_),
    .B(_1463_),
    .X(_1818_));
 sky130_fd_sc_hd__clkbuf_1 _4650_ (.A(_1818_),
    .X(\game.scoring_button_1.next_count[18] ));
 sky130_fd_sc_hd__and2_1 _4651_ (.A(_1791_),
    .B(_1467_),
    .X(_1819_));
 sky130_fd_sc_hd__clkbuf_1 _4652_ (.A(_1819_),
    .X(\game.scoring_button_1.next_count[19] ));
 sky130_fd_sc_hd__and2_1 _4653_ (.A(\game.scoring_button_1.check_hit.in ),
    .B(_1471_),
    .X(_1820_));
 sky130_fd_sc_hd__clkbuf_1 _4654_ (.A(_1820_),
    .X(\game.scoring_button_1.next_count[20] ));
 sky130_fd_sc_hd__and2_1 _4655_ (.A(\game.scoring_button_1.check_hit.in ),
    .B(_1475_),
    .X(_1821_));
 sky130_fd_sc_hd__clkbuf_1 _4656_ (.A(_1821_),
    .X(\game.scoring_button_1.next_count[21] ));
 sky130_fd_sc_hd__and2_1 _4657_ (.A(\game.scoring_button_1.check_hit.in ),
    .B(_1477_),
    .X(_1822_));
 sky130_fd_sc_hd__clkbuf_1 _4658_ (.A(_1822_),
    .X(\game.scoring_button_1.next_count[22] ));
 sky130_fd_sc_hd__or4b_1 _4659_ (.A(\game.scoring_button_1.flash_counter_2[5] ),
    .B(\game.scoring_button_1.flash_counter_2[4] ),
    .C(\game.scoring_button_1.flash_counter_2[7] ),
    .D_N(\game.scoring_button_1.flash_counter_2[6] ),
    .X(_1823_));
 sky130_fd_sc_hd__or4_1 _4660_ (.A(\game.scoring_button_1.flash_counter_2[1] ),
    .B(\game.scoring_button_1.flash_counter_2[0] ),
    .C(\game.scoring_button_1.flash_counter_2[3] ),
    .D(\game.scoring_button_1.flash_counter_2[2] ),
    .X(_1824_));
 sky130_fd_sc_hd__or4b_1 _4661_ (.A(\game.scoring_button_1.flash_counter_2[13] ),
    .B(\game.scoring_button_1.flash_counter_2[12] ),
    .C(\game.scoring_button_1.flash_counter_2[15] ),
    .D_N(\game.scoring_button_1.flash_counter_2[14] ),
    .X(_1825_));
 sky130_fd_sc_hd__or4b_1 _4662_ (.A(\game.scoring_button_1.flash_counter_2[8] ),
    .B(\game.scoring_button_1.flash_counter_2[11] ),
    .C(\game.scoring_button_1.flash_counter_2[10] ),
    .D_N(\game.scoring_button_1.flash_counter_2[9] ),
    .X(_1826_));
 sky130_fd_sc_hd__or3_1 _4663_ (.A(\game.scoring_button_1.flash_counter_2[21] ),
    .B(\game.scoring_button_1.flash_counter_2[20] ),
    .C(\game.scoring_button_1.flash_counter_2[22] ),
    .X(_1827_));
 sky130_fd_sc_hd__and4_1 _4664_ (.A(\game.scoring_button_1.flash_counter_2[17] ),
    .B(\game.scoring_button_1.flash_counter_2[16] ),
    .C(\game.scoring_button_1.flash_counter_2[19] ),
    .D(\game.scoring_button_1.flash_counter_2[18] ),
    .X(_1828_));
 sky130_fd_sc_hd__or4b_1 _4665_ (.A(_1825_),
    .B(_1826_),
    .C(_1827_),
    .D_N(_1828_),
    .X(_1829_));
 sky130_fd_sc_hd__o31a_2 _4666_ (.A1(_1823_),
    .A2(_1824_),
    .A3(_1829_),
    .B1(\game.missed_1 ),
    .X(_1830_));
 sky130_fd_sc_hd__o21bai_1 _4667_ (.A1(_1791_),
    .A2(_1689_),
    .B1_N(_1830_),
    .Y(\game.scoring_button_1.next_missed ));
 sky130_fd_sc_hd__a22o_1 _4668_ (.A1(_1791_),
    .A2(_1495_),
    .B1(_1508_),
    .B2(net127),
    .X(\game.scoring_button_1.next_start_count ));
 sky130_fd_sc_hd__and2b_1 _4669_ (.A_N(\game.scoring_button_1.flash_counter_2[0] ),
    .B(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__clkbuf_1 _4670_ (.A(_1831_),
    .X(\game.scoring_button_1.next_flash_counter_2[0] ));
 sky130_fd_sc_hd__o21ai_1 _4671_ (.A1(net105),
    .A2(\game.scoring_button_1.flash_counter_2[0] ),
    .B1(\game.missed_1 ),
    .Y(_1832_));
 sky130_fd_sc_hd__a21oi_1 _4672_ (.A1(net105),
    .A2(\game.scoring_button_1.flash_counter_2[0] ),
    .B1(_1832_),
    .Y(\game.scoring_button_1.next_flash_counter_2[1] ));
 sky130_fd_sc_hd__and3_1 _4673_ (.A(\game.scoring_button_1.flash_counter_2[1] ),
    .B(\game.scoring_button_1.flash_counter_2[0] ),
    .C(\game.scoring_button_1.flash_counter_2[2] ),
    .X(_1833_));
 sky130_fd_sc_hd__a21o_1 _4674_ (.A1(\game.scoring_button_1.flash_counter_2[1] ),
    .A2(\game.scoring_button_1.flash_counter_2[0] ),
    .B1(\game.scoring_button_1.flash_counter_2[2] ),
    .X(_1834_));
 sky130_fd_sc_hd__and3b_1 _4675_ (.A_N(_1833_),
    .B(\game.missed_1 ),
    .C(_1834_),
    .X(_1835_));
 sky130_fd_sc_hd__clkbuf_1 _4676_ (.A(_1835_),
    .X(\game.scoring_button_1.next_flash_counter_2[2] ));
 sky130_fd_sc_hd__and2_1 _4677_ (.A(\game.scoring_button_1.flash_counter_2[3] ),
    .B(_1833_),
    .X(_1836_));
 sky130_fd_sc_hd__or2_1 _4678_ (.A(\game.scoring_button_1.flash_counter_2[3] ),
    .B(_1833_),
    .X(_1837_));
 sky130_fd_sc_hd__and3b_1 _4679_ (.A_N(_1836_),
    .B(\game.missed_1 ),
    .C(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__clkbuf_1 _4680_ (.A(_1838_),
    .X(\game.scoring_button_1.next_flash_counter_2[3] ));
 sky130_fd_sc_hd__a21boi_1 _4681_ (.A1(net177),
    .A2(_1836_),
    .B1_N(\game.missed_1 ),
    .Y(_1839_));
 sky130_fd_sc_hd__o21a_1 _4682_ (.A1(net177),
    .A2(_1836_),
    .B1(_1839_),
    .X(\game.scoring_button_1.next_flash_counter_2[4] ));
 sky130_fd_sc_hd__and3_1 _4683_ (.A(\game.scoring_button_1.flash_counter_2[5] ),
    .B(\game.scoring_button_1.flash_counter_2[4] ),
    .C(_1836_),
    .X(_1840_));
 sky130_fd_sc_hd__a31o_1 _4684_ (.A1(\game.scoring_button_1.flash_counter_2[3] ),
    .A2(\game.scoring_button_1.flash_counter_2[4] ),
    .A3(_1833_),
    .B1(\game.scoring_button_1.flash_counter_2[5] ),
    .X(_1841_));
 sky130_fd_sc_hd__and3b_1 _4685_ (.A_N(_1840_),
    .B(\game.missed_1 ),
    .C(_1841_),
    .X(_1842_));
 sky130_fd_sc_hd__clkbuf_1 _4686_ (.A(_1842_),
    .X(\game.scoring_button_1.next_flash_counter_2[5] ));
 sky130_fd_sc_hd__and2_1 _4687_ (.A(\game.scoring_button_1.flash_counter_2[6] ),
    .B(_1840_),
    .X(_1843_));
 sky130_fd_sc_hd__or2_1 _4688_ (.A(\game.scoring_button_1.flash_counter_2[6] ),
    .B(_1840_),
    .X(_1844_));
 sky130_fd_sc_hd__and3b_1 _4689_ (.A_N(_1843_),
    .B(_1830_),
    .C(_1844_),
    .X(_1845_));
 sky130_fd_sc_hd__clkbuf_1 _4690_ (.A(_1845_),
    .X(\game.scoring_button_1.next_flash_counter_2[6] ));
 sky130_fd_sc_hd__a21boi_1 _4691_ (.A1(net161),
    .A2(_1843_),
    .B1_N(\game.missed_1 ),
    .Y(_1846_));
 sky130_fd_sc_hd__o21a_1 _4692_ (.A1(net161),
    .A2(_1843_),
    .B1(_1846_),
    .X(\game.scoring_button_1.next_flash_counter_2[7] ));
 sky130_fd_sc_hd__and3_1 _4693_ (.A(\game.scoring_button_1.flash_counter_2[7] ),
    .B(\game.scoring_button_1.flash_counter_2[8] ),
    .C(_1843_),
    .X(_1847_));
 sky130_fd_sc_hd__a31o_1 _4694_ (.A1(\game.scoring_button_1.flash_counter_2[7] ),
    .A2(\game.scoring_button_1.flash_counter_2[6] ),
    .A3(_1840_),
    .B1(\game.scoring_button_1.flash_counter_2[8] ),
    .X(_1848_));
 sky130_fd_sc_hd__and3b_1 _4695_ (.A_N(_1847_),
    .B(\game.missed_1 ),
    .C(_1848_),
    .X(_1849_));
 sky130_fd_sc_hd__clkbuf_1 _4696_ (.A(_1849_),
    .X(\game.scoring_button_1.next_flash_counter_2[8] ));
 sky130_fd_sc_hd__and2_1 _4697_ (.A(\game.scoring_button_1.flash_counter_2[9] ),
    .B(_1847_),
    .X(_1850_));
 sky130_fd_sc_hd__or2_1 _4698_ (.A(\game.scoring_button_1.flash_counter_2[9] ),
    .B(_1847_),
    .X(_1851_));
 sky130_fd_sc_hd__and3b_1 _4699_ (.A_N(_1850_),
    .B(_1830_),
    .C(_1851_),
    .X(_1852_));
 sky130_fd_sc_hd__clkbuf_1 _4700_ (.A(_1852_),
    .X(\game.scoring_button_1.next_flash_counter_2[9] ));
 sky130_fd_sc_hd__a21boi_1 _4701_ (.A1(net158),
    .A2(_1850_),
    .B1_N(\game.missed_1 ),
    .Y(_1853_));
 sky130_fd_sc_hd__o21a_1 _4702_ (.A1(net158),
    .A2(_1850_),
    .B1(_1853_),
    .X(\game.scoring_button_1.next_flash_counter_2[10] ));
 sky130_fd_sc_hd__and3_1 _4703_ (.A(\game.scoring_button_1.flash_counter_2[11] ),
    .B(\game.scoring_button_1.flash_counter_2[10] ),
    .C(_1850_),
    .X(_1854_));
 sky130_fd_sc_hd__a31o_1 _4704_ (.A1(\game.scoring_button_1.flash_counter_2[9] ),
    .A2(\game.scoring_button_1.flash_counter_2[10] ),
    .A3(_1847_),
    .B1(\game.scoring_button_1.flash_counter_2[11] ),
    .X(_1855_));
 sky130_fd_sc_hd__and3b_1 _4705_ (.A_N(_1854_),
    .B(\game.missed_1 ),
    .C(_1855_),
    .X(_1856_));
 sky130_fd_sc_hd__clkbuf_1 _4706_ (.A(_1856_),
    .X(\game.scoring_button_1.next_flash_counter_2[11] ));
 sky130_fd_sc_hd__and2_1 _4707_ (.A(\game.scoring_button_1.flash_counter_2[12] ),
    .B(_1854_),
    .X(_1857_));
 sky130_fd_sc_hd__or2_1 _4708_ (.A(\game.scoring_button_1.flash_counter_2[12] ),
    .B(_1854_),
    .X(_1858_));
 sky130_fd_sc_hd__and3b_1 _4709_ (.A_N(_1857_),
    .B(\game.missed_1 ),
    .C(_1858_),
    .X(_1859_));
 sky130_fd_sc_hd__clkbuf_1 _4710_ (.A(_1859_),
    .X(\game.scoring_button_1.next_flash_counter_2[12] ));
 sky130_fd_sc_hd__a21boi_1 _4711_ (.A1(net184),
    .A2(_1857_),
    .B1_N(\game.missed_1 ),
    .Y(_1860_));
 sky130_fd_sc_hd__o21a_1 _4712_ (.A1(net184),
    .A2(_1857_),
    .B1(_1860_),
    .X(\game.scoring_button_1.next_flash_counter_2[13] ));
 sky130_fd_sc_hd__and3_1 _4713_ (.A(\game.scoring_button_1.flash_counter_2[13] ),
    .B(\game.scoring_button_1.flash_counter_2[14] ),
    .C(_1857_),
    .X(_1861_));
 sky130_fd_sc_hd__a31o_1 _4714_ (.A1(\game.scoring_button_1.flash_counter_2[13] ),
    .A2(\game.scoring_button_1.flash_counter_2[12] ),
    .A3(_1854_),
    .B1(\game.scoring_button_1.flash_counter_2[14] ),
    .X(_1862_));
 sky130_fd_sc_hd__and3b_1 _4715_ (.A_N(_1861_),
    .B(_1830_),
    .C(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__clkbuf_1 _4716_ (.A(_1863_),
    .X(\game.scoring_button_1.next_flash_counter_2[14] ));
 sky130_fd_sc_hd__and2_1 _4717_ (.A(\game.scoring_button_1.flash_counter_2[15] ),
    .B(_1861_),
    .X(_1864_));
 sky130_fd_sc_hd__or2_1 _4718_ (.A(\game.scoring_button_1.flash_counter_2[15] ),
    .B(_1861_),
    .X(_1865_));
 sky130_fd_sc_hd__and3b_1 _4719_ (.A_N(_1864_),
    .B(\game.missed_1 ),
    .C(_1865_),
    .X(_1866_));
 sky130_fd_sc_hd__clkbuf_1 _4720_ (.A(_1866_),
    .X(\game.scoring_button_1.next_flash_counter_2[15] ));
 sky130_fd_sc_hd__a21boi_1 _4721_ (.A1(\game.scoring_button_1.flash_counter_2[16] ),
    .A2(_1864_),
    .B1_N(_1830_),
    .Y(_1867_));
 sky130_fd_sc_hd__o21a_1 _4722_ (.A1(net194),
    .A2(_1864_),
    .B1(_1867_),
    .X(\game.scoring_button_1.next_flash_counter_2[16] ));
 sky130_fd_sc_hd__and3_1 _4723_ (.A(\game.scoring_button_1.flash_counter_2[17] ),
    .B(\game.scoring_button_1.flash_counter_2[16] ),
    .C(_1864_),
    .X(_1868_));
 sky130_fd_sc_hd__a31o_1 _4724_ (.A1(\game.scoring_button_1.flash_counter_2[15] ),
    .A2(\game.scoring_button_1.flash_counter_2[16] ),
    .A3(_1861_),
    .B1(\game.scoring_button_1.flash_counter_2[17] ),
    .X(_1869_));
 sky130_fd_sc_hd__and3b_1 _4725_ (.A_N(_1868_),
    .B(_1830_),
    .C(_1869_),
    .X(_1870_));
 sky130_fd_sc_hd__clkbuf_1 _4726_ (.A(_1870_),
    .X(\game.scoring_button_1.next_flash_counter_2[17] ));
 sky130_fd_sc_hd__and2_1 _4727_ (.A(\game.scoring_button_1.flash_counter_2[18] ),
    .B(_1868_),
    .X(_1871_));
 sky130_fd_sc_hd__or2_1 _4728_ (.A(\game.scoring_button_1.flash_counter_2[18] ),
    .B(_1868_),
    .X(_1872_));
 sky130_fd_sc_hd__and3b_1 _4729_ (.A_N(_1871_),
    .B(_1830_),
    .C(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__clkbuf_1 _4730_ (.A(_1873_),
    .X(\game.scoring_button_1.next_flash_counter_2[18] ));
 sky130_fd_sc_hd__a21boi_1 _4731_ (.A1(net181),
    .A2(_1871_),
    .B1_N(_1830_),
    .Y(_1874_));
 sky130_fd_sc_hd__o21a_1 _4732_ (.A1(net181),
    .A2(_1871_),
    .B1(_1874_),
    .X(\game.scoring_button_1.next_flash_counter_2[19] ));
 sky130_fd_sc_hd__and3_1 _4733_ (.A(\game.scoring_button_1.flash_counter_2[19] ),
    .B(\game.scoring_button_1.flash_counter_2[20] ),
    .C(_1871_),
    .X(_1875_));
 sky130_fd_sc_hd__a31o_1 _4734_ (.A1(\game.scoring_button_1.flash_counter_2[19] ),
    .A2(\game.scoring_button_1.flash_counter_2[18] ),
    .A3(_1868_),
    .B1(\game.scoring_button_1.flash_counter_2[20] ),
    .X(_1876_));
 sky130_fd_sc_hd__and3b_1 _4735_ (.A_N(_1875_),
    .B(\game.missed_1 ),
    .C(_1876_),
    .X(_1877_));
 sky130_fd_sc_hd__clkbuf_1 _4736_ (.A(_1877_),
    .X(\game.scoring_button_1.next_flash_counter_2[20] ));
 sky130_fd_sc_hd__and2_1 _4737_ (.A(\game.scoring_button_1.flash_counter_2[21] ),
    .B(_1875_),
    .X(_1878_));
 sky130_fd_sc_hd__or2_1 _4738_ (.A(\game.scoring_button_1.flash_counter_2[21] ),
    .B(_1875_),
    .X(_1879_));
 sky130_fd_sc_hd__and3b_1 _4739_ (.A_N(_1878_),
    .B(\game.missed_1 ),
    .C(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__clkbuf_1 _4740_ (.A(_1880_),
    .X(\game.scoring_button_1.next_flash_counter_2[21] ));
 sky130_fd_sc_hd__o21ai_1 _4741_ (.A1(net86),
    .A2(_1878_),
    .B1(\game.missed_1 ),
    .Y(_1881_));
 sky130_fd_sc_hd__a21oi_1 _4742_ (.A1(net86),
    .A2(_1878_),
    .B1(_1881_),
    .Y(\game.scoring_button_1.next_flash_counter_2[22] ));
 sky130_fd_sc_hd__and2b_1 _4743_ (.A_N(\game.scoring_button_1.flash_counter_1[0] ),
    .B(_1799_),
    .X(_1882_));
 sky130_fd_sc_hd__clkbuf_1 _4744_ (.A(_1882_),
    .X(\game.scoring_button_1.next_flash_counter_1[0] ));
 sky130_fd_sc_hd__o21ai_1 _4745_ (.A1(net111),
    .A2(\game.scoring_button_1.flash_counter_1[0] ),
    .B1(\game.hit_1 ),
    .Y(_1883_));
 sky130_fd_sc_hd__a21oi_1 _4746_ (.A1(net111),
    .A2(\game.scoring_button_1.flash_counter_1[0] ),
    .B1(_1883_),
    .Y(\game.scoring_button_1.next_flash_counter_1[1] ));
 sky130_fd_sc_hd__and3_1 _4747_ (.A(\game.scoring_button_1.flash_counter_1[1] ),
    .B(\game.scoring_button_1.flash_counter_1[0] ),
    .C(\game.scoring_button_1.flash_counter_1[2] ),
    .X(_1884_));
 sky130_fd_sc_hd__a21o_1 _4748_ (.A1(\game.scoring_button_1.flash_counter_1[1] ),
    .A2(\game.scoring_button_1.flash_counter_1[0] ),
    .B1(\game.scoring_button_1.flash_counter_1[2] ),
    .X(_1885_));
 sky130_fd_sc_hd__and3b_1 _4749_ (.A_N(_1884_),
    .B(\game.hit_1 ),
    .C(_1885_),
    .X(_1886_));
 sky130_fd_sc_hd__clkbuf_1 _4750_ (.A(_1886_),
    .X(\game.scoring_button_1.next_flash_counter_1[2] ));
 sky130_fd_sc_hd__and2_1 _4751_ (.A(\game.scoring_button_1.flash_counter_1[3] ),
    .B(_1884_),
    .X(_1887_));
 sky130_fd_sc_hd__or2_1 _4752_ (.A(\game.scoring_button_1.flash_counter_1[3] ),
    .B(_1884_),
    .X(_1888_));
 sky130_fd_sc_hd__and3b_1 _4753_ (.A_N(_1887_),
    .B(\game.hit_1 ),
    .C(_1888_),
    .X(_1889_));
 sky130_fd_sc_hd__clkbuf_1 _4754_ (.A(_1889_),
    .X(\game.scoring_button_1.next_flash_counter_1[3] ));
 sky130_fd_sc_hd__a21boi_1 _4755_ (.A1(\game.scoring_button_1.flash_counter_1[4] ),
    .A2(_1887_),
    .B1_N(\game.hit_1 ),
    .Y(_1890_));
 sky130_fd_sc_hd__o21a_1 _4756_ (.A1(net207),
    .A2(_1887_),
    .B1(_1890_),
    .X(\game.scoring_button_1.next_flash_counter_1[4] ));
 sky130_fd_sc_hd__and3_1 _4757_ (.A(\game.scoring_button_1.flash_counter_1[5] ),
    .B(\game.scoring_button_1.flash_counter_1[4] ),
    .C(_1887_),
    .X(_1891_));
 sky130_fd_sc_hd__a31o_1 _4758_ (.A1(\game.scoring_button_1.flash_counter_1[3] ),
    .A2(\game.scoring_button_1.flash_counter_1[4] ),
    .A3(_1884_),
    .B1(\game.scoring_button_1.flash_counter_1[5] ),
    .X(_1892_));
 sky130_fd_sc_hd__and3b_1 _4759_ (.A_N(_1891_),
    .B(\game.hit_1 ),
    .C(_1892_),
    .X(_1893_));
 sky130_fd_sc_hd__clkbuf_1 _4760_ (.A(_1893_),
    .X(\game.scoring_button_1.next_flash_counter_1[5] ));
 sky130_fd_sc_hd__and2_1 _4761_ (.A(\game.scoring_button_1.flash_counter_1[6] ),
    .B(_1891_),
    .X(_1894_));
 sky130_fd_sc_hd__or2_1 _4762_ (.A(\game.scoring_button_1.flash_counter_1[6] ),
    .B(_1891_),
    .X(_1895_));
 sky130_fd_sc_hd__and3b_1 _4763_ (.A_N(_1894_),
    .B(_1799_),
    .C(_1895_),
    .X(_1896_));
 sky130_fd_sc_hd__clkbuf_1 _4764_ (.A(_1896_),
    .X(\game.scoring_button_1.next_flash_counter_1[6] ));
 sky130_fd_sc_hd__a21boi_1 _4765_ (.A1(net162),
    .A2(_1894_),
    .B1_N(\game.hit_1 ),
    .Y(_1897_));
 sky130_fd_sc_hd__o21a_1 _4766_ (.A1(net162),
    .A2(_1894_),
    .B1(_1897_),
    .X(\game.scoring_button_1.next_flash_counter_1[7] ));
 sky130_fd_sc_hd__and3_1 _4767_ (.A(\game.scoring_button_1.flash_counter_1[7] ),
    .B(\game.scoring_button_1.flash_counter_1[8] ),
    .C(_1894_),
    .X(_1898_));
 sky130_fd_sc_hd__a31o_1 _4768_ (.A1(\game.scoring_button_1.flash_counter_1[7] ),
    .A2(\game.scoring_button_1.flash_counter_1[6] ),
    .A3(_1891_),
    .B1(\game.scoring_button_1.flash_counter_1[8] ),
    .X(_1899_));
 sky130_fd_sc_hd__and3b_1 _4769_ (.A_N(_1898_),
    .B(\game.hit_1 ),
    .C(_1899_),
    .X(_1900_));
 sky130_fd_sc_hd__clkbuf_1 _4770_ (.A(_1900_),
    .X(\game.scoring_button_1.next_flash_counter_1[8] ));
 sky130_fd_sc_hd__and2_1 _4771_ (.A(\game.scoring_button_1.flash_counter_1[9] ),
    .B(_1898_),
    .X(_1901_));
 sky130_fd_sc_hd__or2_1 _4772_ (.A(\game.scoring_button_1.flash_counter_1[9] ),
    .B(_1898_),
    .X(_1902_));
 sky130_fd_sc_hd__and3b_1 _4773_ (.A_N(_1901_),
    .B(_1799_),
    .C(_1902_),
    .X(_1903_));
 sky130_fd_sc_hd__clkbuf_1 _4774_ (.A(_1903_),
    .X(\game.scoring_button_1.next_flash_counter_1[9] ));
 sky130_fd_sc_hd__a21boi_1 _4775_ (.A1(net157),
    .A2(_1901_),
    .B1_N(\game.hit_1 ),
    .Y(_1904_));
 sky130_fd_sc_hd__o21a_1 _4776_ (.A1(net157),
    .A2(_1901_),
    .B1(_1904_),
    .X(\game.scoring_button_1.next_flash_counter_1[10] ));
 sky130_fd_sc_hd__and3_1 _4777_ (.A(\game.scoring_button_1.flash_counter_1[11] ),
    .B(\game.scoring_button_1.flash_counter_1[10] ),
    .C(_1901_),
    .X(_1905_));
 sky130_fd_sc_hd__a31o_1 _4778_ (.A1(\game.scoring_button_1.flash_counter_1[9] ),
    .A2(\game.scoring_button_1.flash_counter_1[10] ),
    .A3(_1898_),
    .B1(\game.scoring_button_1.flash_counter_1[11] ),
    .X(_1906_));
 sky130_fd_sc_hd__and3b_1 _4779_ (.A_N(_1905_),
    .B(\game.hit_1 ),
    .C(_1906_),
    .X(_1907_));
 sky130_fd_sc_hd__clkbuf_1 _4780_ (.A(_1907_),
    .X(\game.scoring_button_1.next_flash_counter_1[11] ));
 sky130_fd_sc_hd__and2_1 _4781_ (.A(\game.scoring_button_1.flash_counter_1[12] ),
    .B(_1905_),
    .X(_1908_));
 sky130_fd_sc_hd__or2_1 _4782_ (.A(\game.scoring_button_1.flash_counter_1[12] ),
    .B(_1905_),
    .X(_1909_));
 sky130_fd_sc_hd__and3b_1 _4783_ (.A_N(_1908_),
    .B(\game.hit_1 ),
    .C(_1909_),
    .X(_1910_));
 sky130_fd_sc_hd__clkbuf_1 _4784_ (.A(_1910_),
    .X(\game.scoring_button_1.next_flash_counter_1[12] ));
 sky130_fd_sc_hd__a21boi_1 _4785_ (.A1(net155),
    .A2(_1908_),
    .B1_N(\game.hit_1 ),
    .Y(_1911_));
 sky130_fd_sc_hd__o21a_1 _4786_ (.A1(net155),
    .A2(_1908_),
    .B1(_1911_),
    .X(\game.scoring_button_1.next_flash_counter_1[13] ));
 sky130_fd_sc_hd__and3_1 _4787_ (.A(\game.scoring_button_1.flash_counter_1[13] ),
    .B(\game.scoring_button_1.flash_counter_1[14] ),
    .C(_1908_),
    .X(_1912_));
 sky130_fd_sc_hd__a31o_1 _4788_ (.A1(\game.scoring_button_1.flash_counter_1[13] ),
    .A2(\game.scoring_button_1.flash_counter_1[12] ),
    .A3(_1905_),
    .B1(\game.scoring_button_1.flash_counter_1[14] ),
    .X(_1913_));
 sky130_fd_sc_hd__and3b_1 _4789_ (.A_N(_1912_),
    .B(_1799_),
    .C(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__clkbuf_1 _4790_ (.A(_1914_),
    .X(\game.scoring_button_1.next_flash_counter_1[14] ));
 sky130_fd_sc_hd__and2_1 _4791_ (.A(\game.scoring_button_1.flash_counter_1[15] ),
    .B(_1912_),
    .X(_1915_));
 sky130_fd_sc_hd__or2_1 _4792_ (.A(\game.scoring_button_1.flash_counter_1[15] ),
    .B(_1912_),
    .X(_1916_));
 sky130_fd_sc_hd__and3b_1 _4793_ (.A_N(_1915_),
    .B(\game.hit_1 ),
    .C(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__clkbuf_1 _4794_ (.A(_1917_),
    .X(\game.scoring_button_1.next_flash_counter_1[15] ));
 sky130_fd_sc_hd__a21boi_1 _4795_ (.A1(net180),
    .A2(_1915_),
    .B1_N(_1799_),
    .Y(_1918_));
 sky130_fd_sc_hd__o21a_1 _4796_ (.A1(net180),
    .A2(_1915_),
    .B1(_1918_),
    .X(\game.scoring_button_1.next_flash_counter_1[16] ));
 sky130_fd_sc_hd__and3_1 _4797_ (.A(\game.scoring_button_1.flash_counter_1[17] ),
    .B(\game.scoring_button_1.flash_counter_1[16] ),
    .C(_1915_),
    .X(_1919_));
 sky130_fd_sc_hd__a31o_1 _4798_ (.A1(\game.scoring_button_1.flash_counter_1[15] ),
    .A2(\game.scoring_button_1.flash_counter_1[16] ),
    .A3(_1912_),
    .B1(\game.scoring_button_1.flash_counter_1[17] ),
    .X(_1920_));
 sky130_fd_sc_hd__and3b_1 _4799_ (.A_N(_1919_),
    .B(_1799_),
    .C(_1920_),
    .X(_1921_));
 sky130_fd_sc_hd__clkbuf_1 _4800_ (.A(_1921_),
    .X(\game.scoring_button_1.next_flash_counter_1[17] ));
 sky130_fd_sc_hd__and2_1 _4801_ (.A(\game.scoring_button_1.flash_counter_1[18] ),
    .B(_1919_),
    .X(_1922_));
 sky130_fd_sc_hd__or2_1 _4802_ (.A(\game.scoring_button_1.flash_counter_1[18] ),
    .B(_1919_),
    .X(_1923_));
 sky130_fd_sc_hd__and3b_1 _4803_ (.A_N(_1922_),
    .B(_1799_),
    .C(_1923_),
    .X(_1924_));
 sky130_fd_sc_hd__clkbuf_1 _4804_ (.A(_1924_),
    .X(\game.scoring_button_1.next_flash_counter_1[18] ));
 sky130_fd_sc_hd__a21boi_1 _4805_ (.A1(net172),
    .A2(_1922_),
    .B1_N(_1799_),
    .Y(_1925_));
 sky130_fd_sc_hd__o21a_1 _4806_ (.A1(net172),
    .A2(_1922_),
    .B1(_1925_),
    .X(\game.scoring_button_1.next_flash_counter_1[19] ));
 sky130_fd_sc_hd__and3_1 _4807_ (.A(\game.scoring_button_1.flash_counter_1[19] ),
    .B(\game.scoring_button_1.flash_counter_1[20] ),
    .C(_1922_),
    .X(_1926_));
 sky130_fd_sc_hd__a31o_1 _4808_ (.A1(\game.scoring_button_1.flash_counter_1[19] ),
    .A2(\game.scoring_button_1.flash_counter_1[18] ),
    .A3(_1919_),
    .B1(\game.scoring_button_1.flash_counter_1[20] ),
    .X(_1927_));
 sky130_fd_sc_hd__and3b_1 _4809_ (.A_N(_1926_),
    .B(\game.hit_1 ),
    .C(_1927_),
    .X(_1928_));
 sky130_fd_sc_hd__clkbuf_1 _4810_ (.A(_1928_),
    .X(\game.scoring_button_1.next_flash_counter_1[20] ));
 sky130_fd_sc_hd__and2_1 _4811_ (.A(\game.scoring_button_1.flash_counter_1[21] ),
    .B(_1926_),
    .X(_1929_));
 sky130_fd_sc_hd__or2_1 _4812_ (.A(\game.scoring_button_1.flash_counter_1[21] ),
    .B(_1926_),
    .X(_1930_));
 sky130_fd_sc_hd__and3b_1 _4813_ (.A_N(_1929_),
    .B(\game.hit_1 ),
    .C(_1930_),
    .X(_1931_));
 sky130_fd_sc_hd__clkbuf_1 _4814_ (.A(_1931_),
    .X(\game.scoring_button_1.next_flash_counter_1[21] ));
 sky130_fd_sc_hd__o21ai_1 _4815_ (.A1(net85),
    .A2(_1929_),
    .B1(\game.hit_1 ),
    .Y(_1932_));
 sky130_fd_sc_hd__a21oi_1 _4816_ (.A1(net85),
    .A2(_1929_),
    .B1(_1932_),
    .Y(\game.scoring_button_1.next_flash_counter_1[22] ));
 sky130_fd_sc_hd__nor2_1 _4817_ (.A(net109),
    .B(_0032_),
    .Y(_0009_));
 sky130_fd_sc_hd__and2_1 _4818_ (.A(_0248_),
    .B(_1415_),
    .X(_1933_));
 sky130_fd_sc_hd__clkbuf_1 _4819_ (.A(_1933_),
    .X(_0020_));
 sky130_fd_sc_hd__o21a_1 _4820_ (.A1(_0232_),
    .A2(_0254_),
    .B1(_1426_),
    .X(_0028_));
 sky130_fd_sc_hd__and2b_1 _4821_ (.A_N(_0032_),
    .B(_1430_),
    .X(_1934_));
 sky130_fd_sc_hd__clkbuf_1 _4822_ (.A(_1934_),
    .X(_0029_));
 sky130_fd_sc_hd__o21a_1 _4823_ (.A1(_0232_),
    .A2(_0254_),
    .B1(_1432_),
    .X(_0030_));
 sky130_fd_sc_hd__o21a_1 _4824_ (.A1(_0232_),
    .A2(_0254_),
    .B1(_1436_),
    .X(_0031_));
 sky130_fd_sc_hd__and2b_1 _4825_ (.A_N(_0032_),
    .B(_1440_),
    .X(_1935_));
 sky130_fd_sc_hd__clkbuf_1 _4826_ (.A(_1935_),
    .X(_0010_));
 sky130_fd_sc_hd__and3b_1 _4827_ (.A_N(_0032_),
    .B(_1442_),
    .C(_1443_),
    .X(_1936_));
 sky130_fd_sc_hd__clkbuf_1 _4828_ (.A(_1936_),
    .X(_0011_));
 sky130_fd_sc_hd__and2b_1 _4829_ (.A_N(_0032_),
    .B(_1452_),
    .X(_1937_));
 sky130_fd_sc_hd__clkbuf_1 _4830_ (.A(_1937_),
    .X(_0014_));
 sky130_fd_sc_hd__and2b_1 _4831_ (.A_N(_0032_),
    .B(_1454_),
    .X(_1938_));
 sky130_fd_sc_hd__clkbuf_1 _4832_ (.A(_1938_),
    .X(_0015_));
 sky130_fd_sc_hd__and2b_1 _4833_ (.A_N(_0032_),
    .B(_1458_),
    .X(_1939_));
 sky130_fd_sc_hd__clkbuf_1 _4834_ (.A(_1939_),
    .X(_0016_));
 sky130_fd_sc_hd__and2b_1 _4835_ (.A_N(_0032_),
    .B(_1463_),
    .X(_1940_));
 sky130_fd_sc_hd__clkbuf_1 _4836_ (.A(_1940_),
    .X(_0018_));
 sky130_fd_sc_hd__and2b_1 _4837_ (.A_N(_0032_),
    .B(_1467_),
    .X(_1941_));
 sky130_fd_sc_hd__clkbuf_1 _4838_ (.A(_1941_),
    .X(_0019_));
 sky130_fd_sc_hd__and2b_1 _4839_ (.A_N(_0032_),
    .B(_1471_),
    .X(_1942_));
 sky130_fd_sc_hd__clkbuf_1 _4840_ (.A(_1942_),
    .X(_0021_));
 sky130_fd_sc_hd__and2b_1 _4841_ (.A_N(_0032_),
    .B(_1475_),
    .X(_1943_));
 sky130_fd_sc_hd__clkbuf_1 _4842_ (.A(_1943_),
    .X(_0022_));
 sky130_fd_sc_hd__and2b_1 _4843_ (.A_N(_0032_),
    .B(_1477_),
    .X(_1944_));
 sky130_fd_sc_hd__clkbuf_1 _4844_ (.A(_1944_),
    .X(_0023_));
 sky130_fd_sc_hd__o22a_1 _4845_ (.A1(\disp_song.um.idx_note2[0] ),
    .A2(_0325_),
    .B1(_0366_),
    .B2(\disp_song.um.idx_note1[0] ),
    .X(\disp_song.um.next_position[0] ));
 sky130_fd_sc_hd__o22a_1 _4846_ (.A1(\disp_song.um.idx_note2[1] ),
    .A2(_0325_),
    .B1(_0366_),
    .B2(_0179_),
    .X(\disp_song.um.next_position[1] ));
 sky130_fd_sc_hd__o22a_1 _4847_ (.A1(net266),
    .A2(_0325_),
    .B1(_0366_),
    .B2(\disp_song.um.idx_note1[2] ),
    .X(\disp_song.um.next_position[2] ));
 sky130_fd_sc_hd__mux2_1 _4848_ (.A0(\disp_song.um.idx_note1[3] ),
    .A1(\disp_song.um.idx_note2[3] ),
    .S(_2661_),
    .X(_1945_));
 sky130_fd_sc_hd__or2_1 _4849_ (.A(_0352_),
    .B(_1945_),
    .X(_1946_));
 sky130_fd_sc_hd__clkbuf_1 _4850_ (.A(_1946_),
    .X(\disp_song.um.next_position[3] ));
 sky130_fd_sc_hd__or3b_1 _4851_ (.A(_0405_),
    .B(_0352_),
    .C_N(_0316_),
    .X(_1947_));
 sky130_fd_sc_hd__clkbuf_1 _4852_ (.A(_1947_),
    .X(\disp_song.um.next_position[4] ));
 sky130_fd_sc_hd__nor2_2 _4853_ (.A(_2666_),
    .B(_0169_),
    .Y(_1948_));
 sky130_fd_sc_hd__nand2_4 _4854_ (.A(_2677_),
    .B(_0162_),
    .Y(_1949_));
 sky130_fd_sc_hd__nor2_2 _4855_ (.A(_1948_),
    .B(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__nor2_1 _4856_ (.A(\disp_song.um.drum.next_idx2[3] ),
    .B(_1948_),
    .Y(_1951_));
 sky130_fd_sc_hd__nor2_1 _4857_ (.A(_0162_),
    .B(_1951_),
    .Y(_1952_));
 sky130_fd_sc_hd__nor2_1 _4858_ (.A(_1950_),
    .B(_1952_),
    .Y(_1953_));
 sky130_fd_sc_hd__inv_2 _4859_ (.A(\disp_song.um.drum.next_note2[26] ),
    .Y(_1954_));
 sky130_fd_sc_hd__mux2_1 _4860_ (.A0(_1954_),
    .A1(_0343_),
    .S(\disp_song.um.drum.next_idx2[0] ),
    .X(_1955_));
 sky130_fd_sc_hd__clkbuf_8 _4861_ (.A(_2669_),
    .X(_1956_));
 sky130_fd_sc_hd__or2_1 _4862_ (.A(_1956_),
    .B(\disp_song.um.drum.next_note2[25] ),
    .X(_1957_));
 sky130_fd_sc_hd__o21ai_1 _4863_ (.A1(\disp_song.um.drum.next_idx2[0] ),
    .A2(\disp_song.um.drum.next_note2[24] ),
    .B1(_1957_),
    .Y(_1958_));
 sky130_fd_sc_hd__mux2_1 _4864_ (.A0(_1955_),
    .A1(_1958_),
    .S(\disp_song.um.drum.next_idx2[1] ),
    .X(_1959_));
 sky130_fd_sc_hd__nor2_1 _4865_ (.A(_2679_),
    .B(_0169_),
    .Y(_1960_));
 sky130_fd_sc_hd__a21oi_2 _4866_ (.A1(\disp_song.um.drum.next_idx2[1] ),
    .A2(_1960_),
    .B1(_1951_),
    .Y(_1961_));
 sky130_fd_sc_hd__nor2_1 _4867_ (.A(\disp_song.um.drum.next_idx2[1] ),
    .B(_1949_),
    .Y(_1962_));
 sky130_fd_sc_hd__or2_1 _4868_ (.A(_1961_),
    .B(_1962_),
    .X(_1963_));
 sky130_fd_sc_hd__or2_1 _4869_ (.A(_1948_),
    .B(_1949_),
    .X(_1964_));
 sky130_fd_sc_hd__buf_4 _4870_ (.A(_1964_),
    .X(_1965_));
 sky130_fd_sc_hd__mux2_2 _4871_ (.A0(\disp_song.um.drum.next_note2[18] ),
    .A1(\disp_song.um.drum.next_note2[19] ),
    .S(\disp_song.um.drum.next_idx2[0] ),
    .X(_1966_));
 sky130_fd_sc_hd__or2_1 _4872_ (.A(\disp_song.um.drum.next_idx2[2] ),
    .B(_1949_),
    .X(_1967_));
 sky130_fd_sc_hd__clkbuf_4 _4873_ (.A(_1967_),
    .X(_1968_));
 sky130_fd_sc_hd__mux2_1 _4874_ (.A0(\disp_song.um.drum.next_note2[16] ),
    .A1(\disp_song.um.drum.next_note2[17] ),
    .S(_2670_),
    .X(_1969_));
 sky130_fd_sc_hd__and3_1 _4875_ (.A(\disp_song.um.drum.next_idx2[1] ),
    .B(_1968_),
    .C(_1969_),
    .X(_1970_));
 sky130_fd_sc_hd__a31o_1 _4876_ (.A1(_0169_),
    .A2(_1965_),
    .A3(_1966_),
    .B1(_1970_),
    .X(_1971_));
 sky130_fd_sc_hd__a2bb2o_1 _4877_ (.A1_N(_1959_),
    .A2_N(_1963_),
    .B1(_1971_),
    .B2(_1961_),
    .X(_1972_));
 sky130_fd_sc_hd__mux2_1 _4878_ (.A0(\disp_song.um.drum.next_note2[28] ),
    .A1(\disp_song.um.drum.next_note2[29] ),
    .S(_2670_),
    .X(_1973_));
 sky130_fd_sc_hd__and3_1 _4879_ (.A(\disp_song.um.drum.next_idx2[1] ),
    .B(_1968_),
    .C(_1973_),
    .X(_1974_));
 sky130_fd_sc_hd__or2_1 _4880_ (.A(_2670_),
    .B(\disp_song.um.drum.next_note2[30] ),
    .X(_1975_));
 sky130_fd_sc_hd__o21ai_1 _4881_ (.A1(_2669_),
    .A2(\disp_song.um.drum.next_note2[31] ),
    .B1(_1975_),
    .Y(_1976_));
 sky130_fd_sc_hd__and3b_1 _4882_ (.A_N(_1976_),
    .B(_2666_),
    .C(_1965_),
    .X(_1977_));
 sky130_fd_sc_hd__mux2_1 _4883_ (.A0(\disp_song.um.drum.next_note2[22] ),
    .A1(\disp_song.um.drum.next_note2[23] ),
    .S(\disp_song.um.drum.next_idx2[0] ),
    .X(_1978_));
 sky130_fd_sc_hd__mux2_1 _4884_ (.A0(\disp_song.um.drum.next_note2[20] ),
    .A1(\disp_song.um.drum.next_note2[21] ),
    .S(\disp_song.um.drum.next_idx2[0] ),
    .X(_1979_));
 sky130_fd_sc_hd__mux2_1 _4885_ (.A0(_1978_),
    .A1(_1979_),
    .S(\disp_song.um.drum.next_idx2[1] ),
    .X(_1980_));
 sky130_fd_sc_hd__o32a_1 _4886_ (.A1(_1961_),
    .A2(_1974_),
    .A3(_1977_),
    .B1(_1980_),
    .B2(_2679_),
    .X(_1981_));
 sky130_fd_sc_hd__and2_1 _4887_ (.A(_2664_),
    .B(_0169_),
    .X(_1982_));
 sky130_fd_sc_hd__nor2_4 _4888_ (.A(_1948_),
    .B(_1982_),
    .Y(_1983_));
 sky130_fd_sc_hd__mux2_1 _4889_ (.A0(_1972_),
    .A1(_1981_),
    .S(_1983_),
    .X(_1984_));
 sky130_fd_sc_hd__or2_1 _4890_ (.A(\disp_song.um.drum.next_idx2[0] ),
    .B(\disp_song.um.drum.next_note2[10] ),
    .X(_1985_));
 sky130_fd_sc_hd__o21ai_1 _4891_ (.A1(_1956_),
    .A2(\disp_song.um.drum.next_note2[11] ),
    .B1(_1985_),
    .Y(_1986_));
 sky130_fd_sc_hd__or2_1 _4892_ (.A(\disp_song.um.drum.next_idx2[0] ),
    .B(\disp_song.um.drum.next_note2[8] ),
    .X(_1987_));
 sky130_fd_sc_hd__o21ai_1 _4893_ (.A1(_1956_),
    .A2(\disp_song.um.drum.next_note2[9] ),
    .B1(_1987_),
    .Y(_1988_));
 sky130_fd_sc_hd__mux2_1 _4894_ (.A0(_1986_),
    .A1(_1988_),
    .S(\disp_song.um.drum.next_idx2[1] ),
    .X(_1989_));
 sky130_fd_sc_hd__nor2_1 _4895_ (.A(_1962_),
    .B(_1989_),
    .Y(_1990_));
 sky130_fd_sc_hd__mux2_1 _4896_ (.A0(\disp_song.um.drum.next_note2[14] ),
    .A1(\disp_song.um.drum.next_note2[15] ),
    .S(_2670_),
    .X(_1991_));
 sky130_fd_sc_hd__nor2_4 _4897_ (.A(\disp_song.um.drum.next_idx2[2] ),
    .B(_1949_),
    .Y(_1992_));
 sky130_fd_sc_hd__or2_1 _4898_ (.A(_2670_),
    .B(\disp_song.um.drum.next_note2[12] ),
    .X(_1993_));
 sky130_fd_sc_hd__o21ai_1 _4899_ (.A1(_1956_),
    .A2(\disp_song.um.drum.next_note2[13] ),
    .B1(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__or2_1 _4900_ (.A(_2666_),
    .B(_1994_),
    .X(_1995_));
 sky130_fd_sc_hd__nor2_1 _4901_ (.A(_1992_),
    .B(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__a31o_1 _4902_ (.A1(_2666_),
    .A2(_1965_),
    .A3(_1991_),
    .B1(_1996_),
    .X(_1997_));
 sky130_fd_sc_hd__mux2_1 _4903_ (.A0(_1990_),
    .A1(_1997_),
    .S(_1983_),
    .X(_1998_));
 sky130_fd_sc_hd__mux2_1 _4904_ (.A0(\disp_song.um.drum.next_note2[0] ),
    .A1(\disp_song.um.drum.next_note2[1] ),
    .S(_2670_),
    .X(_1999_));
 sky130_fd_sc_hd__nand2_1 _4905_ (.A(\disp_song.um.drum.next_idx2[1] ),
    .B(_1999_),
    .Y(_2000_));
 sky130_fd_sc_hd__mux2_1 _4906_ (.A0(\disp_song.um.drum.next_note2[2] ),
    .A1(\disp_song.um.drum.next_note2[3] ),
    .S(_2670_),
    .X(_2001_));
 sky130_fd_sc_hd__a2bb2o_1 _4907_ (.A1_N(_1992_),
    .A2_N(_2000_),
    .B1(_2001_),
    .B2(_2666_),
    .X(_2002_));
 sky130_fd_sc_hd__mux2_1 _4908_ (.A0(\disp_song.um.drum.next_note2[6] ),
    .A1(\disp_song.um.drum.next_note2[7] ),
    .S(\disp_song.um.drum.next_idx2[0] ),
    .X(_2003_));
 sky130_fd_sc_hd__mux2_1 _4909_ (.A0(\disp_song.um.drum.next_note2[4] ),
    .A1(\disp_song.um.drum.next_note2[5] ),
    .S(\disp_song.um.drum.next_idx2[0] ),
    .X(_2004_));
 sky130_fd_sc_hd__mux2_1 _4910_ (.A0(_2003_),
    .A1(_2004_),
    .S(\disp_song.um.drum.next_idx2[1] ),
    .X(_2005_));
 sky130_fd_sc_hd__mux2_1 _4911_ (.A0(_2002_),
    .A1(_2005_),
    .S(_1983_),
    .X(_2006_));
 sky130_fd_sc_hd__mux2_1 _4912_ (.A0(_1998_),
    .A1(_2006_),
    .S(_1961_),
    .X(_2007_));
 sky130_fd_sc_hd__o211a_1 _4913_ (.A1(_1952_),
    .A2(_2007_),
    .B1(_0214_),
    .C1(_1965_),
    .X(_2008_));
 sky130_fd_sc_hd__o21a_1 _4914_ (.A1(_1953_),
    .A2(_1984_),
    .B1(_2008_),
    .X(\disp_song.um.drum.next_d2[0] ));
 sky130_fd_sc_hd__nand2_2 _4915_ (.A(_2664_),
    .B(_2669_),
    .Y(_2009_));
 sky130_fd_sc_hd__and2_2 _4916_ (.A(\disp_song.um.drum.next_idx2[2] ),
    .B(_2009_),
    .X(_2010_));
 sky130_fd_sc_hd__o21a_1 _4917_ (.A1(\disp_song.um.drum.next_idx2[3] ),
    .A2(_2010_),
    .B1(\disp_song.um.drum.next_idx2[4] ),
    .X(_2011_));
 sky130_fd_sc_hd__nor2_2 _4918_ (.A(\disp_song.um.drum.next_idx2[2] ),
    .B(_2009_),
    .Y(_2012_));
 sky130_fd_sc_hd__or2_2 _4919_ (.A(_2010_),
    .B(_2012_),
    .X(_2013_));
 sky130_fd_sc_hd__mux2_1 _4920_ (.A0(\disp_song.um.drum.next_note2[28] ),
    .A1(\disp_song.um.drum.next_note2[29] ),
    .S(_1956_),
    .X(_2014_));
 sky130_fd_sc_hd__nand2_1 _4921_ (.A(_1968_),
    .B(_2014_),
    .Y(_2015_));
 sky130_fd_sc_hd__nor2_1 _4922_ (.A(_2669_),
    .B(_1992_),
    .Y(_2016_));
 sky130_fd_sc_hd__a32o_1 _4923_ (.A1(_1956_),
    .A2(\disp_song.um.drum.next_note2[31] ),
    .A3(_1965_),
    .B1(_2016_),
    .B2(\disp_song.um.drum.next_note2[30] ),
    .X(_2017_));
 sky130_fd_sc_hd__inv_2 _4924_ (.A(_2017_),
    .Y(_2018_));
 sky130_fd_sc_hd__nand2_2 _4925_ (.A(_2667_),
    .B(_2670_),
    .Y(_2019_));
 sky130_fd_sc_hd__nand2_4 _4926_ (.A(_2009_),
    .B(_2019_),
    .Y(_2020_));
 sky130_fd_sc_hd__mux2_1 _4927_ (.A0(_2015_),
    .A1(_2018_),
    .S(_2020_),
    .X(_2021_));
 sky130_fd_sc_hd__nor2_1 _4928_ (.A(_2013_),
    .B(_2021_),
    .Y(_2022_));
 sky130_fd_sc_hd__or2_1 _4929_ (.A(_1956_),
    .B(\disp_song.um.drum.next_note2[26] ),
    .X(_2023_));
 sky130_fd_sc_hd__nand2_1 _4930_ (.A(_1956_),
    .B(_0343_),
    .Y(_2024_));
 sky130_fd_sc_hd__and2_1 _4931_ (.A(_2009_),
    .B(_2019_),
    .X(_2025_));
 sky130_fd_sc_hd__clkbuf_4 _4932_ (.A(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__a31o_1 _4933_ (.A1(_1965_),
    .A2(_2023_),
    .A3(_2024_),
    .B1(_2026_),
    .X(_2027_));
 sky130_fd_sc_hd__or2_1 _4934_ (.A(\disp_song.note2[24] ),
    .B(_1956_),
    .X(_2028_));
 sky130_fd_sc_hd__or2_1 _4935_ (.A(_1949_),
    .B(_2010_),
    .X(_2029_));
 sky130_fd_sc_hd__a21o_1 _4936_ (.A1(\disp_song.um.drum.next_note2[25] ),
    .A2(_2029_),
    .B1(_2666_),
    .X(_2030_));
 sky130_fd_sc_hd__a21o_1 _4937_ (.A1(_2028_),
    .A2(_2030_),
    .B1(_2020_),
    .X(_2031_));
 sky130_fd_sc_hd__xnor2_1 _4938_ (.A(_2679_),
    .B(_2010_),
    .Y(_2032_));
 sky130_fd_sc_hd__a31o_1 _4939_ (.A1(_2013_),
    .A2(_2027_),
    .A3(_2031_),
    .B1(_2032_),
    .X(_2033_));
 sky130_fd_sc_hd__nor2_2 _4940_ (.A(_2010_),
    .B(_2012_),
    .Y(_2034_));
 sky130_fd_sc_hd__nor2_2 _4941_ (.A(_2666_),
    .B(_2669_),
    .Y(_2035_));
 sky130_fd_sc_hd__or2_1 _4942_ (.A(_2035_),
    .B(_2016_),
    .X(_2036_));
 sky130_fd_sc_hd__a32o_1 _4943_ (.A1(_1956_),
    .A2(\disp_song.um.drum.next_note2[23] ),
    .A3(_1968_),
    .B1(_2036_),
    .B2(\disp_song.um.drum.next_note2[22] ),
    .X(_2037_));
 sky130_fd_sc_hd__and3_1 _4944_ (.A(_2677_),
    .B(_0162_),
    .C(_2012_),
    .X(_2038_));
 sky130_fd_sc_hd__nand2_1 _4945_ (.A(_1956_),
    .B(\disp_song.um.drum.next_note2[21] ),
    .Y(_2039_));
 sky130_fd_sc_hd__a2bb2o_1 _4946_ (.A1_N(_2038_),
    .A2_N(_2039_),
    .B1(\disp_song.note2[20] ),
    .B2(\disp_song.um.drum.next_idx2[0] ),
    .X(_2040_));
 sky130_fd_sc_hd__mux2_1 _4947_ (.A0(_2037_),
    .A1(_2040_),
    .S(_2026_),
    .X(_2041_));
 sky130_fd_sc_hd__nor2_1 _4948_ (.A(_2667_),
    .B(_2669_),
    .Y(_2042_));
 sky130_fd_sc_hd__nand2_4 _4949_ (.A(_1992_),
    .B(_2042_),
    .Y(_2043_));
 sky130_fd_sc_hd__or2_1 _4950_ (.A(\disp_song.note2[17] ),
    .B(_2670_),
    .X(_2044_));
 sky130_fd_sc_hd__o211a_1 _4951_ (.A1(_1956_),
    .A2(\disp_song.um.drum.next_note2[16] ),
    .B1(_2043_),
    .C1(_2044_),
    .X(_2045_));
 sky130_fd_sc_hd__or2_1 _4952_ (.A(\disp_song.um.drum.next_idx2[0] ),
    .B(\disp_song.um.drum.next_note2[19] ),
    .X(_2046_));
 sky130_fd_sc_hd__or2_1 _4953_ (.A(_2669_),
    .B(\disp_song.um.drum.next_note2[18] ),
    .X(_2047_));
 sky130_fd_sc_hd__a31o_1 _4954_ (.A1(_1965_),
    .A2(_2046_),
    .A3(_2047_),
    .B1(_2026_),
    .X(_2048_));
 sky130_fd_sc_hd__o211a_1 _4955_ (.A1(_2020_),
    .A2(_2045_),
    .B1(_2048_),
    .C1(_2013_),
    .X(_2049_));
 sky130_fd_sc_hd__a21oi_1 _4956_ (.A1(_2034_),
    .A2(_2041_),
    .B1(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__a2bb2o_1 _4957_ (.A1_N(_2022_),
    .A2_N(_2033_),
    .B1(_2050_),
    .B2(_2032_),
    .X(_2051_));
 sky130_fd_sc_hd__a21oi_1 _4958_ (.A1(\disp_song.um.drum.next_note2[9] ),
    .A2(_2029_),
    .B1(_2666_),
    .Y(_2052_));
 sky130_fd_sc_hd__nor2_1 _4959_ (.A(\disp_song.note2[8] ),
    .B(_1956_),
    .Y(_2053_));
 sky130_fd_sc_hd__mux2_1 _4960_ (.A0(\disp_song.um.drum.next_note2[10] ),
    .A1(\disp_song.um.drum.next_note2[11] ),
    .S(_1956_),
    .X(_2054_));
 sky130_fd_sc_hd__nand2_1 _4961_ (.A(_2020_),
    .B(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__o32a_1 _4962_ (.A1(_2020_),
    .A2(_2052_),
    .A3(_2053_),
    .B1(_2055_),
    .B2(_1950_),
    .X(_2056_));
 sky130_fd_sc_hd__inv_2 _4963_ (.A(_2056_),
    .Y(_2057_));
 sky130_fd_sc_hd__or2_1 _4964_ (.A(\disp_song.um.drum.next_idx2[0] ),
    .B(\disp_song.um.drum.next_note2[13] ),
    .X(_2058_));
 sky130_fd_sc_hd__o211a_1 _4965_ (.A1(_1956_),
    .A2(\disp_song.um.drum.next_note2[12] ),
    .B1(_1968_),
    .C1(_2058_),
    .X(_2059_));
 sky130_fd_sc_hd__a32o_1 _4966_ (.A1(_1956_),
    .A2(\disp_song.um.drum.next_note2[15] ),
    .A3(_1965_),
    .B1(_2016_),
    .B2(\disp_song.um.drum.next_note2[14] ),
    .X(_2060_));
 sky130_fd_sc_hd__mux2_1 _4967_ (.A0(_2059_),
    .A1(_2060_),
    .S(_2020_),
    .X(_2061_));
 sky130_fd_sc_hd__mux2_1 _4968_ (.A0(_2057_),
    .A1(_2061_),
    .S(_2034_),
    .X(_2062_));
 sky130_fd_sc_hd__mux2_1 _4969_ (.A0(\disp_song.note2[1] ),
    .A1(\disp_song.um.drum.next_note2[0] ),
    .S(\disp_song.um.drum.next_idx2[0] ),
    .X(_2063_));
 sky130_fd_sc_hd__or2_1 _4970_ (.A(_2669_),
    .B(\disp_song.um.drum.next_note2[2] ),
    .X(_2064_));
 sky130_fd_sc_hd__o2111a_1 _4971_ (.A1(\disp_song.um.drum.next_idx2[0] ),
    .A2(\disp_song.um.drum.next_note2[3] ),
    .B1(_1965_),
    .C1(_2020_),
    .D1(_2064_),
    .X(_2065_));
 sky130_fd_sc_hd__a31o_1 _4972_ (.A1(_2026_),
    .A2(_2043_),
    .A3(_2063_),
    .B1(_2065_),
    .X(_2066_));
 sky130_fd_sc_hd__a32o_1 _4973_ (.A1(_1956_),
    .A2(\disp_song.um.drum.next_note2[7] ),
    .A3(_1968_),
    .B1(_2036_),
    .B2(\disp_song.um.drum.next_note2[6] ),
    .X(_2067_));
 sky130_fd_sc_hd__nand2_1 _4974_ (.A(_1956_),
    .B(\disp_song.um.drum.next_note2[5] ),
    .Y(_2068_));
 sky130_fd_sc_hd__a2bb2o_1 _4975_ (.A1_N(_2038_),
    .A2_N(_2068_),
    .B1(\disp_song.note2[4] ),
    .B2(\disp_song.um.drum.next_idx2[0] ),
    .X(_2069_));
 sky130_fd_sc_hd__mux2_1 _4976_ (.A0(_2067_),
    .A1(_2069_),
    .S(_2026_),
    .X(_2070_));
 sky130_fd_sc_hd__mux2_1 _4977_ (.A0(_2066_),
    .A1(_2070_),
    .S(_2034_),
    .X(_2071_));
 sky130_fd_sc_hd__mux2_1 _4978_ (.A0(_2062_),
    .A1(_2071_),
    .S(_2032_),
    .X(_2072_));
 sky130_fd_sc_hd__nor2_1 _4979_ (.A(_2011_),
    .B(_2072_),
    .Y(_2073_));
 sky130_fd_sc_hd__a211oi_1 _4980_ (.A1(_2011_),
    .A2(_2051_),
    .B1(_2073_),
    .C1(_0352_),
    .Y(\disp_song.um.drum.next_d2[1] ));
 sky130_fd_sc_hd__mux2_1 _4981_ (.A0(_1955_),
    .A1(_1958_),
    .S(_2666_),
    .X(_2074_));
 sky130_fd_sc_hd__inv_2 _4982_ (.A(_1973_),
    .Y(_2075_));
 sky130_fd_sc_hd__or2_1 _4983_ (.A(_1992_),
    .B(_1976_),
    .X(_2076_));
 sky130_fd_sc_hd__mux2_1 _4984_ (.A0(_2075_),
    .A1(_2076_),
    .S(_2667_),
    .X(_2077_));
 sky130_fd_sc_hd__or3_1 _4985_ (.A(\disp_song.um.drum.next_idx2[2] ),
    .B(_1962_),
    .C(_2077_),
    .X(_2078_));
 sky130_fd_sc_hd__o21ai_1 _4986_ (.A1(_0169_),
    .A2(_2074_),
    .B1(_2078_),
    .Y(_2079_));
 sky130_fd_sc_hd__mux2_1 _4987_ (.A0(_1986_),
    .A1(_1988_),
    .S(_2666_),
    .X(_2080_));
 sky130_fd_sc_hd__nand2_1 _4988_ (.A(_1968_),
    .B(_1991_),
    .Y(_2081_));
 sky130_fd_sc_hd__mux2_1 _4989_ (.A0(_1994_),
    .A1(_2081_),
    .S(_2667_),
    .X(_2082_));
 sky130_fd_sc_hd__or3_1 _4990_ (.A(\disp_song.um.drum.next_idx2[2] ),
    .B(_1962_),
    .C(_2082_),
    .X(_2083_));
 sky130_fd_sc_hd__o21ai_1 _4991_ (.A1(_0169_),
    .A2(_2080_),
    .B1(_2083_),
    .Y(_2084_));
 sky130_fd_sc_hd__and2_1 _4992_ (.A(_2677_),
    .B(_0169_),
    .X(_2085_));
 sky130_fd_sc_hd__or2_1 _4993_ (.A(_0162_),
    .B(_2085_),
    .X(_2086_));
 sky130_fd_sc_hd__mux2_1 _4994_ (.A0(_2079_),
    .A1(_2084_),
    .S(_2086_),
    .X(_2087_));
 sky130_fd_sc_hd__nand2_1 _4995_ (.A(_2666_),
    .B(_1969_),
    .Y(_2088_));
 sky130_fd_sc_hd__inv_2 _4996_ (.A(_2088_),
    .Y(_2089_));
 sky130_fd_sc_hd__a31o_1 _4997_ (.A1(\disp_song.um.drum.next_idx2[1] ),
    .A2(_1965_),
    .A3(_1966_),
    .B1(_2089_),
    .X(_2090_));
 sky130_fd_sc_hd__mux2_1 _4998_ (.A0(_1978_),
    .A1(_1979_),
    .S(_2666_),
    .X(_2091_));
 sky130_fd_sc_hd__mux2_1 _4999_ (.A0(_2090_),
    .A1(_2091_),
    .S(_0169_),
    .X(_2092_));
 sky130_fd_sc_hd__mux2_1 _5000_ (.A0(_1999_),
    .A1(_2001_),
    .S(_2667_),
    .X(_2093_));
 sky130_fd_sc_hd__mux2_1 _5001_ (.A0(_2003_),
    .A1(_2004_),
    .S(_2666_),
    .X(_2094_));
 sky130_fd_sc_hd__mux2_1 _5002_ (.A0(_2093_),
    .A1(_2094_),
    .S(_0169_),
    .X(_2095_));
 sky130_fd_sc_hd__mux2_1 _5003_ (.A0(_2092_),
    .A1(_2095_),
    .S(_2086_),
    .X(_2096_));
 sky130_fd_sc_hd__nor2_1 _5004_ (.A(_1960_),
    .B(_2085_),
    .Y(_2097_));
 sky130_fd_sc_hd__mux2_1 _5005_ (.A0(_2087_),
    .A1(_2096_),
    .S(_2097_),
    .X(_2098_));
 sky130_fd_sc_hd__and2_1 _5006_ (.A(_0214_),
    .B(_2098_),
    .X(_2099_));
 sky130_fd_sc_hd__clkbuf_1 _5007_ (.A(_2099_),
    .X(\disp_song.um.drum.next_d2[2] ));
 sky130_fd_sc_hd__xnor2_2 _5008_ (.A(\disp_song.um.drum.next_idx2[2] ),
    .B(_2035_),
    .Y(_2100_));
 sky130_fd_sc_hd__mux2_1 _5009_ (.A0(_2059_),
    .A1(_2060_),
    .S(_2026_),
    .X(_2101_));
 sky130_fd_sc_hd__a21oi_1 _5010_ (.A1(\disp_song.um.drum.next_note2[9] ),
    .A2(_1968_),
    .B1(\disp_song.um.drum.next_idx2[1] ),
    .Y(_2102_));
 sky130_fd_sc_hd__nor2_1 _5011_ (.A(_2053_),
    .B(_2102_),
    .Y(_2103_));
 sky130_fd_sc_hd__o211a_1 _5012_ (.A1(\disp_song.um.drum.next_idx2[0] ),
    .A2(_1965_),
    .B1(_2054_),
    .C1(_2043_),
    .X(_2104_));
 sky130_fd_sc_hd__inv_2 _5013_ (.A(_2100_),
    .Y(_2105_));
 sky130_fd_sc_hd__o221a_1 _5014_ (.A1(_2042_),
    .A2(_2103_),
    .B1(_2104_),
    .B2(_2020_),
    .C1(_2105_),
    .X(_2106_));
 sky130_fd_sc_hd__and2_1 _5015_ (.A(_2019_),
    .B(_2085_),
    .X(_2107_));
 sky130_fd_sc_hd__nor2_1 _5016_ (.A(_0162_),
    .B(_2107_),
    .Y(_2108_));
 sky130_fd_sc_hd__a211o_1 _5017_ (.A1(_2100_),
    .A2(_2101_),
    .B1(_2106_),
    .C1(_2108_),
    .X(_2109_));
 sky130_fd_sc_hd__or2_1 _5018_ (.A(_0162_),
    .B(_2107_),
    .X(_2110_));
 sky130_fd_sc_hd__o211a_1 _5019_ (.A1(_1968_),
    .A2(_2035_),
    .B1(_2023_),
    .C1(_2024_),
    .X(_2111_));
 sky130_fd_sc_hd__a21o_1 _5020_ (.A1(\disp_song.um.drum.next_note2[25] ),
    .A2(_1968_),
    .B1(_2667_),
    .X(_2112_));
 sky130_fd_sc_hd__a21o_1 _5021_ (.A1(_2028_),
    .A2(_2112_),
    .B1(_2042_),
    .X(_2113_));
 sky130_fd_sc_hd__o211a_1 _5022_ (.A1(_2020_),
    .A2(_2111_),
    .B1(_2105_),
    .C1(_2113_),
    .X(_2114_));
 sky130_fd_sc_hd__nand2_1 _5023_ (.A(_2020_),
    .B(_2015_),
    .Y(_2115_));
 sky130_fd_sc_hd__o211a_1 _5024_ (.A1(_2020_),
    .A2(_2017_),
    .B1(_2100_),
    .C1(_2115_),
    .X(_2116_));
 sky130_fd_sc_hd__a21oi_1 _5025_ (.A1(_0169_),
    .A2(_2019_),
    .B1(_2679_),
    .Y(_2117_));
 sky130_fd_sc_hd__o32a_1 _5026_ (.A1(_2110_),
    .A2(_2114_),
    .A3(_2116_),
    .B1(_2117_),
    .B2(_2107_),
    .X(_2118_));
 sky130_fd_sc_hd__o211a_1 _5027_ (.A1(\disp_song.note2[3] ),
    .A2(\disp_song.um.drum.next_idx2[0] ),
    .B1(_2043_),
    .C1(_2064_),
    .X(_2119_));
 sky130_fd_sc_hd__mux2_1 _5028_ (.A0(_2067_),
    .A1(_2119_),
    .S(\disp_song.um.drum.next_idx2[2] ),
    .X(_2120_));
 sky130_fd_sc_hd__o211a_1 _5029_ (.A1(\disp_song.note2[19] ),
    .A2(\disp_song.um.drum.next_idx2[0] ),
    .B1(_2047_),
    .C1(_2043_),
    .X(_2121_));
 sky130_fd_sc_hd__mux2_1 _5030_ (.A0(_2037_),
    .A1(_2121_),
    .S(\disp_song.um.drum.next_idx2[2] ),
    .X(_2122_));
 sky130_fd_sc_hd__mux2_1 _5031_ (.A0(_2120_),
    .A1(_2122_),
    .S(_2108_),
    .X(_2123_));
 sky130_fd_sc_hd__mux2_1 _5032_ (.A0(_2040_),
    .A1(_2069_),
    .S(_2110_),
    .X(_2124_));
 sky130_fd_sc_hd__or2_1 _5033_ (.A(_2045_),
    .B(_2110_),
    .X(_2125_));
 sky130_fd_sc_hd__nand2_1 _5034_ (.A(_2043_),
    .B(_2063_),
    .Y(_2126_));
 sky130_fd_sc_hd__a21oi_1 _5035_ (.A1(_2126_),
    .A2(_2110_),
    .B1(_2100_),
    .Y(_2127_));
 sky130_fd_sc_hd__a221o_1 _5036_ (.A1(_2100_),
    .A2(_2124_),
    .B1(_2125_),
    .B2(_2127_),
    .C1(_2026_),
    .X(_2128_));
 sky130_fd_sc_hd__nor2_1 _5037_ (.A(_2107_),
    .B(_2117_),
    .Y(_2129_));
 sky130_fd_sc_hd__o211a_1 _5038_ (.A1(_2020_),
    .A2(_2123_),
    .B1(_2128_),
    .C1(_2129_),
    .X(_2130_));
 sky130_fd_sc_hd__a211o_1 _5039_ (.A1(_2109_),
    .A2(_2118_),
    .B1(_2130_),
    .C1(_1950_),
    .X(_2131_));
 sky130_fd_sc_hd__or2_1 _5040_ (.A(_0169_),
    .B(_1949_),
    .X(_2132_));
 sky130_fd_sc_hd__or3_1 _5041_ (.A(\disp_song.um.drum.next_idx2[1] ),
    .B(_1956_),
    .C(_2132_),
    .X(_2133_));
 sky130_fd_sc_hd__inv_2 _5042_ (.A(_2133_),
    .Y(_2134_));
 sky130_fd_sc_hd__nor2_1 _5043_ (.A(_2009_),
    .B(_2132_),
    .Y(_2135_));
 sky130_fd_sc_hd__a32o_1 _5044_ (.A1(\disp_song.um.drum.next_note2[0] ),
    .A2(_1992_),
    .A3(_2035_),
    .B1(_2135_),
    .B2(\disp_song.um.drum.next_note2[1] ),
    .X(_2136_));
 sky130_fd_sc_hd__a211o_1 _5045_ (.A1(\disp_song.um.drum.next_note2[2] ),
    .A2(_2134_),
    .B1(_2136_),
    .C1(_1965_),
    .X(_2137_));
 sky130_fd_sc_hd__and3_1 _5046_ (.A(_0214_),
    .B(_2131_),
    .C(_2137_),
    .X(_2138_));
 sky130_fd_sc_hd__clkbuf_1 _5047_ (.A(_2138_),
    .X(\disp_song.um.drum.next_d2[3] ));
 sky130_fd_sc_hd__and3_1 _5048_ (.A(_2666_),
    .B(_1968_),
    .C(_1966_),
    .X(_2139_));
 sky130_fd_sc_hd__a21oi_1 _5049_ (.A1(\disp_song.um.drum.next_idx2[1] ),
    .A2(_1969_),
    .B1(_2139_),
    .Y(_2140_));
 sky130_fd_sc_hd__o2bb2a_2 _5050_ (.A1_N(_2666_),
    .A2_N(_2085_),
    .B1(_1982_),
    .B2(_2679_),
    .X(_2141_));
 sky130_fd_sc_hd__mux2_1 _5051_ (.A0(_1959_),
    .A1(_2140_),
    .S(_2141_),
    .X(_2142_));
 sky130_fd_sc_hd__a21oi_1 _5052_ (.A1(_1980_),
    .A2(_2141_),
    .B1(_1983_),
    .Y(_2143_));
 sky130_fd_sc_hd__nor2_1 _5053_ (.A(_2666_),
    .B(_1973_),
    .Y(_2144_));
 sky130_fd_sc_hd__a211o_1 _5054_ (.A1(_2666_),
    .A2(_2076_),
    .B1(_2141_),
    .C1(_2144_),
    .X(_2145_));
 sky130_fd_sc_hd__a22o_1 _5055_ (.A1(_1983_),
    .A2(_2142_),
    .B1(_2143_),
    .B2(_2145_),
    .X(_2146_));
 sky130_fd_sc_hd__o21a_1 _5056_ (.A1(\disp_song.um.drum.next_idx2[1] ),
    .A2(_2081_),
    .B1(_1995_),
    .X(_2147_));
 sky130_fd_sc_hd__mux2_1 _5057_ (.A0(_2147_),
    .A1(_1989_),
    .S(_1983_),
    .X(_2148_));
 sky130_fd_sc_hd__inv_2 _5058_ (.A(_2001_),
    .Y(_2149_));
 sky130_fd_sc_hd__o311a_1 _5059_ (.A1(\disp_song.um.drum.next_idx2[1] ),
    .A2(_1992_),
    .A3(_2149_),
    .B1(_2000_),
    .C1(_1983_),
    .X(_2150_));
 sky130_fd_sc_hd__o21ai_1 _5060_ (.A1(_1983_),
    .A2(_2005_),
    .B1(_2141_),
    .Y(_2151_));
 sky130_fd_sc_hd__o22a_1 _5061_ (.A1(_2141_),
    .A2(_2148_),
    .B1(_2150_),
    .B2(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__a21o_1 _5062_ (.A1(_2666_),
    .A2(_2085_),
    .B1(_0162_),
    .X(_2153_));
 sky130_fd_sc_hd__mux2_1 _5063_ (.A0(_2146_),
    .A1(_2152_),
    .S(_2153_),
    .X(_2154_));
 sky130_fd_sc_hd__nor2_1 _5064_ (.A(_0352_),
    .B(_2154_),
    .Y(\disp_song.um.drum.next_d2[4] ));
 sky130_fd_sc_hd__a21oi_1 _5065_ (.A1(_2679_),
    .A2(_2012_),
    .B1(_0162_),
    .Y(_2155_));
 sky130_fd_sc_hd__inv_2 _5066_ (.A(_2155_),
    .Y(_2156_));
 sky130_fd_sc_hd__xnor2_2 _5067_ (.A(_2679_),
    .B(_2012_),
    .Y(_2157_));
 sky130_fd_sc_hd__o21a_1 _5068_ (.A1(\disp_song.note2[16] ),
    .A2(\disp_song.um.drum.next_idx2[1] ),
    .B1(_2044_),
    .X(_2158_));
 sky130_fd_sc_hd__mux2_1 _5069_ (.A0(_2121_),
    .A1(_2158_),
    .S(_2026_),
    .X(_2159_));
 sky130_fd_sc_hd__mux2_1 _5070_ (.A0(_2041_),
    .A1(_2159_),
    .S(_2034_),
    .X(_2160_));
 sky130_fd_sc_hd__o211a_1 _5071_ (.A1(_2026_),
    .A2(_2111_),
    .B1(_2031_),
    .C1(_2034_),
    .X(_2161_));
 sky130_fd_sc_hd__o21ai_1 _5072_ (.A1(_2034_),
    .A2(_2021_),
    .B1(_2157_),
    .Y(_2162_));
 sky130_fd_sc_hd__o22a_1 _5073_ (.A1(_2157_),
    .A2(_2160_),
    .B1(_2161_),
    .B2(_2162_),
    .X(_2163_));
 sky130_fd_sc_hd__nor2_1 _5074_ (.A(_2034_),
    .B(_2070_),
    .Y(_2164_));
 sky130_fd_sc_hd__o22a_1 _5075_ (.A1(\disp_song.note2[0] ),
    .A2(\disp_song.um.drum.next_idx2[1] ),
    .B1(\disp_song.um.drum.next_idx2[0] ),
    .B2(\disp_song.note2[1] ),
    .X(_2165_));
 sky130_fd_sc_hd__mux2_1 _5076_ (.A0(_2119_),
    .A1(_2165_),
    .S(_2026_),
    .X(_2166_));
 sky130_fd_sc_hd__nor2_1 _5077_ (.A(_2013_),
    .B(_2166_),
    .Y(_2167_));
 sky130_fd_sc_hd__mux2_1 _5078_ (.A0(_2057_),
    .A1(_2061_),
    .S(_2013_),
    .X(_2168_));
 sky130_fd_sc_hd__a21oi_1 _5079_ (.A1(_2157_),
    .A2(_2168_),
    .B1(_2155_),
    .Y(_2169_));
 sky130_fd_sc_hd__o31ai_1 _5080_ (.A1(_2157_),
    .A2(_2164_),
    .A3(_2167_),
    .B1(_2169_),
    .Y(_2170_));
 sky130_fd_sc_hd__o211a_1 _5081_ (.A1(_2156_),
    .A2(_2163_),
    .B1(_2170_),
    .C1(_0214_),
    .X(\disp_song.um.drum.next_d2[5] ));
 sky130_fd_sc_hd__inv_2 _5082_ (.A(_2043_),
    .Y(_2171_));
 sky130_fd_sc_hd__a32o_1 _5083_ (.A1(\disp_song.um.drum.next_note2[3] ),
    .A2(_1992_),
    .A3(_2035_),
    .B1(_2171_),
    .B2(\disp_song.um.drum.next_note2[1] ),
    .X(_2172_));
 sky130_fd_sc_hd__a221o_1 _5084_ (.A1(\disp_song.um.drum.next_note2[5] ),
    .A2(_2134_),
    .B1(_2135_),
    .B2(\disp_song.um.drum.next_note2[4] ),
    .C1(_2172_),
    .X(_2173_));
 sky130_fd_sc_hd__and4b_1 _5085_ (.A_N(_2664_),
    .B(_1956_),
    .C(\disp_song.um.drum.next_note2[2] ),
    .D(_1992_),
    .X(_2174_));
 sky130_fd_sc_hd__a211o_1 _5086_ (.A1(\disp_song.um.drum.next_note2[0] ),
    .A2(_2038_),
    .B1(_2174_),
    .C1(_1965_),
    .X(_2175_));
 sky130_fd_sc_hd__mux2_1 _5087_ (.A0(_2093_),
    .A1(_2094_),
    .S(\disp_song.um.drum.next_idx2[2] ),
    .X(_2176_));
 sky130_fd_sc_hd__a21o_1 _5088_ (.A1(\disp_song.um.drum.next_idx2[1] ),
    .A2(_1966_),
    .B1(_2089_),
    .X(_2177_));
 sky130_fd_sc_hd__mux2_1 _5089_ (.A0(_2091_),
    .A1(_2177_),
    .S(_0169_),
    .X(_2178_));
 sky130_fd_sc_hd__mux2_1 _5090_ (.A0(_2176_),
    .A1(_2178_),
    .S(\disp_song.um.drum.next_idx2[4] ),
    .X(_2179_));
 sky130_fd_sc_hd__mux2_1 _5091_ (.A0(_2074_),
    .A1(_2077_),
    .S(\disp_song.um.drum.next_idx2[2] ),
    .X(_2180_));
 sky130_fd_sc_hd__mux2_1 _5092_ (.A0(_2082_),
    .A1(_2080_),
    .S(_0169_),
    .X(_2181_));
 sky130_fd_sc_hd__mux2_1 _5093_ (.A0(_2180_),
    .A1(_2181_),
    .S(_0162_),
    .X(_2182_));
 sky130_fd_sc_hd__nor2_1 _5094_ (.A(_2677_),
    .B(_2182_),
    .Y(_2183_));
 sky130_fd_sc_hd__a211o_1 _5095_ (.A1(_2677_),
    .A2(_2179_),
    .B1(_2183_),
    .C1(_1950_),
    .X(_2184_));
 sky130_fd_sc_hd__o211a_1 _5096_ (.A1(_2173_),
    .A2(_2175_),
    .B1(_0214_),
    .C1(_2184_),
    .X(\disp_song.um.drum.next_d2[6] ));
 sky130_fd_sc_hd__buf_6 _5097_ (.A(_0199_),
    .X(_2185_));
 sky130_fd_sc_hd__nand2_1 _5098_ (.A(\disp_song.um.drum.next_idx1[2] ),
    .B(\disp_song.um.drum.next_idx1[3] ),
    .Y(_2186_));
 sky130_fd_sc_hd__nand2_2 _5099_ (.A(\disp_song.um.drum.next_idx1[2] ),
    .B(\disp_song.um.drum.next_idx1[1] ),
    .Y(_2187_));
 sky130_fd_sc_hd__a2bb2o_1 _5100_ (.A1_N(_2185_),
    .A2_N(_2186_),
    .B1(_2187_),
    .B2(_0197_),
    .X(_2188_));
 sky130_fd_sc_hd__inv_2 _5101_ (.A(_2188_),
    .Y(_2189_));
 sky130_fd_sc_hd__or3_1 _5102_ (.A(\disp_song.um.drum.next_idx1[4] ),
    .B(\disp_song.um.drum.next_idx1[2] ),
    .C(\disp_song.um.drum.next_idx1[3] ),
    .X(_2190_));
 sky130_fd_sc_hd__clkbuf_4 _5103_ (.A(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__mux2_1 _5104_ (.A0(\disp_song.um.drum.next_note1[12] ),
    .A1(\disp_song.um.drum.next_note1[13] ),
    .S(_0176_),
    .X(_2192_));
 sky130_fd_sc_hd__a21oi_1 _5105_ (.A1(_2191_),
    .A2(_2192_),
    .B1(\disp_song.um.drum.next_idx1[2] ),
    .Y(_2193_));
 sky130_fd_sc_hd__and2_1 _5106_ (.A(_0197_),
    .B(_2187_),
    .X(_2194_));
 sky130_fd_sc_hd__nand2_4 _5107_ (.A(_0185_),
    .B(_2194_),
    .Y(_2195_));
 sky130_fd_sc_hd__mux2_1 _5108_ (.A0(\disp_song.um.drum.next_note1[14] ),
    .A1(\disp_song.um.drum.next_note1[15] ),
    .S(\disp_song.um.drum.next_idx1[0] ),
    .X(_2196_));
 sky130_fd_sc_hd__a21oi_1 _5109_ (.A1(_2195_),
    .A2(_2196_),
    .B1(\disp_song.um.drum.next_idx1[1] ),
    .Y(_2197_));
 sky130_fd_sc_hd__nor2_1 _5110_ (.A(_2193_),
    .B(_2197_),
    .Y(_2198_));
 sky130_fd_sc_hd__mux2_1 _5111_ (.A0(\disp_song.um.drum.next_note1[6] ),
    .A1(\disp_song.um.drum.next_note1[7] ),
    .S(_0176_),
    .X(_2199_));
 sky130_fd_sc_hd__mux2_1 _5112_ (.A0(\disp_song.um.drum.next_note1[4] ),
    .A1(\disp_song.um.drum.next_note1[5] ),
    .S(_0176_),
    .X(_2200_));
 sky130_fd_sc_hd__mux2_1 _5113_ (.A0(_2199_),
    .A1(_2200_),
    .S(\disp_song.um.drum.next_idx1[1] ),
    .X(_2201_));
 sky130_fd_sc_hd__o22a_1 _5114_ (.A1(_2189_),
    .A2(_2198_),
    .B1(_2201_),
    .B2(_0197_),
    .X(_2202_));
 sky130_fd_sc_hd__mux2_1 _5115_ (.A0(\disp_song.um.drum.next_note1[10] ),
    .A1(\disp_song.um.drum.next_note1[11] ),
    .S(\disp_song.um.drum.next_idx1[0] ),
    .X(_2203_));
 sky130_fd_sc_hd__a21o_1 _5116_ (.A1(_2191_),
    .A2(_2203_),
    .B1(\disp_song.um.drum.next_idx1[1] ),
    .X(_2204_));
 sky130_fd_sc_hd__mux2_1 _5117_ (.A0(\disp_song.um.drum.next_note1[8] ),
    .A1(\disp_song.um.drum.next_note1[9] ),
    .S(_0176_),
    .X(_2205_));
 sky130_fd_sc_hd__or2_1 _5118_ (.A(_2185_),
    .B(_2205_),
    .X(_2206_));
 sky130_fd_sc_hd__and3_1 _5119_ (.A(_0185_),
    .B(_0191_),
    .C(_0197_),
    .X(_2207_));
 sky130_fd_sc_hd__clkbuf_2 _5120_ (.A(_2207_),
    .X(_2208_));
 sky130_fd_sc_hd__nor2_1 _5121_ (.A(_0373_),
    .B(_2208_),
    .Y(_2209_));
 sky130_fd_sc_hd__mux2_1 _5122_ (.A0(\disp_song.note1[2] ),
    .A1(_2209_),
    .S(\disp_song.um.drum.next_idx1[0] ),
    .X(_2210_));
 sky130_fd_sc_hd__mux2_1 _5123_ (.A0(\disp_song.um.drum.next_note1[0] ),
    .A1(\disp_song.um.drum.next_note1[1] ),
    .S(_0176_),
    .X(_2211_));
 sky130_fd_sc_hd__or2_1 _5124_ (.A(_2185_),
    .B(_2211_),
    .X(_2212_));
 sky130_fd_sc_hd__o211a_1 _5125_ (.A1(\disp_song.um.drum.next_idx1[1] ),
    .A2(_2210_),
    .B1(_2212_),
    .C1(_2189_),
    .X(_2213_));
 sky130_fd_sc_hd__a31o_1 _5126_ (.A1(_2188_),
    .A2(_2204_),
    .A3(_2206_),
    .B1(_2213_),
    .X(_2214_));
 sky130_fd_sc_hd__nand2_1 _5127_ (.A(_0191_),
    .B(_2185_),
    .Y(_2215_));
 sky130_fd_sc_hd__nand2_1 _5128_ (.A(_2187_),
    .B(_2215_),
    .Y(_2216_));
 sky130_fd_sc_hd__mux2_1 _5129_ (.A0(_2202_),
    .A1(_2214_),
    .S(_2216_),
    .X(_2217_));
 sky130_fd_sc_hd__mux2_1 _5130_ (.A0(\disp_song.um.drum.next_note1[22] ),
    .A1(\disp_song.um.drum.next_note1[23] ),
    .S(\disp_song.um.drum.next_idx1[0] ),
    .X(_2218_));
 sky130_fd_sc_hd__mux2_1 _5131_ (.A0(\disp_song.um.drum.next_note1[20] ),
    .A1(\disp_song.um.drum.next_note1[21] ),
    .S(\disp_song.um.drum.next_idx1[0] ),
    .X(_2219_));
 sky130_fd_sc_hd__mux2_1 _5132_ (.A0(_2218_),
    .A1(_2219_),
    .S(\disp_song.um.drum.next_idx1[1] ),
    .X(_2220_));
 sky130_fd_sc_hd__mux2_1 _5133_ (.A0(\disp_song.um.drum.next_note1[28] ),
    .A1(\disp_song.um.drum.next_note1[29] ),
    .S(\disp_song.um.drum.next_idx1[0] ),
    .X(_2221_));
 sky130_fd_sc_hd__a21oi_1 _5134_ (.A1(_2191_),
    .A2(_2221_),
    .B1(\disp_song.um.drum.next_idx1[2] ),
    .Y(_2222_));
 sky130_fd_sc_hd__mux2_1 _5135_ (.A0(\disp_song.um.drum.next_note1[30] ),
    .A1(\disp_song.um.drum.next_note1[31] ),
    .S(\disp_song.um.drum.next_idx1[0] ),
    .X(_2223_));
 sky130_fd_sc_hd__a21oi_1 _5136_ (.A1(_2195_),
    .A2(_2223_),
    .B1(\disp_song.um.drum.next_idx1[1] ),
    .Y(_2224_));
 sky130_fd_sc_hd__nor2_1 _5137_ (.A(_2222_),
    .B(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__nor2_1 _5138_ (.A(_0415_),
    .B(_2208_),
    .Y(_2226_));
 sky130_fd_sc_hd__mux2_1 _5139_ (.A0(\disp_song.note1[18] ),
    .A1(_2226_),
    .S(\disp_song.um.drum.next_idx1[0] ),
    .X(_2227_));
 sky130_fd_sc_hd__mux2_1 _5140_ (.A0(\disp_song.um.drum.next_note1[16] ),
    .A1(\disp_song.um.drum.next_note1[17] ),
    .S(\disp_song.um.drum.next_idx1[0] ),
    .X(_2228_));
 sky130_fd_sc_hd__mux2_1 _5141_ (.A0(_2227_),
    .A1(_2228_),
    .S(\disp_song.um.drum.next_idx1[1] ),
    .X(_2229_));
 sky130_fd_sc_hd__and2_1 _5142_ (.A(_0198_),
    .B(_2208_),
    .X(_2230_));
 sky130_fd_sc_hd__or2_1 _5143_ (.A(_0430_),
    .B(_2230_),
    .X(_2231_));
 sky130_fd_sc_hd__clkbuf_8 _5144_ (.A(_0175_),
    .X(_2232_));
 sky130_fd_sc_hd__nand2_1 _5145_ (.A(_2232_),
    .B(\disp_song.um.drum.next_note1[26] ),
    .Y(_2233_));
 sky130_fd_sc_hd__and3_1 _5146_ (.A(_0185_),
    .B(_0197_),
    .C(_2187_),
    .X(_2234_));
 sky130_fd_sc_hd__o221a_1 _5147_ (.A1(_0173_),
    .A2(_2231_),
    .B1(_2233_),
    .B2(_2234_),
    .C1(_2185_),
    .X(_2235_));
 sky130_fd_sc_hd__mux2_1 _5148_ (.A0(\disp_song.um.drum.next_note1[24] ),
    .A1(\disp_song.um.drum.next_note1[25] ),
    .S(\disp_song.um.drum.next_idx1[0] ),
    .X(_2236_));
 sky130_fd_sc_hd__nor2_1 _5149_ (.A(_2185_),
    .B(_2236_),
    .Y(_2237_));
 sky130_fd_sc_hd__nor2_1 _5150_ (.A(_2235_),
    .B(_2237_),
    .Y(_2238_));
 sky130_fd_sc_hd__mux4_1 _5151_ (.A0(_2220_),
    .A1(_2225_),
    .A2(_2229_),
    .A3(_2238_),
    .S0(_2188_),
    .S1(_2216_),
    .X(_2239_));
 sky130_fd_sc_hd__nor2_1 _5152_ (.A(_0185_),
    .B(_2194_),
    .Y(_2240_));
 sky130_fd_sc_hd__mux2_1 _5153_ (.A0(_2217_),
    .A1(_2239_),
    .S(_2240_),
    .X(_2241_));
 sky130_fd_sc_hd__and2_1 _5154_ (.A(_0214_),
    .B(_2241_),
    .X(_2242_));
 sky130_fd_sc_hd__clkbuf_1 _5155_ (.A(_2242_),
    .X(\disp_song.um.drum.next_d1[0] ));
 sky130_fd_sc_hd__and3_1 _5156_ (.A(_2654_),
    .B(_0173_),
    .C(_0198_),
    .X(_2243_));
 sky130_fd_sc_hd__buf_2 _5157_ (.A(_2243_),
    .X(_2244_));
 sky130_fd_sc_hd__nor2_1 _5158_ (.A(_0191_),
    .B(_2244_),
    .Y(_2245_));
 sky130_fd_sc_hd__and3_2 _5159_ (.A(_0175_),
    .B(_0191_),
    .C(_0198_),
    .X(_2246_));
 sky130_fd_sc_hd__or2_2 _5160_ (.A(_2245_),
    .B(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__or2_1 _5161_ (.A(_0176_),
    .B(\disp_song.um.drum.next_note1[29] ),
    .X(_2248_));
 sky130_fd_sc_hd__o211a_1 _5162_ (.A1(_0175_),
    .A2(\disp_song.um.drum.next_note1[28] ),
    .B1(_2191_),
    .C1(_2248_),
    .X(_2249_));
 sky130_fd_sc_hd__or2_1 _5163_ (.A(_0176_),
    .B(\disp_song.um.drum.next_note1[31] ),
    .X(_2250_));
 sky130_fd_sc_hd__o211a_1 _5164_ (.A1(_0175_),
    .A2(\disp_song.um.drum.next_note1[30] ),
    .B1(_2195_),
    .C1(_2250_),
    .X(_2251_));
 sky130_fd_sc_hd__nor2_4 _5165_ (.A(_0175_),
    .B(_2185_),
    .Y(_2252_));
 sky130_fd_sc_hd__or2_1 _5166_ (.A(_2244_),
    .B(_2252_),
    .X(_2253_));
 sky130_fd_sc_hd__buf_4 _5167_ (.A(_2253_),
    .X(_2254_));
 sky130_fd_sc_hd__mux2_1 _5168_ (.A0(_2249_),
    .A1(_2251_),
    .S(_2254_),
    .X(_2255_));
 sky130_fd_sc_hd__nor2_4 _5169_ (.A(_2244_),
    .B(_2252_),
    .Y(_2256_));
 sky130_fd_sc_hd__or2_1 _5170_ (.A(\disp_song.um.drum.next_idx1[3] ),
    .B(_2245_),
    .X(_2257_));
 sky130_fd_sc_hd__nor2_2 _5171_ (.A(\disp_song.um.drum.next_idx1[4] ),
    .B(_2257_),
    .Y(_2258_));
 sky130_fd_sc_hd__o21ai_1 _5172_ (.A1(_0430_),
    .A2(_2258_),
    .B1(_0175_),
    .Y(_2259_));
 sky130_fd_sc_hd__o21ai_1 _5173_ (.A1(\disp_song.note1[26] ),
    .A2(_2232_),
    .B1(_2259_),
    .Y(_2260_));
 sky130_fd_sc_hd__inv_2 _5174_ (.A(_2258_),
    .Y(_2261_));
 sky130_fd_sc_hd__a21oi_1 _5175_ (.A1(\disp_song.um.drum.next_note1[25] ),
    .A2(_2261_),
    .B1(_2185_),
    .Y(_2262_));
 sky130_fd_sc_hd__o21ai_1 _5176_ (.A1(\disp_song.note1[24] ),
    .A2(_2232_),
    .B1(_2256_),
    .Y(_2263_));
 sky130_fd_sc_hd__o221a_1 _5177_ (.A1(_2256_),
    .A2(_2260_),
    .B1(_2262_),
    .B2(_2263_),
    .C1(_2247_),
    .X(_2264_));
 sky130_fd_sc_hd__o21ba_1 _5178_ (.A1(_2247_),
    .A2(_2255_),
    .B1_N(_2264_),
    .X(_2265_));
 sky130_fd_sc_hd__nand2_1 _5179_ (.A(_0175_),
    .B(\disp_song.um.drum.next_note1[21] ),
    .Y(_2266_));
 sky130_fd_sc_hd__a2bb2o_1 _5180_ (.A1_N(_2230_),
    .A2_N(_2266_),
    .B1(\disp_song.note1[20] ),
    .B2(\disp_song.um.drum.next_idx1[0] ),
    .X(_2267_));
 sky130_fd_sc_hd__nor2_1 _5181_ (.A(_0175_),
    .B(_2230_),
    .Y(_2268_));
 sky130_fd_sc_hd__a32o_1 _5182_ (.A1(_0175_),
    .A2(\disp_song.um.drum.next_note1[23] ),
    .A3(_2191_),
    .B1(_2268_),
    .B2(\disp_song.um.drum.next_note1[22] ),
    .X(_2269_));
 sky130_fd_sc_hd__mux2_1 _5183_ (.A0(_2267_),
    .A1(_2269_),
    .S(_2254_),
    .X(_2270_));
 sky130_fd_sc_hd__or2_1 _5184_ (.A(_0175_),
    .B(\disp_song.um.drum.next_note1[16] ),
    .X(_2271_));
 sky130_fd_sc_hd__and2_1 _5185_ (.A(\disp_song.um.drum.next_note1[17] ),
    .B(_2191_),
    .X(_2272_));
 sky130_fd_sc_hd__or2_1 _5186_ (.A(_2268_),
    .B(_2272_),
    .X(_2273_));
 sky130_fd_sc_hd__nor2_2 _5187_ (.A(_2245_),
    .B(_2246_),
    .Y(_2274_));
 sky130_fd_sc_hd__a31o_1 _5188_ (.A1(_2256_),
    .A2(_2271_),
    .A3(_2273_),
    .B1(_2274_),
    .X(_2275_));
 sky130_fd_sc_hd__o21ai_1 _5189_ (.A1(_0415_),
    .A2(_2258_),
    .B1(_2232_),
    .Y(_2276_));
 sky130_fd_sc_hd__o21ai_1 _5190_ (.A1(\disp_song.note1[18] ),
    .A2(_2232_),
    .B1(_2276_),
    .Y(_2277_));
 sky130_fd_sc_hd__nor2_1 _5191_ (.A(_2256_),
    .B(_2277_),
    .Y(_2278_));
 sky130_fd_sc_hd__o22a_1 _5192_ (.A1(_2247_),
    .A2(_2270_),
    .B1(_2275_),
    .B2(_2278_),
    .X(_2279_));
 sky130_fd_sc_hd__o21a_1 _5193_ (.A1(_2186_),
    .A2(_2244_),
    .B1(_2257_),
    .X(_2280_));
 sky130_fd_sc_hd__mux2_1 _5194_ (.A0(_2265_),
    .A1(_2279_),
    .S(_2280_),
    .X(_2281_));
 sky130_fd_sc_hd__or2_1 _5195_ (.A(_0175_),
    .B(\disp_song.um.drum.next_note1[12] ),
    .X(_2282_));
 sky130_fd_sc_hd__o211a_1 _5196_ (.A1(\disp_song.um.drum.next_idx1[0] ),
    .A2(\disp_song.um.drum.next_note1[13] ),
    .B1(_2191_),
    .C1(_2282_),
    .X(_2283_));
 sky130_fd_sc_hd__or2_1 _5197_ (.A(_0176_),
    .B(\disp_song.um.drum.next_note1[15] ),
    .X(_2284_));
 sky130_fd_sc_hd__o211a_1 _5198_ (.A1(_2232_),
    .A2(\disp_song.um.drum.next_note1[14] ),
    .B1(_2195_),
    .C1(_2284_),
    .X(_2285_));
 sky130_fd_sc_hd__mux2_1 _5199_ (.A0(_2283_),
    .A1(_2285_),
    .S(_2254_),
    .X(_2286_));
 sky130_fd_sc_hd__a21o_1 _5200_ (.A1(\disp_song.um.drum.next_note1[11] ),
    .A2(_2261_),
    .B1(_0176_),
    .X(_2287_));
 sky130_fd_sc_hd__o21ai_1 _5201_ (.A1(\disp_song.note1[10] ),
    .A2(_2232_),
    .B1(_2287_),
    .Y(_2288_));
 sky130_fd_sc_hd__a21oi_1 _5202_ (.A1(\disp_song.um.drum.next_note1[9] ),
    .A2(_2261_),
    .B1(_2185_),
    .Y(_2289_));
 sky130_fd_sc_hd__or2_1 _5203_ (.A(\disp_song.note1[8] ),
    .B(_0175_),
    .X(_2290_));
 sky130_fd_sc_hd__nand2_1 _5204_ (.A(_2256_),
    .B(_2290_),
    .Y(_2291_));
 sky130_fd_sc_hd__o221a_1 _5205_ (.A1(_2256_),
    .A2(_2288_),
    .B1(_2289_),
    .B2(_2291_),
    .C1(_2247_),
    .X(_2292_));
 sky130_fd_sc_hd__o21ba_1 _5206_ (.A1(_2247_),
    .A2(_2286_),
    .B1_N(_2292_),
    .X(_2293_));
 sky130_fd_sc_hd__nand2_1 _5207_ (.A(_0175_),
    .B(\disp_song.um.drum.next_note1[5] ),
    .Y(_2294_));
 sky130_fd_sc_hd__a2bb2o_1 _5208_ (.A1_N(_2230_),
    .A2_N(_2294_),
    .B1(\disp_song.note1[4] ),
    .B2(\disp_song.um.drum.next_idx1[0] ),
    .X(_2295_));
 sky130_fd_sc_hd__a32o_1 _5209_ (.A1(_2232_),
    .A2(\disp_song.um.drum.next_note1[7] ),
    .A3(_2191_),
    .B1(_2268_),
    .B2(\disp_song.um.drum.next_note1[6] ),
    .X(_2296_));
 sky130_fd_sc_hd__mux2_1 _5210_ (.A0(_2295_),
    .A1(_2296_),
    .S(_2254_),
    .X(_2297_));
 sky130_fd_sc_hd__a21oi_1 _5211_ (.A1(\disp_song.um.drum.next_note1[1] ),
    .A2(_2191_),
    .B1(\disp_song.um.drum.next_idx1[0] ),
    .Y(_2298_));
 sky130_fd_sc_hd__nor2_1 _5212_ (.A(_2232_),
    .B(\disp_song.um.drum.next_note1[0] ),
    .Y(_2299_));
 sky130_fd_sc_hd__a211o_1 _5213_ (.A1(\disp_song.um.drum.next_idx1[0] ),
    .A2(_2230_),
    .B1(_2298_),
    .C1(_2299_),
    .X(_2300_));
 sky130_fd_sc_hd__o21ai_1 _5214_ (.A1(_2254_),
    .A2(_2300_),
    .B1(_2247_),
    .Y(_2301_));
 sky130_fd_sc_hd__o21ai_1 _5215_ (.A1(_0373_),
    .A2(_2258_),
    .B1(_2232_),
    .Y(_2302_));
 sky130_fd_sc_hd__o21ai_1 _5216_ (.A1(\disp_song.note1[2] ),
    .A2(_2232_),
    .B1(_2302_),
    .Y(_2303_));
 sky130_fd_sc_hd__nor2_1 _5217_ (.A(_2256_),
    .B(_2303_),
    .Y(_2304_));
 sky130_fd_sc_hd__o22a_1 _5218_ (.A1(_2247_),
    .A2(_2297_),
    .B1(_2301_),
    .B2(_2304_),
    .X(_2305_));
 sky130_fd_sc_hd__mux2_1 _5219_ (.A0(_2293_),
    .A1(_2305_),
    .S(_2280_),
    .X(_2306_));
 sky130_fd_sc_hd__nand2_1 _5220_ (.A(\disp_song.um.drum.next_idx1[4] ),
    .B(_2257_),
    .Y(_2307_));
 sky130_fd_sc_hd__mux2_1 _5221_ (.A0(_2281_),
    .A1(_2306_),
    .S(_2307_),
    .X(_2308_));
 sky130_fd_sc_hd__and2_1 _5222_ (.A(_0214_),
    .B(_2308_),
    .X(_2309_));
 sky130_fd_sc_hd__clkbuf_1 _5223_ (.A(_2309_),
    .X(\disp_song.um.drum.next_d1[1] ));
 sky130_fd_sc_hd__nor2_1 _5224_ (.A(_0173_),
    .B(\disp_song.um.drum.next_idx1[1] ),
    .Y(_2310_));
 sky130_fd_sc_hd__or4b_1 _5225_ (.A(\disp_song.um.drum.next_idx1[4] ),
    .B(_0191_),
    .C(\disp_song.um.drum.next_idx1[3] ),
    .D_N(_2310_),
    .X(_2311_));
 sky130_fd_sc_hd__inv_2 _5226_ (.A(_2311_),
    .Y(_2312_));
 sky130_fd_sc_hd__or4b_1 _5227_ (.A(\disp_song.um.drum.next_idx1[4] ),
    .B(_0191_),
    .C(\disp_song.um.drum.next_idx1[3] ),
    .D_N(_2244_),
    .X(_2313_));
 sky130_fd_sc_hd__inv_2 _5228_ (.A(_2313_),
    .Y(_2314_));
 sky130_fd_sc_hd__a22o_1 _5229_ (.A1(\disp_song.um.drum.next_note1[1] ),
    .A2(_2312_),
    .B1(_2314_),
    .B2(\disp_song.um.drum.next_note1[0] ),
    .X(_2315_));
 sky130_fd_sc_hd__o21ai_1 _5230_ (.A1(_2232_),
    .A2(_0430_),
    .B1(_2233_),
    .Y(_2316_));
 sky130_fd_sc_hd__mux2_1 _5231_ (.A0(_2236_),
    .A1(_2316_),
    .S(\disp_song.um.drum.next_idx1[1] ),
    .X(_2317_));
 sky130_fd_sc_hd__mux2_1 _5232_ (.A0(_2218_),
    .A1(_2219_),
    .S(_2185_),
    .X(_2318_));
 sky130_fd_sc_hd__o21a_1 _5233_ (.A1(\disp_song.um.drum.next_idx1[2] ),
    .A2(_2318_),
    .B1(\disp_song.um.drum.next_idx1[4] ),
    .X(_2319_));
 sky130_fd_sc_hd__mux2_1 _5234_ (.A0(_2227_),
    .A1(_2228_),
    .S(_2185_),
    .X(_2320_));
 sky130_fd_sc_hd__a21o_1 _5235_ (.A1(\disp_song.um.drum.next_idx1[2] ),
    .A2(_2320_),
    .B1(\disp_song.um.drum.next_idx1[3] ),
    .X(_2321_));
 sky130_fd_sc_hd__o311a_1 _5236_ (.A1(_0191_),
    .A2(_0197_),
    .A3(_2317_),
    .B1(_2319_),
    .C1(_2321_),
    .X(_2322_));
 sky130_fd_sc_hd__nand2_1 _5237_ (.A(_0191_),
    .B(_0197_),
    .Y(_2323_));
 sky130_fd_sc_hd__mux2_1 _5238_ (.A0(_2199_),
    .A1(_2200_),
    .S(_2185_),
    .X(_2324_));
 sky130_fd_sc_hd__mux2_1 _5239_ (.A0(_2203_),
    .A1(_2205_),
    .S(_2185_),
    .X(_2325_));
 sky130_fd_sc_hd__mux2_1 _5240_ (.A0(_2192_),
    .A1(_2196_),
    .S(\disp_song.um.drum.next_idx1[1] ),
    .X(_2326_));
 sky130_fd_sc_hd__mux2_1 _5241_ (.A0(_2210_),
    .A1(_2211_),
    .S(_2185_),
    .X(_2327_));
 sky130_fd_sc_hd__mux4_1 _5242_ (.A0(_2324_),
    .A1(_2325_),
    .A2(_2326_),
    .A3(_2327_),
    .S0(\disp_song.um.drum.next_idx1[2] ),
    .S1(_0197_),
    .X(_2328_));
 sky130_fd_sc_hd__a21boi_1 _5243_ (.A1(\disp_song.um.drum.next_idx1[4] ),
    .A2(_2323_),
    .B1_N(_2328_),
    .Y(_2329_));
 sky130_fd_sc_hd__or3_1 _5244_ (.A(_2234_),
    .B(_2322_),
    .C(_2329_),
    .X(_2330_));
 sky130_fd_sc_hd__o211a_1 _5245_ (.A1(_2195_),
    .A2(_2315_),
    .B1(_2330_),
    .C1(_0214_),
    .X(\disp_song.um.drum.next_d1[2] ));
 sky130_fd_sc_hd__and2_1 _5246_ (.A(\disp_song.um.drum.next_note1[1] ),
    .B(_2314_),
    .X(_2331_));
 sky130_fd_sc_hd__a32o_1 _5247_ (.A1(\disp_song.um.drum.next_note1[0] ),
    .A2(_2208_),
    .A3(_2252_),
    .B1(_2312_),
    .B2(\disp_song.um.drum.next_note1[2] ),
    .X(_2332_));
 sky130_fd_sc_hd__o21ai_1 _5248_ (.A1(_2252_),
    .A2(_2323_),
    .B1(\disp_song.um.drum.next_idx1[4] ),
    .Y(_2333_));
 sky130_fd_sc_hd__mux2_1 _5249_ (.A0(_2283_),
    .A1(_2285_),
    .S(_2256_),
    .X(_2334_));
 sky130_fd_sc_hd__inv_2 _5250_ (.A(_2288_),
    .Y(_2335_));
 sky130_fd_sc_hd__nand2_1 _5251_ (.A(_2208_),
    .B(_2244_),
    .Y(_2336_));
 sky130_fd_sc_hd__o211a_1 _5252_ (.A1(\disp_song.um.drum.next_idx1[0] ),
    .A2(\disp_song.um.drum.next_note1[9] ),
    .B1(_2290_),
    .C1(_2336_),
    .X(_2337_));
 sky130_fd_sc_hd__mux2_1 _5253_ (.A0(_2335_),
    .A1(_2337_),
    .S(_2254_),
    .X(_2338_));
 sky130_fd_sc_hd__o22a_2 _5254_ (.A1(_0175_),
    .A2(_2187_),
    .B1(_2252_),
    .B2(\disp_song.um.drum.next_idx1[2] ),
    .X(_2339_));
 sky130_fd_sc_hd__mux2_1 _5255_ (.A0(_2334_),
    .A1(_2338_),
    .S(_2339_),
    .X(_2340_));
 sky130_fd_sc_hd__mux2_1 _5256_ (.A0(_2295_),
    .A1(_2296_),
    .S(_2256_),
    .X(_2341_));
 sky130_fd_sc_hd__nor2_1 _5257_ (.A(_2254_),
    .B(_2303_),
    .Y(_2342_));
 sky130_fd_sc_hd__o21ai_1 _5258_ (.A1(_2256_),
    .A2(_2300_),
    .B1(_2339_),
    .Y(_2343_));
 sky130_fd_sc_hd__o22a_1 _5259_ (.A1(_2339_),
    .A2(_2341_),
    .B1(_2342_),
    .B2(_2343_),
    .X(_2344_));
 sky130_fd_sc_hd__nor2_1 _5260_ (.A(\disp_song.um.drum.next_idx1[2] ),
    .B(_2252_),
    .Y(_2345_));
 sky130_fd_sc_hd__o22a_1 _5261_ (.A1(_2252_),
    .A2(_2323_),
    .B1(_2345_),
    .B2(_0197_),
    .X(_2346_));
 sky130_fd_sc_hd__mux2_1 _5262_ (.A0(_2340_),
    .A1(_2344_),
    .S(_2346_),
    .X(_2347_));
 sky130_fd_sc_hd__mux2_1 _5263_ (.A0(_2249_),
    .A1(_2251_),
    .S(_2256_),
    .X(_2348_));
 sky130_fd_sc_hd__mux2_1 _5264_ (.A0(\disp_song.note1[24] ),
    .A1(\disp_song.um.drum.next_note1[25] ),
    .S(_0175_),
    .X(_2349_));
 sky130_fd_sc_hd__nor2_1 _5265_ (.A(_2254_),
    .B(_2260_),
    .Y(_2350_));
 sky130_fd_sc_hd__a31o_1 _5266_ (.A1(_2254_),
    .A2(_2336_),
    .A3(_2349_),
    .B1(_2350_),
    .X(_2351_));
 sky130_fd_sc_hd__mux2_1 _5267_ (.A0(_2348_),
    .A1(_2351_),
    .S(_2339_),
    .X(_2352_));
 sky130_fd_sc_hd__mux2_1 _5268_ (.A0(_2267_),
    .A1(_2269_),
    .S(_2256_),
    .X(_2353_));
 sky130_fd_sc_hd__o211ai_1 _5269_ (.A1(_2268_),
    .A2(_2272_),
    .B1(_2271_),
    .C1(_2254_),
    .Y(_2354_));
 sky130_fd_sc_hd__o211a_1 _5270_ (.A1(_2254_),
    .A2(_2277_),
    .B1(_2339_),
    .C1(_2354_),
    .X(_2355_));
 sky130_fd_sc_hd__o21ba_1 _5271_ (.A1(_2339_),
    .A2(_2353_),
    .B1_N(_2355_),
    .X(_2356_));
 sky130_fd_sc_hd__mux2_1 _5272_ (.A0(_2352_),
    .A1(_2356_),
    .S(_2346_),
    .X(_2357_));
 sky130_fd_sc_hd__and2b_1 _5273_ (.A_N(_2333_),
    .B(_2357_),
    .X(_2358_));
 sky130_fd_sc_hd__a211o_1 _5274_ (.A1(_2333_),
    .A2(_2347_),
    .B1(_2358_),
    .C1(_2234_),
    .X(_2359_));
 sky130_fd_sc_hd__o311a_1 _5275_ (.A1(_2195_),
    .A2(_2331_),
    .A3(_2332_),
    .B1(_2359_),
    .C1(_0214_),
    .X(\disp_song.um.drum.next_d1[3] ));
 sky130_fd_sc_hd__nor2_1 _5276_ (.A(\disp_song.um.drum.next_idx1[1] ),
    .B(_2323_),
    .Y(_2360_));
 sky130_fd_sc_hd__or2_1 _5277_ (.A(_0185_),
    .B(_2360_),
    .X(_2361_));
 sky130_fd_sc_hd__nor2_1 _5278_ (.A(_2232_),
    .B(_0373_),
    .Y(_2362_));
 sky130_fd_sc_hd__a211o_1 _5279_ (.A1(\disp_song.note1[2] ),
    .A2(_2232_),
    .B1(_0191_),
    .C1(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__mux2_1 _5280_ (.A0(\disp_song.note1[18] ),
    .A1(\disp_song.um.drum.next_note1[19] ),
    .S(\disp_song.um.drum.next_idx1[0] ),
    .X(_2364_));
 sky130_fd_sc_hd__inv_2 _5281_ (.A(_2361_),
    .Y(_2365_));
 sky130_fd_sc_hd__o221a_1 _5282_ (.A1(_2185_),
    .A2(_2228_),
    .B1(_2364_),
    .B2(_0191_),
    .C1(_2365_),
    .X(_2366_));
 sky130_fd_sc_hd__a31o_1 _5283_ (.A1(_2212_),
    .A2(_2361_),
    .A3(_2363_),
    .B1(_2366_),
    .X(_2367_));
 sky130_fd_sc_hd__o21a_1 _5284_ (.A1(_0191_),
    .A2(_2203_),
    .B1(_2206_),
    .X(_2368_));
 sky130_fd_sc_hd__o21ba_1 _5285_ (.A1(_0191_),
    .A2(_2316_),
    .B1_N(_2237_),
    .X(_2369_));
 sky130_fd_sc_hd__mux2_1 _5286_ (.A0(_2368_),
    .A1(_2369_),
    .S(_2365_),
    .X(_2370_));
 sky130_fd_sc_hd__mux2_1 _5287_ (.A0(_2201_),
    .A1(_2220_),
    .S(_2365_),
    .X(_2371_));
 sky130_fd_sc_hd__o21ba_1 _5288_ (.A1(_2185_),
    .A2(_2192_),
    .B1_N(_2197_),
    .X(_2372_));
 sky130_fd_sc_hd__o21ba_1 _5289_ (.A1(_2185_),
    .A2(_2221_),
    .B1_N(_2224_),
    .X(_2373_));
 sky130_fd_sc_hd__mux2_1 _5290_ (.A0(_2372_),
    .A1(_2373_),
    .S(_2365_),
    .X(_2374_));
 sky130_fd_sc_hd__and2_1 _5291_ (.A(\disp_song.um.drum.next_idx1[3] ),
    .B(_2215_),
    .X(_2375_));
 sky130_fd_sc_hd__or2_1 _5292_ (.A(_2360_),
    .B(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__mux4_1 _5293_ (.A0(_2367_),
    .A1(_2370_),
    .A2(_2371_),
    .A3(_2374_),
    .S0(_2376_),
    .S1(_2216_),
    .X(_2377_));
 sky130_fd_sc_hd__and2_1 _5294_ (.A(_0214_),
    .B(_2377_),
    .X(_2378_));
 sky130_fd_sc_hd__clkbuf_1 _5295_ (.A(_2378_),
    .X(\disp_song.um.drum.next_d1[4] ));
 sky130_fd_sc_hd__a31o_1 _5296_ (.A1(_0191_),
    .A2(_0197_),
    .A3(_2244_),
    .B1(_0185_),
    .X(_2379_));
 sky130_fd_sc_hd__o22a_1 _5297_ (.A1(\disp_song.note1[18] ),
    .A2(_2232_),
    .B1(\disp_song.um.drum.next_idx1[1] ),
    .B2(_2226_),
    .X(_2380_));
 sky130_fd_sc_hd__o21a_1 _5298_ (.A1(\disp_song.note1[17] ),
    .A2(_2185_),
    .B1(_2271_),
    .X(_2381_));
 sky130_fd_sc_hd__o22a_1 _5299_ (.A1(_2310_),
    .A2(_2380_),
    .B1(_2381_),
    .B2(_2254_),
    .X(_2382_));
 sky130_fd_sc_hd__mux2_1 _5300_ (.A0(_2270_),
    .A1(_2382_),
    .S(_2274_),
    .X(_2383_));
 sky130_fd_sc_hd__o2bb2a_1 _5301_ (.A1_N(_2185_),
    .A2_N(_2231_),
    .B1(\disp_song.note1[26] ),
    .B2(_2232_),
    .X(_2384_));
 sky130_fd_sc_hd__o22a_1 _5302_ (.A1(_2254_),
    .A2(_2349_),
    .B1(_2384_),
    .B2(_2310_),
    .X(_2385_));
 sky130_fd_sc_hd__mux2_1 _5303_ (.A0(_2255_),
    .A1(_2385_),
    .S(_2274_),
    .X(_2386_));
 sky130_fd_sc_hd__xnor2_2 _5304_ (.A(_0197_),
    .B(_2246_),
    .Y(_2387_));
 sky130_fd_sc_hd__mux2_1 _5305_ (.A0(_2383_),
    .A1(_2386_),
    .S(_2387_),
    .X(_2388_));
 sky130_fd_sc_hd__a21o_1 _5306_ (.A1(\disp_song.um.drum.next_note1[11] ),
    .A2(_2191_),
    .B1(\disp_song.um.drum.next_idx1[1] ),
    .X(_2389_));
 sky130_fd_sc_hd__o21a_1 _5307_ (.A1(\disp_song.note1[10] ),
    .A2(_2232_),
    .B1(_2389_),
    .X(_2390_));
 sky130_fd_sc_hd__o22a_1 _5308_ (.A1(_2254_),
    .A2(_2337_),
    .B1(_2390_),
    .B2(_2310_),
    .X(_2391_));
 sky130_fd_sc_hd__or2_1 _5309_ (.A(_2247_),
    .B(_2391_),
    .X(_2392_));
 sky130_fd_sc_hd__o211a_1 _5310_ (.A1(_2274_),
    .A2(_2286_),
    .B1(_2387_),
    .C1(_2392_),
    .X(_2393_));
 sky130_fd_sc_hd__o22a_1 _5311_ (.A1(\disp_song.note1[2] ),
    .A2(_2232_),
    .B1(\disp_song.um.drum.next_idx1[1] ),
    .B2(_2209_),
    .X(_2394_));
 sky130_fd_sc_hd__o22a_1 _5312_ (.A1(\disp_song.note1[1] ),
    .A2(_2185_),
    .B1(\disp_song.um.drum.next_note1[0] ),
    .B2(_2232_),
    .X(_2395_));
 sky130_fd_sc_hd__o22a_1 _5313_ (.A1(_2310_),
    .A2(_2394_),
    .B1(_2395_),
    .B2(_2254_),
    .X(_2396_));
 sky130_fd_sc_hd__mux2_1 _5314_ (.A0(_2297_),
    .A1(_2396_),
    .S(_2274_),
    .X(_2397_));
 sky130_fd_sc_hd__inv_2 _5315_ (.A(_2397_),
    .Y(_2398_));
 sky130_fd_sc_hd__o21ai_1 _5316_ (.A1(_2387_),
    .A2(_2398_),
    .B1(_2379_),
    .Y(_2399_));
 sky130_fd_sc_hd__o221a_1 _5317_ (.A1(_2379_),
    .A2(_2388_),
    .B1(_2393_),
    .B2(_2399_),
    .C1(_0214_),
    .X(\disp_song.um.drum.next_d1[5] ));
 sky130_fd_sc_hd__a32o_1 _5318_ (.A1(\disp_song.um.drum.next_note1[3] ),
    .A2(_2208_),
    .A3(_2252_),
    .B1(_2314_),
    .B2(\disp_song.um.drum.next_note1[4] ),
    .X(_2400_));
 sky130_fd_sc_hd__a41o_1 _5319_ (.A1(_0179_),
    .A2(_2232_),
    .A3(\disp_song.um.drum.next_note1[2] ),
    .A4(_2208_),
    .B1(_2400_),
    .X(_2401_));
 sky130_fd_sc_hd__a221o_1 _5320_ (.A1(\disp_song.um.drum.next_note1[5] ),
    .A2(_2312_),
    .B1(_2360_),
    .B2(_2211_),
    .C1(_2195_),
    .X(_2402_));
 sky130_fd_sc_hd__mux2_1 _5321_ (.A0(_2228_),
    .A1(_2364_),
    .S(\disp_song.um.drum.next_idx1[1] ),
    .X(_2403_));
 sky130_fd_sc_hd__mux2_1 _5322_ (.A0(_2318_),
    .A1(_2403_),
    .S(_0191_),
    .X(_2404_));
 sky130_fd_sc_hd__mux2_1 _5323_ (.A0(_2221_),
    .A1(_2223_),
    .S(\disp_song.um.drum.next_idx1[1] ),
    .X(_2405_));
 sky130_fd_sc_hd__mux2_1 _5324_ (.A0(_2317_),
    .A1(_2405_),
    .S(\disp_song.um.drum.next_idx1[2] ),
    .X(_2406_));
 sky130_fd_sc_hd__or2_1 _5325_ (.A(_2187_),
    .B(_2199_),
    .X(_2407_));
 sky130_fd_sc_hd__mux2_1 _5326_ (.A0(_2325_),
    .A1(_2326_),
    .S(\disp_song.um.drum.next_idx1[2] ),
    .X(_2408_));
 sky130_fd_sc_hd__mux4_1 _5327_ (.A0(_2404_),
    .A1(_2406_),
    .A2(_2407_),
    .A3(_2408_),
    .S0(\disp_song.um.drum.next_idx1[3] ),
    .S1(_0185_),
    .X(_2409_));
 sky130_fd_sc_hd__o211a_1 _5328_ (.A1(_2401_),
    .A2(_2402_),
    .B1(_2409_),
    .C1(_0214_),
    .X(\disp_song.um.drum.next_d1[6] ));
 sky130_fd_sc_hd__inv_2 _5329_ (.A(_0366_),
    .Y(\disp_song.next_green ));
 sky130_fd_sc_hd__nand3_1 _5330_ (.A(_0209_),
    .B(_2658_),
    .C(_1302_),
    .Y(_2410_));
 sky130_fd_sc_hd__inv_2 _5331_ (.A(_2410_),
    .Y(_2411_));
 sky130_fd_sc_hd__or2_1 _5332_ (.A(net252),
    .B(_2411_),
    .X(_2412_));
 sky130_fd_sc_hd__clkbuf_1 _5333_ (.A(_2412_),
    .X(_0033_));
 sky130_fd_sc_hd__and2_1 _5334_ (.A(\game.scoring_button_2.acc[2] ),
    .B(_2410_),
    .X(_2413_));
 sky130_fd_sc_hd__clkbuf_1 _5335_ (.A(_2413_),
    .X(_0034_));
 sky130_fd_sc_hd__nand2_1 _5336_ (.A(_1021_),
    .B(_1022_),
    .Y(_2414_));
 sky130_fd_sc_hd__o31a_1 _5337_ (.A1(_1028_),
    .A2(_1029_),
    .A3(_1030_),
    .B1(\highest_score.highest_score[1] ),
    .X(_2415_));
 sky130_fd_sc_hd__o21ai_1 _5338_ (.A1(_1012_),
    .A2(_1028_),
    .B1(_1057_),
    .Y(_2416_));
 sky130_fd_sc_hd__or4_1 _5339_ (.A(\highest_score.highest_score[1] ),
    .B(_1028_),
    .C(_1029_),
    .D(_1030_),
    .X(_2417_));
 sky130_fd_sc_hd__o221a_1 _5340_ (.A1(\highest_score.highest_score[2] ),
    .A2(_2414_),
    .B1(_2415_),
    .B2(_2416_),
    .C1(_2417_),
    .X(_2418_));
 sky130_fd_sc_hd__a22o_1 _5341_ (.A1(\highest_score.highest_score[2] ),
    .A2(_2414_),
    .B1(_1024_),
    .B2(\highest_score.highest_score[3] ),
    .X(_2419_));
 sky130_fd_sc_hd__o22a_1 _5342_ (.A1(\highest_score.highest_score[4] ),
    .A2(_0855_),
    .B1(_1024_),
    .B2(\highest_score.highest_score[3] ),
    .X(_2420_));
 sky130_fd_sc_hd__a22o_1 _5343_ (.A1(\highest_score.highest_score[5] ),
    .A2(_0840_),
    .B1(_0855_),
    .B2(\highest_score.highest_score[4] ),
    .X(_2421_));
 sky130_fd_sc_hd__inv_2 _5344_ (.A(_2421_),
    .Y(_2422_));
 sky130_fd_sc_hd__and3_1 _5345_ (.A(\highest_score.highest_score[7] ),
    .B(_0841_),
    .C(_0847_),
    .X(_2423_));
 sky130_fd_sc_hd__a21o_1 _5346_ (.A1(_0841_),
    .A2(_0847_),
    .B1(\highest_score.highest_score[7] ),
    .X(_2424_));
 sky130_fd_sc_hd__xnor2_1 _5347_ (.A(\highest_score.highest_score[6] ),
    .B(_0858_),
    .Y(_2425_));
 sky130_fd_sc_hd__or2_1 _5348_ (.A(\highest_score.highest_score[5] ),
    .B(_0840_),
    .X(_2426_));
 sky130_fd_sc_hd__and4b_1 _5349_ (.A_N(_2423_),
    .B(_2424_),
    .C(_2425_),
    .D(_2426_),
    .X(_2427_));
 sky130_fd_sc_hd__o2111a_1 _5350_ (.A1(_2418_),
    .A2(_2419_),
    .B1(_2420_),
    .C1(_2422_),
    .D1(_2427_),
    .X(_2428_));
 sky130_fd_sc_hd__and3b_1 _5351_ (.A_N(_2423_),
    .B(_2424_),
    .C(_2425_),
    .X(_2429_));
 sky130_fd_sc_hd__and2_1 _5352_ (.A(_2426_),
    .B(_2421_),
    .X(_2430_));
 sky130_fd_sc_hd__and4b_1 _5353_ (.A_N(_2423_),
    .B(\highest_score.highest_score[6] ),
    .C(_0835_),
    .D(_2424_),
    .X(_2431_));
 sky130_fd_sc_hd__a2111oi_1 _5354_ (.A1(_2429_),
    .A2(_2430_),
    .B1(_2431_),
    .C1(_0921_),
    .D1(_2423_),
    .Y(_2432_));
 sky130_fd_sc_hd__or3b_1 _5355_ (.A(net42),
    .B(_2428_),
    .C_N(_2432_),
    .X(_2433_));
 sky130_fd_sc_hd__buf_2 _5356_ (.A(_2433_),
    .X(_2434_));
 sky130_fd_sc_hd__mux2_1 _5357_ (.A0(_1034_),
    .A1(\highest_score.highest_score[0] ),
    .S(_2434_),
    .X(_2435_));
 sky130_fd_sc_hd__clkbuf_1 _5358_ (.A(_2435_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _5359_ (.A0(_1035_),
    .A1(\highest_score.highest_score[1] ),
    .S(_2434_),
    .X(_2436_));
 sky130_fd_sc_hd__clkbuf_1 _5360_ (.A(_2436_),
    .X(_0036_));
 sky130_fd_sc_hd__and2_1 _5361_ (.A(_1021_),
    .B(_1022_),
    .X(_2437_));
 sky130_fd_sc_hd__mux2_1 _5362_ (.A0(_2437_),
    .A1(\highest_score.highest_score[2] ),
    .S(_2434_),
    .X(_2438_));
 sky130_fd_sc_hd__clkbuf_1 _5363_ (.A(_2438_),
    .X(_0037_));
 sky130_fd_sc_hd__inv_2 _5364_ (.A(_1024_),
    .Y(_2439_));
 sky130_fd_sc_hd__mux2_1 _5365_ (.A0(_2439_),
    .A1(\highest_score.highest_score[3] ),
    .S(_2434_),
    .X(_2440_));
 sky130_fd_sc_hd__clkbuf_1 _5366_ (.A(_2440_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _5367_ (.A0(_0946_),
    .A1(\highest_score.highest_score[4] ),
    .S(_2434_),
    .X(_2441_));
 sky130_fd_sc_hd__clkbuf_1 _5368_ (.A(_2441_),
    .X(_0039_));
 sky130_fd_sc_hd__nor2_1 _5369_ (.A(_0830_),
    .B(_0838_),
    .Y(_2442_));
 sky130_fd_sc_hd__a211o_1 _5370_ (.A1(_0830_),
    .A2(_0791_),
    .B1(_0857_),
    .C1(_2442_),
    .X(_2443_));
 sky130_fd_sc_hd__inv_2 _5371_ (.A(_2443_),
    .Y(_2444_));
 sky130_fd_sc_hd__mux2_1 _5372_ (.A0(_2444_),
    .A1(\highest_score.highest_score[5] ),
    .S(_2434_),
    .X(_2445_));
 sky130_fd_sc_hd__clkbuf_1 _5373_ (.A(_2445_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _5374_ (.A0(_0858_),
    .A1(\highest_score.highest_score[6] ),
    .S(_2434_),
    .X(_2446_));
 sky130_fd_sc_hd__clkbuf_1 _5375_ (.A(_2446_),
    .X(_0041_));
 sky130_fd_sc_hd__o21ai_1 _5376_ (.A1(_0848_),
    .A2(_2434_),
    .B1(_0899_),
    .Y(_0042_));
 sky130_fd_sc_hd__or2b_1 _5377_ (.A(\game.beat_clk ),
    .B_N(_0206_),
    .X(_2447_));
 sky130_fd_sc_hd__nand2_1 _5378_ (.A(net179),
    .B(_2447_),
    .Y(_2448_));
 sky130_fd_sc_hd__o21a_1 _5379_ (.A1(net179),
    .A2(net123),
    .B1(_2448_),
    .X(_0043_));
 sky130_fd_sc_hd__nand3_1 _5380_ (.A(\pulseout.fin_pulse[0] ),
    .B(\pulseout.fin_pulse[1] ),
    .C(\game.beat_clk ),
    .Y(_2449_));
 sky130_fd_sc_hd__a21o_1 _5381_ (.A1(\pulseout.fin_pulse[0] ),
    .A2(\game.beat_clk ),
    .B1(\pulseout.fin_pulse[1] ),
    .X(_2450_));
 sky130_fd_sc_hd__and3_1 _5382_ (.A(_0206_),
    .B(_2449_),
    .C(_2450_),
    .X(_2451_));
 sky130_fd_sc_hd__clkbuf_1 _5383_ (.A(_2451_),
    .X(_0044_));
 sky130_fd_sc_hd__xnor2_1 _5384_ (.A(net128),
    .B(_2449_),
    .Y(_0045_));
 sky130_fd_sc_hd__a41o_1 _5385_ (.A1(\pulseout.fin_pulse[0] ),
    .A2(\pulseout.fin_pulse[1] ),
    .A3(\pulseout.fin_pulse[2] ),
    .A4(\game.beat_clk ),
    .B1(\pulseout.fin_pulse[3] ),
    .X(_2452_));
 sky130_fd_sc_hd__and4_1 _5386_ (.A(\pulseout.fin_pulse[0] ),
    .B(\pulseout.fin_pulse[1] ),
    .C(\pulseout.fin_pulse[2] ),
    .D(\pulseout.fin_pulse[3] ),
    .X(_2453_));
 sky130_fd_sc_hd__nand2_1 _5387_ (.A(_2447_),
    .B(_2453_),
    .Y(_2454_));
 sky130_fd_sc_hd__and3_1 _5388_ (.A(_0206_),
    .B(_2452_),
    .C(_2454_),
    .X(_2455_));
 sky130_fd_sc_hd__clkbuf_1 _5389_ (.A(_2455_),
    .X(_0046_));
 sky130_fd_sc_hd__xnor2_1 _5390_ (.A(net147),
    .B(_2454_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _5391_ (.A(\pulseout.fin_pulse[4] ),
    .Y(_2456_));
 sky130_fd_sc_hd__a31o_1 _5392_ (.A1(\pulseout.fin_pulse[4] ),
    .A2(\game.beat_clk ),
    .A3(_2453_),
    .B1(net265),
    .X(_2457_));
 sky130_fd_sc_hd__o311a_1 _5393_ (.A1(_2456_),
    .A2(_0204_),
    .A3(_2454_),
    .B1(_2457_),
    .C1(_0206_),
    .X(_0048_));
 sky130_fd_sc_hd__o22a_1 _5394_ (.A1(\game.scoring_button_2.check_hit.edge_1 ),
    .A2(_1287_),
    .B1(net131),
    .B2(_2411_),
    .X(_0049_));
 sky130_fd_sc_hd__and2b_1 _5395_ (.A_N(_0209_),
    .B(\modetrans.mode[5] ),
    .X(_2458_));
 sky130_fd_sc_hd__and2_1 _5396_ (.A(\game.beat_clk ),
    .B(_0209_),
    .X(_2459_));
 sky130_fd_sc_hd__buf_4 _5397_ (.A(_2459_),
    .X(_2460_));
 sky130_fd_sc_hd__nor2_1 _5398_ (.A(_2458_),
    .B(_2460_),
    .Y(_2461_));
 sky130_fd_sc_hd__buf_6 _5399_ (.A(_2461_),
    .X(_2462_));
 sky130_fd_sc_hd__a22o_1 _5400_ (.A1(\disp_song.note2[0] ),
    .A2(_2458_),
    .B1(_2462_),
    .B2(net91),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _5401_ (.A0(\disp_song.note2[1] ),
    .A1(\game.padded_notes2[0] ),
    .S(_0219_),
    .X(_2463_));
 sky130_fd_sc_hd__mux2_1 _5402_ (.A0(_2463_),
    .A1(\game.padded_notes2[1] ),
    .S(_2462_),
    .X(_2464_));
 sky130_fd_sc_hd__clkbuf_1 _5403_ (.A(_2464_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _5404_ (.A0(\disp_song.note2[2] ),
    .A1(\game.padded_notes2[1] ),
    .S(_0219_),
    .X(_2465_));
 sky130_fd_sc_hd__mux2_1 _5405_ (.A0(_2465_),
    .A1(net242),
    .S(_2462_),
    .X(_2466_));
 sky130_fd_sc_hd__clkbuf_1 _5406_ (.A(_2466_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _5407_ (.A0(\disp_song.note2[3] ),
    .A1(\game.padded_notes2[2] ),
    .S(_0219_),
    .X(_2467_));
 sky130_fd_sc_hd__mux2_1 _5408_ (.A0(_2467_),
    .A1(\game.padded_notes2[3] ),
    .S(_2462_),
    .X(_2468_));
 sky130_fd_sc_hd__clkbuf_1 _5409_ (.A(_2468_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _5410_ (.A0(\disp_song.note2[4] ),
    .A1(\game.padded_notes2[3] ),
    .S(_0219_),
    .X(_2469_));
 sky130_fd_sc_hd__mux2_1 _5411_ (.A0(_2469_),
    .A1(net254),
    .S(_2462_),
    .X(_2470_));
 sky130_fd_sc_hd__clkbuf_1 _5412_ (.A(_2470_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _5413_ (.A0(\disp_song.note2[5] ),
    .A1(\game.padded_notes2[4] ),
    .S(_0219_),
    .X(_2471_));
 sky130_fd_sc_hd__buf_8 _5414_ (.A(_2461_),
    .X(_2472_));
 sky130_fd_sc_hd__buf_8 _5415_ (.A(_2472_),
    .X(_2473_));
 sky130_fd_sc_hd__mux2_1 _5416_ (.A0(_2471_),
    .A1(\game.padded_notes2[5] ),
    .S(_2473_),
    .X(_2474_));
 sky130_fd_sc_hd__clkbuf_1 _5417_ (.A(_2474_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _5418_ (.A0(\disp_song.note2[6] ),
    .A1(\game.padded_notes2[5] ),
    .S(_0219_),
    .X(_2475_));
 sky130_fd_sc_hd__mux2_1 _5419_ (.A0(_2475_),
    .A1(net227),
    .S(_2473_),
    .X(_2476_));
 sky130_fd_sc_hd__clkbuf_1 _5420_ (.A(_2476_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _5421_ (.A0(\disp_song.note2[7] ),
    .A1(\game.padded_notes2[6] ),
    .S(_0219_),
    .X(_2477_));
 sky130_fd_sc_hd__mux2_1 _5422_ (.A0(_2477_),
    .A1(\game.padded_notes2[7] ),
    .S(_2473_),
    .X(_2478_));
 sky130_fd_sc_hd__clkbuf_1 _5423_ (.A(_2478_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _5424_ (.A0(\disp_song.note2[8] ),
    .A1(\game.padded_notes2[7] ),
    .S(_0219_),
    .X(_2479_));
 sky130_fd_sc_hd__mux2_1 _5425_ (.A0(_2479_),
    .A1(net209),
    .S(_2473_),
    .X(_2480_));
 sky130_fd_sc_hd__clkbuf_1 _5426_ (.A(_2480_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _5427_ (.A0(\disp_song.note2[9] ),
    .A1(\game.padded_notes2[8] ),
    .S(_0219_),
    .X(_2481_));
 sky130_fd_sc_hd__mux2_1 _5428_ (.A0(_2481_),
    .A1(\game.padded_notes2[9] ),
    .S(_2473_),
    .X(_2482_));
 sky130_fd_sc_hd__clkbuf_1 _5429_ (.A(_2482_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _5430_ (.A0(\disp_song.note2[10] ),
    .A1(\game.padded_notes2[9] ),
    .S(_0219_),
    .X(_2483_));
 sky130_fd_sc_hd__mux2_1 _5431_ (.A0(_2483_),
    .A1(net229),
    .S(_2473_),
    .X(_2484_));
 sky130_fd_sc_hd__clkbuf_1 _5432_ (.A(_2484_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _5433_ (.A0(\disp_song.note2[11] ),
    .A1(\game.padded_notes2[10] ),
    .S(_0219_),
    .X(_2485_));
 sky130_fd_sc_hd__mux2_1 _5434_ (.A0(_2485_),
    .A1(\game.padded_notes2[11] ),
    .S(_2473_),
    .X(_2486_));
 sky130_fd_sc_hd__clkbuf_1 _5435_ (.A(_2486_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _5436_ (.A0(\disp_song.note2[12] ),
    .A1(\game.padded_notes2[11] ),
    .S(_0219_),
    .X(_2487_));
 sky130_fd_sc_hd__mux2_1 _5437_ (.A0(_2487_),
    .A1(net235),
    .S(_2473_),
    .X(_2488_));
 sky130_fd_sc_hd__clkbuf_1 _5438_ (.A(_2488_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _5439_ (.A0(\disp_song.note2[13] ),
    .A1(\game.padded_notes2[12] ),
    .S(_0219_),
    .X(_2489_));
 sky130_fd_sc_hd__mux2_1 _5440_ (.A0(_2489_),
    .A1(\game.padded_notes2[13] ),
    .S(_2473_),
    .X(_2490_));
 sky130_fd_sc_hd__clkbuf_1 _5441_ (.A(_2490_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _5442_ (.A0(\disp_song.note2[14] ),
    .A1(\game.padded_notes2[13] ),
    .S(_0219_),
    .X(_2491_));
 sky130_fd_sc_hd__mux2_1 _5443_ (.A0(_2491_),
    .A1(net231),
    .S(_2473_),
    .X(_2492_));
 sky130_fd_sc_hd__clkbuf_1 _5444_ (.A(_2492_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _5445_ (.A0(\disp_song.note2[15] ),
    .A1(\game.padded_notes2[14] ),
    .S(_0219_),
    .X(_2493_));
 sky130_fd_sc_hd__mux2_1 _5446_ (.A0(_2493_),
    .A1(\game.padded_notes2[15] ),
    .S(_2473_),
    .X(_2494_));
 sky130_fd_sc_hd__clkbuf_1 _5447_ (.A(_2494_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _5448_ (.A0(\disp_song.note2[16] ),
    .A1(\game.padded_notes2[15] ),
    .S(_0219_),
    .X(_2495_));
 sky130_fd_sc_hd__mux2_1 _5449_ (.A0(_2495_),
    .A1(net261),
    .S(_2473_),
    .X(_2496_));
 sky130_fd_sc_hd__clkbuf_1 _5450_ (.A(_2496_),
    .X(_0066_));
 sky130_fd_sc_hd__buf_8 _5451_ (.A(_0209_),
    .X(_2497_));
 sky130_fd_sc_hd__mux2_1 _5452_ (.A0(\disp_song.note2[17] ),
    .A1(\game.padded_notes2[16] ),
    .S(_2497_),
    .X(_2498_));
 sky130_fd_sc_hd__mux2_1 _5453_ (.A0(_2498_),
    .A1(\game.padded_notes2[17] ),
    .S(_2473_),
    .X(_2499_));
 sky130_fd_sc_hd__clkbuf_1 _5454_ (.A(_2499_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _5455_ (.A0(\disp_song.note2[18] ),
    .A1(\game.padded_notes2[17] ),
    .S(_2497_),
    .X(_2500_));
 sky130_fd_sc_hd__mux2_1 _5456_ (.A0(_2500_),
    .A1(net230),
    .S(_2473_),
    .X(_2501_));
 sky130_fd_sc_hd__clkbuf_1 _5457_ (.A(_2501_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _5458_ (.A0(\disp_song.note2[19] ),
    .A1(\game.padded_notes2[18] ),
    .S(_2497_),
    .X(_2502_));
 sky130_fd_sc_hd__mux2_1 _5459_ (.A0(_2502_),
    .A1(\game.padded_notes2[19] ),
    .S(_2473_),
    .X(_2503_));
 sky130_fd_sc_hd__clkbuf_1 _5460_ (.A(_2503_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _5461_ (.A0(\disp_song.note2[20] ),
    .A1(\game.padded_notes2[19] ),
    .S(_2497_),
    .X(_2504_));
 sky130_fd_sc_hd__mux2_1 _5462_ (.A0(_2504_),
    .A1(net251),
    .S(_2473_),
    .X(_2505_));
 sky130_fd_sc_hd__clkbuf_1 _5463_ (.A(_2505_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _5464_ (.A0(\disp_song.note2[21] ),
    .A1(\game.padded_notes2[20] ),
    .S(_2497_),
    .X(_2506_));
 sky130_fd_sc_hd__mux2_1 _5465_ (.A0(_2506_),
    .A1(\game.padded_notes2[21] ),
    .S(_2473_),
    .X(_2507_));
 sky130_fd_sc_hd__clkbuf_1 _5466_ (.A(_2507_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _5467_ (.A0(\disp_song.note2[22] ),
    .A1(\game.padded_notes2[21] ),
    .S(_2497_),
    .X(_2508_));
 sky130_fd_sc_hd__mux2_1 _5468_ (.A0(_2508_),
    .A1(net211),
    .S(_2473_),
    .X(_2509_));
 sky130_fd_sc_hd__clkbuf_1 _5469_ (.A(_2509_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _5470_ (.A0(\disp_song.note2[23] ),
    .A1(\game.padded_notes2[22] ),
    .S(_2497_),
    .X(_2510_));
 sky130_fd_sc_hd__mux2_1 _5471_ (.A0(_2510_),
    .A1(\game.padded_notes2[23] ),
    .S(_2473_),
    .X(_2511_));
 sky130_fd_sc_hd__clkbuf_1 _5472_ (.A(_2511_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _5473_ (.A0(\disp_song.note2[24] ),
    .A1(\game.padded_notes2[23] ),
    .S(_2497_),
    .X(_2512_));
 sky130_fd_sc_hd__mux2_1 _5474_ (.A0(_2512_),
    .A1(net221),
    .S(_2473_),
    .X(_2513_));
 sky130_fd_sc_hd__clkbuf_1 _5475_ (.A(_2513_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _5476_ (.A0(\disp_song.note2[25] ),
    .A1(\game.padded_notes2[24] ),
    .S(_2497_),
    .X(_2514_));
 sky130_fd_sc_hd__buf_8 _5477_ (.A(_2472_),
    .X(_2515_));
 sky130_fd_sc_hd__mux2_1 _5478_ (.A0(_2514_),
    .A1(\game.padded_notes2[25] ),
    .S(_2515_),
    .X(_2516_));
 sky130_fd_sc_hd__clkbuf_1 _5479_ (.A(_2516_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _5480_ (.A0(\disp_song.note2[26] ),
    .A1(\game.padded_notes2[25] ),
    .S(_2497_),
    .X(_2517_));
 sky130_fd_sc_hd__mux2_1 _5481_ (.A0(_2517_),
    .A1(net239),
    .S(_2515_),
    .X(_2518_));
 sky130_fd_sc_hd__clkbuf_1 _5482_ (.A(_2518_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _5483_ (.A0(\disp_song.note2[27] ),
    .A1(\game.padded_notes2[26] ),
    .S(_2497_),
    .X(_2519_));
 sky130_fd_sc_hd__mux2_1 _5484_ (.A0(_2519_),
    .A1(\game.padded_notes2[27] ),
    .S(_2515_),
    .X(_2520_));
 sky130_fd_sc_hd__clkbuf_1 _5485_ (.A(_2520_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _5486_ (.A0(\disp_song.note2[28] ),
    .A1(\game.padded_notes2[27] ),
    .S(_2497_),
    .X(_2521_));
 sky130_fd_sc_hd__mux2_1 _5487_ (.A0(_2521_),
    .A1(net233),
    .S(_2515_),
    .X(_2522_));
 sky130_fd_sc_hd__clkbuf_1 _5488_ (.A(_2522_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _5489_ (.A0(\disp_song.note2[29] ),
    .A1(\game.padded_notes2[28] ),
    .S(_2497_),
    .X(_2523_));
 sky130_fd_sc_hd__mux2_1 _5490_ (.A0(_2523_),
    .A1(\game.padded_notes2[29] ),
    .S(_2515_),
    .X(_2524_));
 sky130_fd_sc_hd__clkbuf_1 _5491_ (.A(_2524_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _5492_ (.A0(\disp_song.note2[30] ),
    .A1(\game.padded_notes2[29] ),
    .S(_2497_),
    .X(_2525_));
 sky130_fd_sc_hd__mux2_1 _5493_ (.A0(_2525_),
    .A1(net234),
    .S(_2515_),
    .X(_2526_));
 sky130_fd_sc_hd__clkbuf_1 _5494_ (.A(_2526_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _5495_ (.A0(\disp_song.note2[31] ),
    .A1(\game.padded_notes2[30] ),
    .S(_2497_),
    .X(_2527_));
 sky130_fd_sc_hd__mux2_1 _5496_ (.A0(_2527_),
    .A1(\game.padded_notes2[31] ),
    .S(_2515_),
    .X(_2528_));
 sky130_fd_sc_hd__clkbuf_1 _5497_ (.A(_2528_),
    .X(_0081_));
 sky130_fd_sc_hd__a22o_1 _5498_ (.A1(\game.padded_notes2[31] ),
    .A2(_2460_),
    .B1(_2462_),
    .B2(net133),
    .X(_0082_));
 sky130_fd_sc_hd__a22o_1 _5499_ (.A1(net133),
    .A2(_2460_),
    .B1(_2462_),
    .B2(net143),
    .X(_0083_));
 sky130_fd_sc_hd__a22o_1 _5500_ (.A1(\game.out[8] ),
    .A2(_2460_),
    .B1(_2462_),
    .B2(net140),
    .X(_0084_));
 sky130_fd_sc_hd__a22o_1 _5501_ (.A1(net140),
    .A2(_2460_),
    .B1(_2462_),
    .B2(net145),
    .X(_0085_));
 sky130_fd_sc_hd__a22o_1 _5502_ (.A1(\game.out[10] ),
    .A2(_2460_),
    .B1(_2462_),
    .B2(net117),
    .X(_0086_));
 sky130_fd_sc_hd__a22o_1 _5503_ (.A1(net117),
    .A2(_2460_),
    .B1(_2462_),
    .B2(\game.out[12] ),
    .X(_0087_));
 sky130_fd_sc_hd__a22o_1 _5504_ (.A1(net269),
    .A2(_2460_),
    .B1(_2462_),
    .B2(net110),
    .X(_0088_));
 sky130_fd_sc_hd__nand3_1 _5505_ (.A(_0209_),
    .B(_2656_),
    .C(_1688_),
    .Y(_2529_));
 sky130_fd_sc_hd__inv_2 _5506_ (.A(_2529_),
    .Y(_2530_));
 sky130_fd_sc_hd__o21a_1 _5507_ (.A1(net170),
    .A2(_2530_),
    .B1(_1673_),
    .X(_0089_));
 sky130_fd_sc_hd__a22o_1 _5508_ (.A1(net97),
    .A2(_2458_),
    .B1(_2462_),
    .B2(\game.padded_notes1[0] ),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _5509_ (.A0(\disp_song.note1[1] ),
    .A1(\game.padded_notes1[0] ),
    .S(_2497_),
    .X(_2531_));
 sky130_fd_sc_hd__mux2_1 _5510_ (.A0(_2531_),
    .A1(net232),
    .S(_2515_),
    .X(_2532_));
 sky130_fd_sc_hd__clkbuf_1 _5511_ (.A(_2532_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _5512_ (.A0(\disp_song.note1[2] ),
    .A1(\game.padded_notes1[1] ),
    .S(_2497_),
    .X(_2533_));
 sky130_fd_sc_hd__mux2_1 _5513_ (.A0(_2533_),
    .A1(\game.padded_notes1[2] ),
    .S(_2515_),
    .X(_2534_));
 sky130_fd_sc_hd__clkbuf_1 _5514_ (.A(_2534_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _5515_ (.A0(\disp_song.note1[3] ),
    .A1(\game.padded_notes1[2] ),
    .S(_2497_),
    .X(_2535_));
 sky130_fd_sc_hd__mux2_1 _5516_ (.A0(_2535_),
    .A1(\game.padded_notes1[3] ),
    .S(_2515_),
    .X(_2536_));
 sky130_fd_sc_hd__clkbuf_1 _5517_ (.A(_2536_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _5518_ (.A0(\disp_song.note1[4] ),
    .A1(\game.padded_notes1[3] ),
    .S(_2497_),
    .X(_2537_));
 sky130_fd_sc_hd__mux2_1 _5519_ (.A0(_2537_),
    .A1(net218),
    .S(_2515_),
    .X(_2538_));
 sky130_fd_sc_hd__clkbuf_1 _5520_ (.A(_2538_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _5521_ (.A0(\disp_song.note1[5] ),
    .A1(\game.padded_notes1[4] ),
    .S(_2497_),
    .X(_2539_));
 sky130_fd_sc_hd__mux2_1 _5522_ (.A0(_2539_),
    .A1(net256),
    .S(_2515_),
    .X(_2540_));
 sky130_fd_sc_hd__clkbuf_1 _5523_ (.A(_2540_),
    .X(_0095_));
 sky130_fd_sc_hd__buf_6 _5524_ (.A(_0209_),
    .X(_2541_));
 sky130_fd_sc_hd__mux2_1 _5525_ (.A0(\disp_song.note1[6] ),
    .A1(\game.padded_notes1[5] ),
    .S(_2541_),
    .X(_2542_));
 sky130_fd_sc_hd__mux2_1 _5526_ (.A0(_2542_),
    .A1(\game.padded_notes1[6] ),
    .S(_2515_),
    .X(_2543_));
 sky130_fd_sc_hd__clkbuf_1 _5527_ (.A(_2543_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _5528_ (.A0(\disp_song.note1[7] ),
    .A1(\game.padded_notes1[6] ),
    .S(_2541_),
    .X(_2544_));
 sky130_fd_sc_hd__mux2_1 _5529_ (.A0(_2544_),
    .A1(\game.padded_notes1[7] ),
    .S(_2515_),
    .X(_2545_));
 sky130_fd_sc_hd__clkbuf_1 _5530_ (.A(_2545_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _5531_ (.A0(\disp_song.note1[8] ),
    .A1(\game.padded_notes1[7] ),
    .S(_2541_),
    .X(_2546_));
 sky130_fd_sc_hd__mux2_1 _5532_ (.A0(_2546_),
    .A1(net224),
    .S(_2515_),
    .X(_2547_));
 sky130_fd_sc_hd__clkbuf_1 _5533_ (.A(_2547_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _5534_ (.A0(\disp_song.note1[9] ),
    .A1(\game.padded_notes1[8] ),
    .S(_2541_),
    .X(_2548_));
 sky130_fd_sc_hd__mux2_1 _5535_ (.A0(_2548_),
    .A1(net214),
    .S(_2515_),
    .X(_2549_));
 sky130_fd_sc_hd__clkbuf_1 _5536_ (.A(_2549_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _5537_ (.A0(\disp_song.note1[10] ),
    .A1(\game.padded_notes1[9] ),
    .S(_2541_),
    .X(_2550_));
 sky130_fd_sc_hd__mux2_1 _5538_ (.A0(_2550_),
    .A1(\game.padded_notes1[10] ),
    .S(_2515_),
    .X(_2551_));
 sky130_fd_sc_hd__clkbuf_1 _5539_ (.A(_2551_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _5540_ (.A0(\disp_song.note1[11] ),
    .A1(\game.padded_notes1[10] ),
    .S(_2541_),
    .X(_2552_));
 sky130_fd_sc_hd__mux2_1 _5541_ (.A0(_2552_),
    .A1(\game.padded_notes1[11] ),
    .S(_2515_),
    .X(_2553_));
 sky130_fd_sc_hd__clkbuf_1 _5542_ (.A(_2553_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _5543_ (.A0(\disp_song.note1[12] ),
    .A1(\game.padded_notes1[11] ),
    .S(_2541_),
    .X(_2554_));
 sky130_fd_sc_hd__mux2_1 _5544_ (.A0(_2554_),
    .A1(net241),
    .S(_2515_),
    .X(_2555_));
 sky130_fd_sc_hd__clkbuf_1 _5545_ (.A(_2555_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _5546_ (.A0(\disp_song.note1[13] ),
    .A1(\game.padded_notes1[12] ),
    .S(_2541_),
    .X(_2556_));
 sky130_fd_sc_hd__mux2_1 _5547_ (.A0(_2556_),
    .A1(net243),
    .S(_2515_),
    .X(_2557_));
 sky130_fd_sc_hd__clkbuf_1 _5548_ (.A(_2557_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _5549_ (.A0(\disp_song.note1[14] ),
    .A1(\game.padded_notes1[13] ),
    .S(_2541_),
    .X(_2558_));
 sky130_fd_sc_hd__mux2_1 _5550_ (.A0(_2558_),
    .A1(\game.padded_notes1[14] ),
    .S(_2472_),
    .X(_2559_));
 sky130_fd_sc_hd__clkbuf_1 _5551_ (.A(_2559_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _5552_ (.A0(\disp_song.note1[15] ),
    .A1(\game.padded_notes1[14] ),
    .S(_2541_),
    .X(_2560_));
 sky130_fd_sc_hd__mux2_1 _5553_ (.A0(_2560_),
    .A1(\game.padded_notes1[15] ),
    .S(_2472_),
    .X(_2561_));
 sky130_fd_sc_hd__clkbuf_1 _5554_ (.A(_2561_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _5555_ (.A0(\disp_song.note1[16] ),
    .A1(\game.padded_notes1[15] ),
    .S(_2541_),
    .X(_2562_));
 sky130_fd_sc_hd__mux2_1 _5556_ (.A0(_2562_),
    .A1(net226),
    .S(_2472_),
    .X(_2563_));
 sky130_fd_sc_hd__clkbuf_1 _5557_ (.A(_2563_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _5558_ (.A0(\disp_song.note1[17] ),
    .A1(\game.padded_notes1[16] ),
    .S(_2541_),
    .X(_2564_));
 sky130_fd_sc_hd__mux2_1 _5559_ (.A0(_2564_),
    .A1(net238),
    .S(_2472_),
    .X(_2565_));
 sky130_fd_sc_hd__clkbuf_1 _5560_ (.A(_2565_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _5561_ (.A0(\disp_song.note1[18] ),
    .A1(\game.padded_notes1[17] ),
    .S(_2541_),
    .X(_2566_));
 sky130_fd_sc_hd__mux2_1 _5562_ (.A0(_2566_),
    .A1(\game.padded_notes1[18] ),
    .S(_2472_),
    .X(_2567_));
 sky130_fd_sc_hd__clkbuf_1 _5563_ (.A(_2567_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _5564_ (.A0(\disp_song.note1[19] ),
    .A1(\game.padded_notes1[18] ),
    .S(_2541_),
    .X(_2568_));
 sky130_fd_sc_hd__mux2_1 _5565_ (.A0(_2568_),
    .A1(\game.padded_notes1[19] ),
    .S(_2472_),
    .X(_2569_));
 sky130_fd_sc_hd__clkbuf_1 _5566_ (.A(_2569_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _5567_ (.A0(\disp_song.note1[20] ),
    .A1(\game.padded_notes1[19] ),
    .S(_2541_),
    .X(_2570_));
 sky130_fd_sc_hd__mux2_1 _5568_ (.A0(_2570_),
    .A1(net222),
    .S(_2472_),
    .X(_2571_));
 sky130_fd_sc_hd__clkbuf_1 _5569_ (.A(_2571_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _5570_ (.A0(\disp_song.note1[21] ),
    .A1(\game.padded_notes1[20] ),
    .S(_2541_),
    .X(_2572_));
 sky130_fd_sc_hd__mux2_1 _5571_ (.A0(_2572_),
    .A1(net225),
    .S(_2472_),
    .X(_2573_));
 sky130_fd_sc_hd__clkbuf_1 _5572_ (.A(_2573_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _5573_ (.A0(\disp_song.note1[22] ),
    .A1(\game.padded_notes1[21] ),
    .S(_2541_),
    .X(_2574_));
 sky130_fd_sc_hd__mux2_1 _5574_ (.A0(_2574_),
    .A1(\game.padded_notes1[22] ),
    .S(_2472_),
    .X(_2575_));
 sky130_fd_sc_hd__clkbuf_1 _5575_ (.A(_2575_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _5576_ (.A0(\disp_song.note1[23] ),
    .A1(\game.padded_notes1[22] ),
    .S(_2541_),
    .X(_2576_));
 sky130_fd_sc_hd__mux2_1 _5577_ (.A0(_2576_),
    .A1(\game.padded_notes1[23] ),
    .S(_2472_),
    .X(_2577_));
 sky130_fd_sc_hd__clkbuf_1 _5578_ (.A(_2577_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _5579_ (.A0(\disp_song.note1[24] ),
    .A1(\game.padded_notes1[23] ),
    .S(_2541_),
    .X(_2578_));
 sky130_fd_sc_hd__mux2_1 _5580_ (.A0(_2578_),
    .A1(net210),
    .S(_2472_),
    .X(_2579_));
 sky130_fd_sc_hd__clkbuf_1 _5581_ (.A(_2579_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _5582_ (.A0(\disp_song.note1[25] ),
    .A1(\game.padded_notes1[24] ),
    .S(_2541_),
    .X(_2580_));
 sky130_fd_sc_hd__mux2_1 _5583_ (.A0(_2580_),
    .A1(net217),
    .S(_2472_),
    .X(_2581_));
 sky130_fd_sc_hd__clkbuf_1 _5584_ (.A(_2581_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _5585_ (.A0(\disp_song.note1[26] ),
    .A1(\game.padded_notes1[25] ),
    .S(_0209_),
    .X(_2582_));
 sky130_fd_sc_hd__mux2_1 _5586_ (.A0(_2582_),
    .A1(\game.padded_notes1[26] ),
    .S(_2472_),
    .X(_2583_));
 sky130_fd_sc_hd__clkbuf_1 _5587_ (.A(_2583_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _5588_ (.A0(\disp_song.note1[27] ),
    .A1(\game.padded_notes1[26] ),
    .S(_0209_),
    .X(_2584_));
 sky130_fd_sc_hd__mux2_1 _5589_ (.A0(_2584_),
    .A1(\game.padded_notes1[27] ),
    .S(_2472_),
    .X(_2585_));
 sky130_fd_sc_hd__clkbuf_1 _5590_ (.A(_2585_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _5591_ (.A0(\disp_song.note1[28] ),
    .A1(\game.padded_notes1[27] ),
    .S(_0209_),
    .X(_2586_));
 sky130_fd_sc_hd__mux2_1 _5592_ (.A0(_2586_),
    .A1(net212),
    .S(_2472_),
    .X(_2587_));
 sky130_fd_sc_hd__clkbuf_1 _5593_ (.A(_2587_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _5594_ (.A0(\disp_song.note1[29] ),
    .A1(\game.padded_notes1[28] ),
    .S(_0209_),
    .X(_2588_));
 sky130_fd_sc_hd__mux2_1 _5595_ (.A0(_2588_),
    .A1(net223),
    .S(_2472_),
    .X(_2589_));
 sky130_fd_sc_hd__clkbuf_1 _5596_ (.A(_2589_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _5597_ (.A0(\disp_song.note1[30] ),
    .A1(\game.padded_notes1[29] ),
    .S(_0209_),
    .X(_2590_));
 sky130_fd_sc_hd__mux2_1 _5598_ (.A0(_2590_),
    .A1(\game.padded_notes1[30] ),
    .S(_2472_),
    .X(_2591_));
 sky130_fd_sc_hd__clkbuf_1 _5599_ (.A(_2591_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _5600_ (.A0(\disp_song.note1[31] ),
    .A1(\game.padded_notes1[30] ),
    .S(_0209_),
    .X(_2592_));
 sky130_fd_sc_hd__mux2_1 _5601_ (.A0(_2592_),
    .A1(\game.padded_notes1[31] ),
    .S(_2472_),
    .X(_2593_));
 sky130_fd_sc_hd__clkbuf_1 _5602_ (.A(_2593_),
    .X(_0121_));
 sky130_fd_sc_hd__a22o_1 _5603_ (.A1(\game.padded_notes1[31] ),
    .A2(_2460_),
    .B1(_2462_),
    .B2(net138),
    .X(_0122_));
 sky130_fd_sc_hd__a22o_1 _5604_ (.A1(\game.out[0] ),
    .A2(_2460_),
    .B1(_2462_),
    .B2(net119),
    .X(_0123_));
 sky130_fd_sc_hd__a22o_1 _5605_ (.A1(net119),
    .A2(_2460_),
    .B1(_2462_),
    .B2(net101),
    .X(_0124_));
 sky130_fd_sc_hd__a22o_1 _5606_ (.A1(net101),
    .A2(_2460_),
    .B1(_2462_),
    .B2(\game.out[3] ),
    .X(_0125_));
 sky130_fd_sc_hd__a22o_1 _5607_ (.A1(\game.out[3] ),
    .A2(_2460_),
    .B1(_2462_),
    .B2(net115),
    .X(_0126_));
 sky130_fd_sc_hd__a22o_1 _5608_ (.A1(net115),
    .A2(_2460_),
    .B1(_2462_),
    .B2(net127),
    .X(_0127_));
 sky130_fd_sc_hd__a22o_1 _5609_ (.A1(\game.out[5] ),
    .A2(_2460_),
    .B1(_2462_),
    .B2(net93),
    .X(_0128_));
 sky130_fd_sc_hd__xnor2_1 _5610_ (.A(net124),
    .B(_0830_),
    .Y(_0129_));
 sky130_fd_sc_hd__and3_1 _5611_ (.A(\game.flash_counter[1] ),
    .B(\game.flash_counter[0] ),
    .C(_0842_),
    .X(_2594_));
 sky130_fd_sc_hd__clkbuf_2 _5612_ (.A(_2594_),
    .X(_2595_));
 sky130_fd_sc_hd__a21oi_1 _5613_ (.A1(\game.flash_counter[0] ),
    .A2(_0842_),
    .B1(net99),
    .Y(_2596_));
 sky130_fd_sc_hd__nor2_1 _5614_ (.A(_2595_),
    .B(net100),
    .Y(_0130_));
 sky130_fd_sc_hd__xor2_1 _5615_ (.A(net113),
    .B(_2595_),
    .X(_0131_));
 sky130_fd_sc_hd__and3_1 _5616_ (.A(\game.flash_counter[3] ),
    .B(\game.flash_counter[2] ),
    .C(_2595_),
    .X(_2597_));
 sky130_fd_sc_hd__a21o_1 _5617_ (.A1(\game.flash_counter[2] ),
    .A2(_2595_),
    .B1(\game.flash_counter[3] ),
    .X(_2598_));
 sky130_fd_sc_hd__and2b_1 _5618_ (.A_N(_2597_),
    .B(_2598_),
    .X(_2599_));
 sky130_fd_sc_hd__clkbuf_1 _5619_ (.A(_2599_),
    .X(_0132_));
 sky130_fd_sc_hd__nand2_1 _5620_ (.A(_0868_),
    .B(_2595_),
    .Y(_2600_));
 sky130_fd_sc_hd__o21a_1 _5621_ (.A1(net96),
    .A2(_2597_),
    .B1(_2600_),
    .X(_0133_));
 sky130_fd_sc_hd__xnor2_1 _5622_ (.A(net146),
    .B(_2600_),
    .Y(_0134_));
 sky130_fd_sc_hd__and2_1 _5623_ (.A(_0868_),
    .B(_2595_),
    .X(_2601_));
 sky130_fd_sc_hd__nand2_1 _5624_ (.A(\game.flash_counter[5] ),
    .B(_2601_),
    .Y(_2602_));
 sky130_fd_sc_hd__xnor2_1 _5625_ (.A(net142),
    .B(_2602_),
    .Y(_0135_));
 sky130_fd_sc_hd__a31oi_1 _5626_ (.A1(\game.flash_counter[6] ),
    .A2(\game.flash_counter[5] ),
    .A3(_2601_),
    .B1(\game.flash_counter[7] ),
    .Y(_2603_));
 sky130_fd_sc_hd__or2b_1 _5627_ (.A(\game.flash_counter[21] ),
    .B_N(\game.flash_counter[20] ),
    .X(_2604_));
 sky130_fd_sc_hd__or4b_1 _5628_ (.A(\game.flash_counter[22] ),
    .B(\game.flash_counter[17] ),
    .C(\game.flash_counter[16] ),
    .D_N(\game.flash_counter[23] ),
    .X(_2605_));
 sky130_fd_sc_hd__or4bb_1 _5629_ (.A(\game.flash_counter[8] ),
    .B(\game.flash_counter[7] ),
    .C_N(\game.flash_counter[6] ),
    .D_N(\game.flash_counter[9] ),
    .X(_2606_));
 sky130_fd_sc_hd__or4bb_1 _5630_ (.A(\game.flash_counter[13] ),
    .B(\game.flash_counter[11] ),
    .C_N(\game.flash_counter[10] ),
    .D_N(\game.flash_counter[12] ),
    .X(_2607_));
 sky130_fd_sc_hd__or4bb_1 _5631_ (.A(\game.flash_counter[18] ),
    .B(\game.flash_counter[14] ),
    .C_N(\game.flash_counter[15] ),
    .D_N(\game.flash_counter[19] ),
    .X(_2608_));
 sky130_fd_sc_hd__or3_1 _5632_ (.A(_2606_),
    .B(_2607_),
    .C(_2608_),
    .X(_2609_));
 sky130_fd_sc_hd__nor4_1 _5633_ (.A(_2602_),
    .B(_2604_),
    .C(_2605_),
    .D(_2609_),
    .Y(_2610_));
 sky130_fd_sc_hd__and4_1 _5634_ (.A(\game.flash_counter[6] ),
    .B(\game.flash_counter[7] ),
    .C(\game.flash_counter[5] ),
    .D(_2601_),
    .X(_2611_));
 sky130_fd_sc_hd__clkbuf_2 _5635_ (.A(_2611_),
    .X(_2612_));
 sky130_fd_sc_hd__nor3_1 _5636_ (.A(_2603_),
    .B(net37),
    .C(_2612_),
    .Y(_0136_));
 sky130_fd_sc_hd__xor2_1 _5637_ (.A(net187),
    .B(_2612_),
    .X(_0137_));
 sky130_fd_sc_hd__a21oi_1 _5638_ (.A1(\game.flash_counter[8] ),
    .A2(_2612_),
    .B1(\game.flash_counter[9] ),
    .Y(_2613_));
 sky130_fd_sc_hd__a311oi_1 _5639_ (.A1(net129),
    .A2(\game.flash_counter[8] ),
    .A3(_2612_),
    .B1(_2613_),
    .C1(net37),
    .Y(_0138_));
 sky130_fd_sc_hd__or4_2 _5640_ (.A(_2602_),
    .B(_2604_),
    .C(_2605_),
    .D(_2609_),
    .X(_2614_));
 sky130_fd_sc_hd__a31o_1 _5641_ (.A1(\game.flash_counter[9] ),
    .A2(\game.flash_counter[8] ),
    .A3(_2612_),
    .B1(\game.flash_counter[10] ),
    .X(_2615_));
 sky130_fd_sc_hd__and4_1 _5642_ (.A(\game.flash_counter[10] ),
    .B(\game.flash_counter[9] ),
    .C(\game.flash_counter[8] ),
    .D(_2612_),
    .X(_2616_));
 sky130_fd_sc_hd__inv_2 _5643_ (.A(_2616_),
    .Y(_2617_));
 sky130_fd_sc_hd__and3_1 _5644_ (.A(_2614_),
    .B(_2615_),
    .C(_2617_),
    .X(_2618_));
 sky130_fd_sc_hd__clkbuf_1 _5645_ (.A(_2618_),
    .X(_0139_));
 sky130_fd_sc_hd__xor2_1 _5646_ (.A(net126),
    .B(_2616_),
    .X(_0140_));
 sky130_fd_sc_hd__a21oi_1 _5647_ (.A1(\game.flash_counter[11] ),
    .A2(_2616_),
    .B1(\game.flash_counter[12] ),
    .Y(_2619_));
 sky130_fd_sc_hd__and3_1 _5648_ (.A(\game.flash_counter[10] ),
    .B(\game.flash_counter[6] ),
    .C(\game.flash_counter[7] ),
    .X(_2620_));
 sky130_fd_sc_hd__and3_1 _5649_ (.A(\game.flash_counter[12] ),
    .B(\game.flash_counter[11] ),
    .C(_2620_),
    .X(_2621_));
 sky130_fd_sc_hd__and3_1 _5650_ (.A(_0868_),
    .B(_0870_),
    .C(_2621_),
    .X(_2622_));
 sky130_fd_sc_hd__and2_1 _5651_ (.A(_0842_),
    .B(_2622_),
    .X(_2623_));
 sky130_fd_sc_hd__nor3_1 _5652_ (.A(_2610_),
    .B(_2619_),
    .C(_2623_),
    .Y(_0141_));
 sky130_fd_sc_hd__nand2_1 _5653_ (.A(\game.flash_counter[13] ),
    .B(_2623_),
    .Y(_2624_));
 sky130_fd_sc_hd__or2_1 _5654_ (.A(\game.flash_counter[13] ),
    .B(_2623_),
    .X(_2625_));
 sky130_fd_sc_hd__and2_1 _5655_ (.A(_2624_),
    .B(_2625_),
    .X(_2626_));
 sky130_fd_sc_hd__clkbuf_1 _5656_ (.A(_2626_),
    .X(_0142_));
 sky130_fd_sc_hd__xnor2_1 _5657_ (.A(net121),
    .B(_2624_),
    .Y(_0143_));
 sky130_fd_sc_hd__and3_1 _5658_ (.A(\game.flash_counter[15] ),
    .B(\game.flash_counter[14] ),
    .C(\game.flash_counter[13] ),
    .X(_2627_));
 sky130_fd_sc_hd__and3_1 _5659_ (.A(_0842_),
    .B(_2622_),
    .C(_2627_),
    .X(_2628_));
 sky130_fd_sc_hd__buf_2 _5660_ (.A(_2628_),
    .X(_2629_));
 sky130_fd_sc_hd__a31o_1 _5661_ (.A1(\game.flash_counter[14] ),
    .A2(\game.flash_counter[13] ),
    .A3(_2623_),
    .B1(\game.flash_counter[15] ),
    .X(_2630_));
 sky130_fd_sc_hd__nand2_1 _5662_ (.A(_2614_),
    .B(_2630_),
    .Y(_2631_));
 sky130_fd_sc_hd__nor2_1 _5663_ (.A(_2629_),
    .B(_2631_),
    .Y(_0144_));
 sky130_fd_sc_hd__or2_1 _5664_ (.A(\game.flash_counter[16] ),
    .B(_2629_),
    .X(_2632_));
 sky130_fd_sc_hd__nand2_1 _5665_ (.A(\game.flash_counter[16] ),
    .B(_2629_),
    .Y(_2633_));
 sky130_fd_sc_hd__and2_1 _5666_ (.A(_2632_),
    .B(_2633_),
    .X(_2634_));
 sky130_fd_sc_hd__clkbuf_1 _5667_ (.A(_2634_),
    .X(_0145_));
 sky130_fd_sc_hd__xnor2_1 _5668_ (.A(net137),
    .B(_2633_),
    .Y(_0146_));
 sky130_fd_sc_hd__a31oi_1 _5669_ (.A1(\game.flash_counter[17] ),
    .A2(\game.flash_counter[16] ),
    .A3(_2629_),
    .B1(net263),
    .Y(_2635_));
 sky130_fd_sc_hd__and4_1 _5670_ (.A(\game.flash_counter[18] ),
    .B(\game.flash_counter[17] ),
    .C(\game.flash_counter[16] ),
    .D(_2629_),
    .X(_2636_));
 sky130_fd_sc_hd__nor2_1 _5671_ (.A(net264),
    .B(_2636_),
    .Y(_0147_));
 sky130_fd_sc_hd__or2_1 _5672_ (.A(\game.flash_counter[19] ),
    .B(_2636_),
    .X(_2637_));
 sky130_fd_sc_hd__nand2_1 _5673_ (.A(\game.flash_counter[19] ),
    .B(_2636_),
    .Y(_2638_));
 sky130_fd_sc_hd__and3_1 _5674_ (.A(_2614_),
    .B(_2637_),
    .C(_2638_),
    .X(_2639_));
 sky130_fd_sc_hd__clkbuf_1 _5675_ (.A(_2639_),
    .X(_0148_));
 sky130_fd_sc_hd__and2_1 _5676_ (.A(\game.flash_counter[19] ),
    .B(_2636_),
    .X(_2640_));
 sky130_fd_sc_hd__or2_1 _5677_ (.A(\game.flash_counter[20] ),
    .B(_2640_),
    .X(_2641_));
 sky130_fd_sc_hd__nand2_1 _5678_ (.A(\game.flash_counter[20] ),
    .B(_2640_),
    .Y(_2642_));
 sky130_fd_sc_hd__and3_1 _5679_ (.A(_2614_),
    .B(_2641_),
    .C(_2642_),
    .X(_2643_));
 sky130_fd_sc_hd__clkbuf_1 _5680_ (.A(_2643_),
    .X(_0149_));
 sky130_fd_sc_hd__a2bb2o_1 _5681_ (.A1_N(_2604_),
    .A2_N(_2638_),
    .B1(_2642_),
    .B2(net175),
    .X(_0150_));
 sky130_fd_sc_hd__and4_1 _5682_ (.A(\game.flash_counter[19] ),
    .B(\game.flash_counter[18] ),
    .C(\game.flash_counter[17] ),
    .D(\game.flash_counter[16] ),
    .X(_2644_));
 sky130_fd_sc_hd__and3_1 _5683_ (.A(\game.flash_counter[20] ),
    .B(\game.flash_counter[21] ),
    .C(_2644_),
    .X(_2645_));
 sky130_fd_sc_hd__nand2_1 _5684_ (.A(_2629_),
    .B(_2645_),
    .Y(_2646_));
 sky130_fd_sc_hd__xnor2_1 _5685_ (.A(net125),
    .B(_2646_),
    .Y(_0151_));
 sky130_fd_sc_hd__nand4_1 _5686_ (.A(\game.flash_counter[22] ),
    .B(\game.flash_counter[23] ),
    .C(_2629_),
    .D(_2645_),
    .Y(_2647_));
 sky130_fd_sc_hd__a31o_1 _5687_ (.A1(\game.flash_counter[22] ),
    .A2(_2629_),
    .A3(_2645_),
    .B1(\game.flash_counter[23] ),
    .X(_2648_));
 sky130_fd_sc_hd__and3_1 _5688_ (.A(_2614_),
    .B(_2647_),
    .C(_2648_),
    .X(_2649_));
 sky130_fd_sc_hd__clkbuf_1 _5689_ (.A(_2649_),
    .X(_0152_));
 sky130_fd_sc_hd__and2b_1 _5690_ (.A_N(\disp_song.um.boton2e.edge_2 ),
    .B(\disp_song.um.boton2e.edge_1 ),
    .X(_2650_));
 sky130_fd_sc_hd__mux2_1 _5691_ (.A0(\disp_song.next_red ),
    .A1(\disp_song.next_green ),
    .S(_2650_),
    .X(_2651_));
 sky130_fd_sc_hd__clkbuf_1 _5692_ (.A(_2651_),
    .X(_0153_));
 sky130_fd_sc_hd__or2_1 _5693_ (.A(net203),
    .B(_2530_),
    .X(_2652_));
 sky130_fd_sc_hd__clkbuf_1 _5694_ (.A(_2652_),
    .X(_0154_));
 sky130_fd_sc_hd__and2_1 _5695_ (.A(\game.scoring_button_1.acc[2] ),
    .B(_2529_),
    .X(_2653_));
 sky130_fd_sc_hd__clkbuf_1 _5696_ (.A(_2653_),
    .X(_0155_));
 sky130_fd_sc_hd__dfrtp_1 _5697_ (.CLK(clknet_leaf_0_clk),
    .D(_0033_),
    .RESET_B(net48),
    .Q(\game.scoring_button_2.acc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5698_ (.CLK(clknet_leaf_1_clk),
    .D(_0034_),
    .RESET_B(net48),
    .Q(\game.scoring_button_2.acc[2] ));
 sky130_fd_sc_hd__dfrtp_2 _5699_ (.CLK(clknet_leaf_62_clk),
    .D(_0035_),
    .RESET_B(net53),
    .Q(\highest_score.highest_score[0] ));
 sky130_fd_sc_hd__dfrtp_4 _5700_ (.CLK(clknet_leaf_62_clk),
    .D(_0036_),
    .RESET_B(net53),
    .Q(\highest_score.highest_score[1] ));
 sky130_fd_sc_hd__dfrtp_2 _5701_ (.CLK(clknet_leaf_62_clk),
    .D(_0037_),
    .RESET_B(net53),
    .Q(\highest_score.highest_score[2] ));
 sky130_fd_sc_hd__dfrtp_2 _5702_ (.CLK(clknet_leaf_61_clk),
    .D(_0038_),
    .RESET_B(net53),
    .Q(\highest_score.highest_score[3] ));
 sky130_fd_sc_hd__dfrtp_4 _5703_ (.CLK(clknet_leaf_60_clk),
    .D(_0039_),
    .RESET_B(net50),
    .Q(\highest_score.highest_score[4] ));
 sky130_fd_sc_hd__dfrtp_4 _5704_ (.CLK(clknet_leaf_60_clk),
    .D(_0040_),
    .RESET_B(net50),
    .Q(\highest_score.highest_score[5] ));
 sky130_fd_sc_hd__dfrtp_4 _5705_ (.CLK(clknet_leaf_60_clk),
    .D(_0041_),
    .RESET_B(net50),
    .Q(\highest_score.highest_score[6] ));
 sky130_fd_sc_hd__dfrtp_1 _5706_ (.CLK(clknet_leaf_60_clk),
    .D(_0042_),
    .RESET_B(net51),
    .Q(\highest_score.highest_score[7] ));
 sky130_fd_sc_hd__dfrtp_1 _5707_ (.CLK(clknet_leaf_23_clk),
    .D(net77),
    .RESET_B(net65),
    .Q(\modetrans.u3.Q1 ));
 sky130_fd_sc_hd__dfrtp_1 _5708_ (.CLK(clknet_leaf_43_clk),
    .D(net80),
    .RESET_B(net65),
    .Q(\modetrans.u3.Q2 ));
 sky130_fd_sc_hd__dfrtp_1 _5709_ (.CLK(clknet_leaf_23_clk),
    .D(\modetrans.pushed_4 ),
    .RESET_B(net64),
    .Q(\modetrans.u3.sync_pb ));
 sky130_fd_sc_hd__dfrtp_2 _5710_ (.CLK(clknet_leaf_39_clk),
    .D(net75),
    .RESET_B(net66),
    .Q(\modetrans.u2.Q1 ));
 sky130_fd_sc_hd__dfrtp_1 _5711_ (.CLK(clknet_leaf_23_clk),
    .D(net82),
    .RESET_B(net65),
    .Q(\modetrans.u2.Q2 ));
 sky130_fd_sc_hd__dfrtp_1 _5712_ (.CLK(clknet_leaf_39_clk),
    .D(\modetrans.pushed_3 ),
    .RESET_B(net66),
    .Q(\modetrans.u2.sync_pb ));
 sky130_fd_sc_hd__dfstp_2 _5713_ (.CLK(clknet_leaf_5_clk),
    .D(_0003_),
    .SET_B(net49),
    .Q(\modetrans.mode[0] ));
 sky130_fd_sc_hd__dfrtp_1 _5714_ (.CLK(clknet_leaf_22_clk),
    .D(_0004_),
    .RESET_B(net59),
    .Q(\modetrans.mode[1] ));
 sky130_fd_sc_hd__dfrtp_4 _5715_ (.CLK(clknet_leaf_23_clk),
    .D(_0005_),
    .RESET_B(net65),
    .Q(\modetrans.mode[2] ));
 sky130_fd_sc_hd__dfrtp_4 _5716_ (.CLK(clknet_leaf_22_clk),
    .D(_0006_),
    .RESET_B(net65),
    .Q(\modetrans.mode[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5717_ (.CLK(clknet_leaf_5_clk),
    .D(_0007_),
    .RESET_B(net59),
    .Q(\modetrans.mode[4] ));
 sky130_fd_sc_hd__dfrtp_4 _5718_ (.CLK(clknet_leaf_22_clk),
    .D(_0008_),
    .RESET_B(net59),
    .Q(\modetrans.mode[5] ));
 sky130_fd_sc_hd__dfrtp_1 _5719_ (.CLK(clknet_leaf_7_clk),
    .D(_0043_),
    .RESET_B(net59),
    .Q(\pulseout.fin_pulse[0] ));
 sky130_fd_sc_hd__dfrtp_1 _5720_ (.CLK(clknet_leaf_6_clk),
    .D(_0044_),
    .RESET_B(net59),
    .Q(\pulseout.fin_pulse[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5721_ (.CLK(clknet_leaf_7_clk),
    .D(_0045_),
    .RESET_B(net59),
    .Q(\pulseout.fin_pulse[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5722_ (.CLK(clknet_leaf_6_clk),
    .D(_0046_),
    .RESET_B(net59),
    .Q(\pulseout.fin_pulse[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5723_ (.CLK(clknet_leaf_6_clk),
    .D(_0047_),
    .RESET_B(net59),
    .Q(\pulseout.fin_pulse[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5724_ (.CLK(clknet_leaf_6_clk),
    .D(_0048_),
    .RESET_B(net59),
    .Q(\pulseout.fin_pulse[5] ));
 sky130_fd_sc_hd__dfstp_2 _5725_ (.CLK(clknet_leaf_4_clk),
    .D(_0000_),
    .SET_B(net49),
    .Q(\lvls.level[0] ));
 sky130_fd_sc_hd__dfrtp_4 _5726_ (.CLK(clknet_leaf_4_clk),
    .D(_0001_),
    .RESET_B(net49),
    .Q(\lvls.level[1] ));
 sky130_fd_sc_hd__dfrtp_4 _5727_ (.CLK(clknet_leaf_4_clk),
    .D(_0002_),
    .RESET_B(net49),
    .Q(\lvls.level[2] ));
 sky130_fd_sc_hd__dfrtp_4 _5728_ (.CLK(clknet_leaf_0_clk),
    .D(\game.scoring_button_2.next_num_misses[0] ),
    .RESET_B(net48),
    .Q(\game.addmisses.add1.b[0] ));
 sky130_fd_sc_hd__dfrtp_4 _5729_ (.CLK(clknet_leaf_0_clk),
    .D(\game.scoring_button_2.next_num_misses[1] ),
    .RESET_B(net48),
    .Q(\game.addmisses.add1.b[1] ));
 sky130_fd_sc_hd__dfrtp_2 _5730_ (.CLK(clknet_leaf_73_clk),
    .D(\game.scoring_button_2.next_num_misses[2] ),
    .RESET_B(net48),
    .Q(\game.addmisses.add1.b[2] ));
 sky130_fd_sc_hd__dfrtp_4 _5731_ (.CLK(clknet_leaf_73_clk),
    .D(\game.scoring_button_2.next_num_misses[3] ),
    .RESET_B(net48),
    .Q(\game.addmisses.add1.b[3] ));
 sky130_fd_sc_hd__dfrtp_4 _5732_ (.CLK(clknet_leaf_73_clk),
    .D(\game.scoring_button_2.next_num_misses[4] ),
    .RESET_B(net48),
    .Q(\game.addmisses.add2.b[0] ));
 sky130_fd_sc_hd__dfrtp_4 _5733_ (.CLK(clknet_leaf_72_clk),
    .D(\game.scoring_button_2.next_num_misses[5] ),
    .RESET_B(net48),
    .Q(\game.addmisses.add2.b[1] ));
 sky130_fd_sc_hd__dfrtp_4 _5734_ (.CLK(clknet_leaf_73_clk),
    .D(\game.scoring_button_2.next_num_misses[6] ),
    .RESET_B(net48),
    .Q(\game.addmisses.add2.b[2] ));
 sky130_fd_sc_hd__dfrtp_4 _5735_ (.CLK(clknet_leaf_72_clk),
    .D(\game.scoring_button_2.next_num_misses[7] ),
    .RESET_B(net48),
    .Q(\game.addmisses.add2.b[3] ));
 sky130_fd_sc_hd__dfrtp_4 _5736_ (.CLK(clknet_leaf_70_clk),
    .D(\game.scoring_button_2.next_num_misses[8] ),
    .RESET_B(net46),
    .Q(\game.addmisses.add3.b[0] ));
 sky130_fd_sc_hd__dfrtp_4 _5737_ (.CLK(clknet_leaf_70_clk),
    .D(\game.scoring_button_2.next_num_misses[9] ),
    .RESET_B(net46),
    .Q(\game.addmisses.add3.b[1] ));
 sky130_fd_sc_hd__dfrtp_4 _5738_ (.CLK(clknet_leaf_70_clk),
    .D(\game.scoring_button_2.next_num_misses[10] ),
    .RESET_B(net46),
    .Q(\game.addmisses.add3.b[2] ));
 sky130_fd_sc_hd__dfrtp_2 _5739_ (.CLK(clknet_leaf_70_clk),
    .D(\game.scoring_button_2.next_num_misses[11] ),
    .RESET_B(net46),
    .Q(\game.addmisses.add3.b[3] ));
 sky130_fd_sc_hd__dfrtp_2 _5740_ (.CLK(clknet_leaf_70_clk),
    .D(\game.scoring_button_2.next_num_misses[12] ),
    .RESET_B(net46),
    .Q(\game.addmisses.add4.b[0] ));
 sky130_fd_sc_hd__dfrtp_2 _5741_ (.CLK(clknet_leaf_69_clk),
    .D(\game.scoring_button_2.next_num_misses[13] ),
    .RESET_B(net46),
    .Q(\game.addmisses.add4.b[1] ));
 sky130_fd_sc_hd__dfrtp_4 _5742_ (.CLK(clknet_leaf_69_clk),
    .D(\game.scoring_button_2.next_num_misses[14] ),
    .RESET_B(net46),
    .Q(\game.addmisses.add4.b[2] ));
 sky130_fd_sc_hd__dfrtp_4 _5743_ (.CLK(clknet_leaf_69_clk),
    .D(\game.scoring_button_2.next_num_misses[15] ),
    .RESET_B(net46),
    .Q(\game.addmisses.add4.b[3] ));
 sky130_fd_sc_hd__dfrtp_4 _5744_ (.CLK(clknet_leaf_1_clk),
    .D(\game.scoring_button_2.next_num_hits[0] ),
    .RESET_B(net48),
    .Q(\game.addhits.add1.b[0] ));
 sky130_fd_sc_hd__dfrtp_4 _5745_ (.CLK(clknet_leaf_1_clk),
    .D(\game.scoring_button_2.next_num_hits[1] ),
    .RESET_B(net49),
    .Q(\game.addhits.add1.b[1] ));
 sky130_fd_sc_hd__dfrtp_2 _5746_ (.CLK(clknet_leaf_3_clk),
    .D(\game.scoring_button_2.next_num_hits[2] ),
    .RESET_B(net49),
    .Q(\game.addhits.add1.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5747_ (.CLK(clknet_leaf_3_clk),
    .D(\game.scoring_button_2.next_num_hits[3] ),
    .RESET_B(net49),
    .Q(\game.addhits.add1.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5748_ (.CLK(clknet_leaf_3_clk),
    .D(\game.scoring_button_2.next_num_hits[4] ),
    .RESET_B(net49),
    .Q(\game.addhits.add2.b[0] ));
 sky130_fd_sc_hd__dfrtp_4 _5749_ (.CLK(clknet_leaf_3_clk),
    .D(\game.scoring_button_2.next_num_hits[5] ),
    .RESET_B(net49),
    .Q(\game.addhits.add2.b[1] ));
 sky130_fd_sc_hd__dfrtp_2 _5750_ (.CLK(clknet_leaf_2_clk),
    .D(\game.scoring_button_2.next_num_hits[6] ),
    .RESET_B(net48),
    .Q(\game.addhits.add2.b[2] ));
 sky130_fd_sc_hd__dfrtp_2 _5751_ (.CLK(clknet_leaf_3_clk),
    .D(\game.scoring_button_2.next_num_hits[7] ),
    .RESET_B(net49),
    .Q(\game.addhits.add2.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5752_ (.CLK(clknet_leaf_66_clk),
    .D(\game.scoring_button_2.next_num_hits[8] ),
    .RESET_B(net46),
    .Q(\game.addhits.add3.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _5753_ (.CLK(clknet_leaf_66_clk),
    .D(\game.scoring_button_2.next_num_hits[9] ),
    .RESET_B(net47),
    .Q(\game.addhits.add3.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5754_ (.CLK(clknet_leaf_68_clk),
    .D(\game.scoring_button_2.next_num_hits[10] ),
    .RESET_B(net46),
    .Q(\game.addhits.add3.b[2] ));
 sky130_fd_sc_hd__dfrtp_2 _5755_ (.CLK(clknet_leaf_68_clk),
    .D(\game.scoring_button_2.next_num_hits[11] ),
    .RESET_B(net46),
    .Q(\game.addhits.add3.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5756_ (.CLK(clknet_leaf_65_clk),
    .D(\game.scoring_button_2.next_num_hits[12] ),
    .RESET_B(net47),
    .Q(\game.addhits.add4.b[0] ));
 sky130_fd_sc_hd__dfrtp_2 _5757_ (.CLK(clknet_leaf_64_clk),
    .D(\game.scoring_button_2.next_num_hits[13] ),
    .RESET_B(net47),
    .Q(\game.addhits.add4.b[1] ));
 sky130_fd_sc_hd__dfrtp_2 _5758_ (.CLK(clknet_leaf_65_clk),
    .D(\game.scoring_button_2.next_num_hits[14] ),
    .RESET_B(net47),
    .Q(\game.addhits.add4.b[2] ));
 sky130_fd_sc_hd__dfrtp_4 _5759_ (.CLK(clknet_leaf_64_clk),
    .D(\game.scoring_button_2.next_num_hits[15] ),
    .RESET_B(net47),
    .Q(\game.addhits.add4.b[3] ));
 sky130_fd_sc_hd__dfrtp_4 _5760_ (.CLK(clknet_leaf_47_clk),
    .D(\game.scoring_button_2.next_missed ),
    .RESET_B(net56),
    .Q(\game.missed_2 ));
 sky130_fd_sc_hd__dfrtp_4 _5761_ (.CLK(clknet_leaf_62_clk),
    .D(\game.scoring_button_2.next_good ),
    .RESET_B(net53),
    .Q(\game.hit_2 ));
 sky130_fd_sc_hd__dfrtp_1 _5762_ (.CLK(clknet_leaf_0_clk),
    .D(net132),
    .RESET_B(net48),
    .Q(\game.scoring_button_2.hit ));
 sky130_fd_sc_hd__dfrtp_1 _5763_ (.CLK(clknet_leaf_16_clk),
    .D(\game.scoring_button_2.next_count[0] ),
    .RESET_B(net62),
    .Q(\game.scoring_button_2.counts[0] ));
 sky130_fd_sc_hd__dfrtp_1 _5764_ (.CLK(clknet_leaf_16_clk),
    .D(\game.scoring_button_2.next_count[1] ),
    .RESET_B(net62),
    .Q(\game.scoring_button_2.counts[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5765_ (.CLK(clknet_leaf_16_clk),
    .D(\game.scoring_button_2.next_count[2] ),
    .RESET_B(net62),
    .Q(\game.scoring_button_2.counts[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5766_ (.CLK(clknet_leaf_16_clk),
    .D(\game.scoring_button_2.next_count[3] ),
    .RESET_B(net62),
    .Q(\game.scoring_button_2.counts[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5767_ (.CLK(clknet_leaf_15_clk),
    .D(\game.scoring_button_2.next_count[4] ),
    .RESET_B(net62),
    .Q(\game.scoring_button_2.counts[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5768_ (.CLK(clknet_leaf_17_clk),
    .D(\game.scoring_button_2.next_count[5] ),
    .RESET_B(net62),
    .Q(\game.scoring_button_2.counts[5] ));
 sky130_fd_sc_hd__dfrtp_1 _5769_ (.CLK(clknet_leaf_17_clk),
    .D(\game.scoring_button_2.next_count[6] ),
    .RESET_B(net62),
    .Q(\game.scoring_button_2.counts[6] ));
 sky130_fd_sc_hd__dfrtp_1 _5770_ (.CLK(clknet_leaf_11_clk),
    .D(\game.scoring_button_2.next_count[7] ),
    .RESET_B(net57),
    .Q(\game.scoring_button_2.counts[7] ));
 sky130_fd_sc_hd__dfrtp_1 _5771_ (.CLK(clknet_leaf_10_clk),
    .D(\game.scoring_button_2.next_count[8] ),
    .RESET_B(net57),
    .Q(\game.scoring_button_2.counts[8] ));
 sky130_fd_sc_hd__dfrtp_1 _5772_ (.CLK(clknet_leaf_10_clk),
    .D(\game.scoring_button_2.next_count[9] ),
    .RESET_B(net57),
    .Q(\game.scoring_button_2.counts[9] ));
 sky130_fd_sc_hd__dfrtp_1 _5773_ (.CLK(clknet_leaf_10_clk),
    .D(\game.scoring_button_2.next_count[10] ),
    .RESET_B(net57),
    .Q(\game.scoring_button_2.counts[10] ));
 sky130_fd_sc_hd__dfrtp_1 _5774_ (.CLK(clknet_leaf_7_clk),
    .D(\game.scoring_button_2.next_count[11] ),
    .RESET_B(net57),
    .Q(\game.scoring_button_2.counts[11] ));
 sky130_fd_sc_hd__dfrtp_1 _5775_ (.CLK(clknet_leaf_7_clk),
    .D(\game.scoring_button_2.next_count[12] ),
    .RESET_B(net59),
    .Q(\game.scoring_button_2.counts[12] ));
 sky130_fd_sc_hd__dfrtp_1 _5776_ (.CLK(clknet_leaf_7_clk),
    .D(\game.scoring_button_2.next_count[13] ),
    .RESET_B(net59),
    .Q(\game.scoring_button_2.counts[13] ));
 sky130_fd_sc_hd__dfrtp_1 _5777_ (.CLK(clknet_leaf_7_clk),
    .D(\game.scoring_button_2.next_count[14] ),
    .RESET_B(net59),
    .Q(\game.scoring_button_2.counts[14] ));
 sky130_fd_sc_hd__dfrtp_1 _5778_ (.CLK(clknet_leaf_11_clk),
    .D(\game.scoring_button_2.next_count[15] ),
    .RESET_B(net57),
    .Q(\game.scoring_button_2.counts[15] ));
 sky130_fd_sc_hd__dfrtp_1 _5779_ (.CLK(clknet_leaf_11_clk),
    .D(\game.scoring_button_2.next_count[16] ),
    .RESET_B(net57),
    .Q(\game.scoring_button_2.counts[16] ));
 sky130_fd_sc_hd__dfrtp_1 _5780_ (.CLK(clknet_leaf_11_clk),
    .D(\game.scoring_button_2.next_count[17] ),
    .RESET_B(net57),
    .Q(\game.scoring_button_2.counts[17] ));
 sky130_fd_sc_hd__dfrtp_1 _5781_ (.CLK(clknet_leaf_11_clk),
    .D(\game.scoring_button_2.next_count[18] ),
    .RESET_B(net57),
    .Q(\game.scoring_button_2.counts[18] ));
 sky130_fd_sc_hd__dfrtp_1 _5782_ (.CLK(clknet_leaf_11_clk),
    .D(\game.scoring_button_2.next_count[19] ),
    .RESET_B(net57),
    .Q(\game.scoring_button_2.counts[19] ));
 sky130_fd_sc_hd__dfrtp_1 _5783_ (.CLK(clknet_leaf_11_clk),
    .D(\game.scoring_button_2.next_count[20] ),
    .RESET_B(net57),
    .Q(\game.scoring_button_2.counts[20] ));
 sky130_fd_sc_hd__dfrtp_1 _5784_ (.CLK(clknet_leaf_11_clk),
    .D(\game.scoring_button_2.next_count[21] ),
    .RESET_B(net57),
    .Q(\game.scoring_button_2.counts[21] ));
 sky130_fd_sc_hd__dfrtp_1 _5785_ (.CLK(clknet_leaf_11_clk),
    .D(\game.scoring_button_2.next_count[22] ),
    .RESET_B(net57),
    .Q(\game.scoring_button_2.counts[22] ));
 sky130_fd_sc_hd__dfrtp_2 _5786_ (.CLK(clknet_leaf_55_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[0] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _5787_ (.CLK(clknet_leaf_55_clk),
    .D(net104),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5788_ (.CLK(clknet_leaf_55_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[2] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5789_ (.CLK(clknet_leaf_54_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[3] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5790_ (.CLK(clknet_leaf_54_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[4] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5791_ (.CLK(clknet_leaf_54_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[5] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _5792_ (.CLK(clknet_leaf_55_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[6] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _5793_ (.CLK(clknet_leaf_53_clk),
    .D(net193),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _5794_ (.CLK(clknet_leaf_53_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[8] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _5795_ (.CLK(clknet_leaf_53_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[9] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _5796_ (.CLK(clknet_leaf_53_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[10] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _5797_ (.CLK(clknet_leaf_53_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[11] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _5798_ (.CLK(clknet_leaf_53_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[12] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _5799_ (.CLK(clknet_leaf_56_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[13] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _5800_ (.CLK(clknet_leaf_55_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[14] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _5801_ (.CLK(clknet_leaf_55_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[15] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _5802_ (.CLK(clknet_leaf_56_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[16] ),
    .RESET_B(net51),
    .Q(\game.scoring_button_2.flash_counter_1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _5803_ (.CLK(clknet_leaf_56_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[17] ),
    .RESET_B(net51),
    .Q(\game.scoring_button_2.flash_counter_1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _5804_ (.CLK(clknet_leaf_56_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[18] ),
    .RESET_B(net51),
    .Q(\game.scoring_button_2.flash_counter_1[18] ));
 sky130_fd_sc_hd__dfrtp_1 _5805_ (.CLK(clknet_leaf_57_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[19] ),
    .RESET_B(net50),
    .Q(\game.scoring_button_2.flash_counter_1[19] ));
 sky130_fd_sc_hd__dfrtp_1 _5806_ (.CLK(clknet_leaf_55_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[20] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[20] ));
 sky130_fd_sc_hd__dfrtp_1 _5807_ (.CLK(clknet_leaf_55_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[21] ),
    .RESET_B(net52),
    .Q(\game.scoring_button_2.flash_counter_1[21] ));
 sky130_fd_sc_hd__dfrtp_1 _5808_ (.CLK(clknet_leaf_55_clk),
    .D(\game.scoring_button_2.next_flash_counter_1[22] ),
    .RESET_B(net73),
    .Q(\game.scoring_button_2.flash_counter_1[22] ));
 sky130_fd_sc_hd__dfrtp_2 _5809_ (.CLK(clknet_leaf_47_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[0] ),
    .RESET_B(net56),
    .Q(\game.scoring_button_2.flash_counter_2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _5810_ (.CLK(clknet_leaf_47_clk),
    .D(net108),
    .RESET_B(net55),
    .Q(\game.scoring_button_2.flash_counter_2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5811_ (.CLK(clknet_leaf_47_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[2] ),
    .RESET_B(net56),
    .Q(\game.scoring_button_2.flash_counter_2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5812_ (.CLK(clknet_leaf_47_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[3] ),
    .RESET_B(net56),
    .Q(\game.scoring_button_2.flash_counter_2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5813_ (.CLK(clknet_leaf_48_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[4] ),
    .RESET_B(net56),
    .Q(\game.scoring_button_2.flash_counter_2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5814_ (.CLK(clknet_leaf_50_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[5] ),
    .RESET_B(net56),
    .Q(\game.scoring_button_2.flash_counter_2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _5815_ (.CLK(clknet_leaf_49_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[6] ),
    .RESET_B(net56),
    .Q(\game.scoring_button_2.flash_counter_2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _5816_ (.CLK(clknet_leaf_49_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[7] ),
    .RESET_B(net56),
    .Q(\game.scoring_button_2.flash_counter_2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _5817_ (.CLK(clknet_leaf_50_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[8] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_2.flash_counter_2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _5818_ (.CLK(clknet_leaf_50_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[9] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_2.flash_counter_2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _5819_ (.CLK(clknet_leaf_50_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[10] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_2.flash_counter_2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _5820_ (.CLK(clknet_leaf_50_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[11] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_2.flash_counter_2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _5821_ (.CLK(clknet_leaf_51_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[12] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_2.flash_counter_2[12] ));
 sky130_fd_sc_hd__dfrtp_1 _5822_ (.CLK(clknet_leaf_51_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[13] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_2.flash_counter_2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _5823_ (.CLK(clknet_leaf_51_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[14] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_2.flash_counter_2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _5824_ (.CLK(clknet_leaf_51_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[15] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_2.flash_counter_2[15] ));
 sky130_fd_sc_hd__dfrtp_1 _5825_ (.CLK(clknet_leaf_52_clk),
    .D(net186),
    .RESET_B(net55),
    .Q(\game.scoring_button_2.flash_counter_2[16] ));
 sky130_fd_sc_hd__dfrtp_1 _5826_ (.CLK(clknet_leaf_52_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[17] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_2.flash_counter_2[17] ));
 sky130_fd_sc_hd__dfrtp_1 _5827_ (.CLK(clknet_leaf_50_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[18] ),
    .RESET_B(net56),
    .Q(\game.scoring_button_2.flash_counter_2[18] ));
 sky130_fd_sc_hd__dfrtp_1 _5828_ (.CLK(clknet_leaf_50_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[19] ),
    .RESET_B(net56),
    .Q(\game.scoring_button_2.flash_counter_2[19] ));
 sky130_fd_sc_hd__dfrtp_1 _5829_ (.CLK(clknet_leaf_52_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[20] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_2.flash_counter_2[20] ));
 sky130_fd_sc_hd__dfrtp_1 _5830_ (.CLK(clknet_leaf_46_clk),
    .D(\game.scoring_button_2.next_flash_counter_2[21] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_2.flash_counter_2[21] ));
 sky130_fd_sc_hd__dfrtp_1 _5831_ (.CLK(clknet_leaf_52_clk),
    .D(net88),
    .RESET_B(net55),
    .Q(\game.scoring_button_2.flash_counter_2[22] ));
 sky130_fd_sc_hd__dfrtp_4 _5832_ (.CLK(clknet_leaf_10_clk),
    .D(\game.scoring_button_2.next_start_count ),
    .RESET_B(net57),
    .Q(\game.scoring_button_2.check_hit.in ));
 sky130_fd_sc_hd__dfrtp_1 _5833_ (.CLK(clknet_leaf_0_clk),
    .D(net84),
    .RESET_B(net48),
    .Q(\game.scoring_button_2.check_hit.edge_2 ));
 sky130_fd_sc_hd__dfrtp_1 _5834_ (.CLK(clknet_leaf_11_clk),
    .D(net90),
    .RESET_B(net57),
    .Q(\game.scoring_button_2.check_hit.edge_1 ));
 sky130_fd_sc_hd__dfrtp_4 _5835_ (.CLK(clknet_leaf_0_clk),
    .D(\game.scoring_button_1.next_num_misses[0] ),
    .RESET_B(net49),
    .Q(\game.addmisses.a[0] ));
 sky130_fd_sc_hd__dfrtp_4 _5836_ (.CLK(clknet_leaf_0_clk),
    .D(\game.scoring_button_1.next_num_misses[1] ),
    .RESET_B(net49),
    .Q(\game.addmisses.a[1] ));
 sky130_fd_sc_hd__dfrtp_2 _5837_ (.CLK(clknet_leaf_73_clk),
    .D(\game.scoring_button_1.next_num_misses[2] ),
    .RESET_B(net49),
    .Q(\game.addmisses.a[2] ));
 sky130_fd_sc_hd__dfrtp_4 _5838_ (.CLK(clknet_leaf_2_clk),
    .D(\game.scoring_button_1.next_num_misses[3] ),
    .RESET_B(net49),
    .Q(\game.addmisses.a[3] ));
 sky130_fd_sc_hd__dfrtp_4 _5839_ (.CLK(clknet_leaf_2_clk),
    .D(\game.scoring_button_1.next_num_misses[4] ),
    .RESET_B(net48),
    .Q(\game.addmisses.a[4] ));
 sky130_fd_sc_hd__dfrtp_4 _5840_ (.CLK(clknet_leaf_71_clk),
    .D(\game.scoring_button_1.next_num_misses[5] ),
    .RESET_B(net48),
    .Q(\game.addmisses.a[5] ));
 sky130_fd_sc_hd__dfrtp_4 _5841_ (.CLK(clknet_leaf_73_clk),
    .D(\game.scoring_button_1.next_num_misses[6] ),
    .RESET_B(net48),
    .Q(\game.addmisses.a[6] ));
 sky130_fd_sc_hd__dfrtp_4 _5842_ (.CLK(clknet_leaf_72_clk),
    .D(\game.scoring_button_1.next_num_misses[7] ),
    .RESET_B(net48),
    .Q(\game.addmisses.a[7] ));
 sky130_fd_sc_hd__dfrtp_4 _5843_ (.CLK(clknet_leaf_72_clk),
    .D(\game.scoring_button_1.next_num_misses[8] ),
    .RESET_B(net48),
    .Q(\game.addmisses.a[8] ));
 sky130_fd_sc_hd__dfrtp_4 _5844_ (.CLK(clknet_leaf_70_clk),
    .D(\game.scoring_button_1.next_num_misses[9] ),
    .RESET_B(net46),
    .Q(\game.addmisses.a[9] ));
 sky130_fd_sc_hd__dfrtp_4 _5845_ (.CLK(clknet_leaf_71_clk),
    .D(\game.scoring_button_1.next_num_misses[10] ),
    .RESET_B(net46),
    .Q(\game.addmisses.a[10] ));
 sky130_fd_sc_hd__dfrtp_2 _5846_ (.CLK(clknet_leaf_71_clk),
    .D(\game.scoring_button_1.next_num_misses[11] ),
    .RESET_B(net46),
    .Q(\game.addmisses.a[11] ));
 sky130_fd_sc_hd__dfrtp_2 _5847_ (.CLK(clknet_3_0__leaf_clk),
    .D(\game.scoring_button_1.next_num_misses[12] ),
    .RESET_B(net46),
    .Q(\game.addmisses.a[12] ));
 sky130_fd_sc_hd__dfrtp_2 _5848_ (.CLK(clknet_leaf_69_clk),
    .D(\game.scoring_button_1.next_num_misses[13] ),
    .RESET_B(net46),
    .Q(\game.addmisses.a[13] ));
 sky130_fd_sc_hd__dfrtp_4 _5849_ (.CLK(clknet_leaf_69_clk),
    .D(\game.scoring_button_1.next_num_misses[14] ),
    .RESET_B(net46),
    .Q(\game.addmisses.a[14] ));
 sky130_fd_sc_hd__dfrtp_4 _5850_ (.CLK(clknet_leaf_68_clk),
    .D(\game.scoring_button_1.next_num_misses[15] ),
    .RESET_B(net46),
    .Q(\game.addmisses.a[15] ));
 sky130_fd_sc_hd__dfrtp_4 _5851_ (.CLK(clknet_leaf_4_clk),
    .D(\game.scoring_button_1.next_num_hits[0] ),
    .RESET_B(net49),
    .Q(\game.addhits.a[0] ));
 sky130_fd_sc_hd__dfrtp_4 _5852_ (.CLK(clknet_leaf_4_clk),
    .D(\game.scoring_button_1.next_num_hits[1] ),
    .RESET_B(net49),
    .Q(\game.addhits.a[1] ));
 sky130_fd_sc_hd__dfrtp_2 _5853_ (.CLK(clknet_leaf_4_clk),
    .D(\game.scoring_button_1.next_num_hits[2] ),
    .RESET_B(net49),
    .Q(\game.addhits.a[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5854_ (.CLK(clknet_leaf_4_clk),
    .D(\game.scoring_button_1.next_num_hits[3] ),
    .RESET_B(net49),
    .Q(\game.addhits.a[3] ));
 sky130_fd_sc_hd__dfrtp_2 _5855_ (.CLK(clknet_3_1__leaf_clk),
    .D(\game.scoring_button_1.next_num_hits[4] ),
    .RESET_B(net48),
    .Q(\game.addhits.a[4] ));
 sky130_fd_sc_hd__dfrtp_4 _5856_ (.CLK(clknet_leaf_66_clk),
    .D(\game.scoring_button_1.next_num_hits[5] ),
    .RESET_B(net47),
    .Q(\game.addhits.a[5] ));
 sky130_fd_sc_hd__dfrtp_2 _5857_ (.CLK(clknet_leaf_71_clk),
    .D(\game.scoring_button_1.next_num_hits[6] ),
    .RESET_B(net46),
    .Q(\game.addhits.a[6] ));
 sky130_fd_sc_hd__dfrtp_2 _5858_ (.CLK(clknet_leaf_66_clk),
    .D(\game.scoring_button_1.next_num_hits[7] ),
    .RESET_B(net46),
    .Q(\game.addhits.a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _5859_ (.CLK(clknet_leaf_66_clk),
    .D(\game.scoring_button_1.next_num_hits[8] ),
    .RESET_B(net47),
    .Q(\game.addhits.a[8] ));
 sky130_fd_sc_hd__dfrtp_1 _5860_ (.CLK(clknet_leaf_65_clk),
    .D(\game.scoring_button_1.next_num_hits[9] ),
    .RESET_B(net47),
    .Q(\game.addhits.a[9] ));
 sky130_fd_sc_hd__dfrtp_2 _5861_ (.CLK(clknet_leaf_65_clk),
    .D(\game.scoring_button_1.next_num_hits[10] ),
    .RESET_B(net47),
    .Q(\game.addhits.a[10] ));
 sky130_fd_sc_hd__dfrtp_2 _5862_ (.CLK(clknet_leaf_65_clk),
    .D(\game.scoring_button_1.next_num_hits[11] ),
    .RESET_B(net47),
    .Q(\game.addhits.a[11] ));
 sky130_fd_sc_hd__dfrtp_1 _5863_ (.CLK(clknet_leaf_65_clk),
    .D(\game.scoring_button_1.next_num_hits[12] ),
    .RESET_B(net47),
    .Q(\game.addhits.a[12] ));
 sky130_fd_sc_hd__dfrtp_2 _5864_ (.CLK(clknet_leaf_59_clk),
    .D(\game.scoring_button_1.next_num_hits[13] ),
    .RESET_B(net47),
    .Q(\game.addhits.a[13] ));
 sky130_fd_sc_hd__dfrtp_2 _5865_ (.CLK(clknet_leaf_64_clk),
    .D(\game.scoring_button_1.next_num_hits[14] ),
    .RESET_B(net47),
    .Q(\game.addhits.a[14] ));
 sky130_fd_sc_hd__dfrtp_4 _5866_ (.CLK(clknet_leaf_64_clk),
    .D(\game.scoring_button_1.next_num_hits[15] ),
    .RESET_B(net50),
    .Q(\game.addhits.a[15] ));
 sky130_fd_sc_hd__dfrtp_1 _5867_ (.CLK(clknet_leaf_23_clk),
    .D(net92),
    .RESET_B(net64),
    .Q(\game.padded_notes2[0] ));
 sky130_fd_sc_hd__dfstp_1 _5868_ (.CLK(clknet_leaf_22_clk),
    .D(_0051_),
    .SET_B(net65),
    .Q(\game.padded_notes2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5869_ (.CLK(clknet_leaf_22_clk),
    .D(_0052_),
    .RESET_B(net59),
    .Q(\game.padded_notes2[2] ));
 sky130_fd_sc_hd__dfstp_1 _5870_ (.CLK(clknet_leaf_22_clk),
    .D(_0053_),
    .SET_B(net60),
    .Q(\game.padded_notes2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5871_ (.CLK(clknet_leaf_22_clk),
    .D(_0054_),
    .RESET_B(net64),
    .Q(\game.padded_notes2[4] ));
 sky130_fd_sc_hd__dfstp_1 _5872_ (.CLK(clknet_leaf_29_clk),
    .D(_0055_),
    .SET_B(net69),
    .Q(\game.padded_notes2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _5873_ (.CLK(clknet_leaf_20_clk),
    .D(_0056_),
    .RESET_B(net63),
    .Q(\game.padded_notes2[6] ));
 sky130_fd_sc_hd__dfstp_1 _5874_ (.CLK(clknet_leaf_19_clk),
    .D(_0057_),
    .SET_B(net63),
    .Q(\game.padded_notes2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _5875_ (.CLK(clknet_leaf_19_clk),
    .D(_0058_),
    .RESET_B(net63),
    .Q(\game.padded_notes2[8] ));
 sky130_fd_sc_hd__dfstp_1 _5876_ (.CLK(clknet_leaf_19_clk),
    .D(_0059_),
    .SET_B(net63),
    .Q(\game.padded_notes2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _5877_ (.CLK(clknet_leaf_19_clk),
    .D(_0060_),
    .RESET_B(net63),
    .Q(\game.padded_notes2[10] ));
 sky130_fd_sc_hd__dfstp_1 _5878_ (.CLK(clknet_leaf_19_clk),
    .D(_0061_),
    .SET_B(net63),
    .Q(\game.padded_notes2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _5879_ (.CLK(clknet_leaf_19_clk),
    .D(_0062_),
    .RESET_B(net63),
    .Q(\game.padded_notes2[12] ));
 sky130_fd_sc_hd__dfstp_1 _5880_ (.CLK(clknet_leaf_20_clk),
    .D(_0063_),
    .SET_B(net63),
    .Q(\game.padded_notes2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _5881_ (.CLK(clknet_leaf_20_clk),
    .D(_0064_),
    .RESET_B(net69),
    .Q(\game.padded_notes2[14] ));
 sky130_fd_sc_hd__dfstp_1 _5882_ (.CLK(clknet_leaf_30_clk),
    .D(_0065_),
    .SET_B(net69),
    .Q(\game.padded_notes2[15] ));
 sky130_fd_sc_hd__dfrtp_1 _5883_ (.CLK(clknet_leaf_30_clk),
    .D(_0066_),
    .RESET_B(net69),
    .Q(\game.padded_notes2[16] ));
 sky130_fd_sc_hd__dfstp_1 _5884_ (.CLK(clknet_leaf_29_clk),
    .D(_0067_),
    .SET_B(net69),
    .Q(\game.padded_notes2[17] ));
 sky130_fd_sc_hd__dfrtp_1 _5885_ (.CLK(clknet_leaf_29_clk),
    .D(_0068_),
    .RESET_B(net69),
    .Q(\game.padded_notes2[18] ));
 sky130_fd_sc_hd__dfstp_1 _5886_ (.CLK(clknet_leaf_30_clk),
    .D(_0069_),
    .SET_B(net69),
    .Q(\game.padded_notes2[19] ));
 sky130_fd_sc_hd__dfrtp_1 _5887_ (.CLK(clknet_leaf_30_clk),
    .D(_0070_),
    .RESET_B(net69),
    .Q(\game.padded_notes2[20] ));
 sky130_fd_sc_hd__dfstp_1 _5888_ (.CLK(clknet_leaf_30_clk),
    .D(_0071_),
    .SET_B(net69),
    .Q(\game.padded_notes2[21] ));
 sky130_fd_sc_hd__dfrtp_1 _5889_ (.CLK(clknet_leaf_31_clk),
    .D(_0072_),
    .RESET_B(net69),
    .Q(\game.padded_notes2[22] ));
 sky130_fd_sc_hd__dfstp_1 _5890_ (.CLK(clknet_leaf_32_clk),
    .D(_0073_),
    .SET_B(net69),
    .Q(\game.padded_notes2[23] ));
 sky130_fd_sc_hd__dfrtp_1 _5891_ (.CLK(clknet_leaf_27_clk),
    .D(_0074_),
    .RESET_B(net68),
    .Q(\game.padded_notes2[24] ));
 sky130_fd_sc_hd__dfstp_1 _5892_ (.CLK(clknet_leaf_26_clk),
    .D(_0075_),
    .SET_B(net68),
    .Q(\game.padded_notes2[25] ));
 sky130_fd_sc_hd__dfrtp_1 _5893_ (.CLK(clknet_leaf_26_clk),
    .D(_0076_),
    .RESET_B(net68),
    .Q(\game.padded_notes2[26] ));
 sky130_fd_sc_hd__dfstp_1 _5894_ (.CLK(clknet_leaf_32_clk),
    .D(_0077_),
    .SET_B(net68),
    .Q(\game.padded_notes2[27] ));
 sky130_fd_sc_hd__dfrtp_1 _5895_ (.CLK(clknet_leaf_32_clk),
    .D(_0078_),
    .RESET_B(net68),
    .Q(\game.padded_notes2[28] ));
 sky130_fd_sc_hd__dfstp_1 _5896_ (.CLK(clknet_leaf_32_clk),
    .D(_0079_),
    .SET_B(net68),
    .Q(\game.padded_notes2[29] ));
 sky130_fd_sc_hd__dfrtp_1 _5897_ (.CLK(clknet_leaf_31_clk),
    .D(_0080_),
    .RESET_B(net69),
    .Q(\game.padded_notes2[30] ));
 sky130_fd_sc_hd__dfstp_1 _5898_ (.CLK(clknet_leaf_26_clk),
    .D(_0081_),
    .SET_B(net68),
    .Q(\game.padded_notes2[31] ));
 sky130_fd_sc_hd__dfrtp_1 _5899_ (.CLK(clknet_leaf_44_clk),
    .D(net134),
    .RESET_B(net53),
    .Q(\game.out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _5900_ (.CLK(clknet_leaf_44_clk),
    .D(_0083_),
    .RESET_B(net53),
    .Q(\game.out[8] ));
 sky130_fd_sc_hd__dfrtp_1 _5901_ (.CLK(clknet_leaf_44_clk),
    .D(net141),
    .RESET_B(net53),
    .Q(\game.out[9] ));
 sky130_fd_sc_hd__dfrtp_1 _5902_ (.CLK(clknet_leaf_44_clk),
    .D(_0085_),
    .RESET_B(net53),
    .Q(\game.out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _5903_ (.CLK(clknet_leaf_44_clk),
    .D(net118),
    .RESET_B(net53),
    .Q(\game.out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _5904_ (.CLK(clknet_leaf_44_clk),
    .D(net136),
    .RESET_B(net54),
    .Q(\game.out[12] ));
 sky130_fd_sc_hd__dfrtp_1 _5905_ (.CLK(clknet_leaf_44_clk),
    .D(_0088_),
    .RESET_B(net54),
    .Q(\game.out[13] ));
 sky130_fd_sc_hd__dfrtp_4 _5906_ (.CLK(clknet_leaf_25_clk),
    .D(\game.scoring_button_1.next_missed ),
    .RESET_B(net64),
    .Q(\game.missed_1 ));
 sky130_fd_sc_hd__dfrtp_4 _5907_ (.CLK(clknet_leaf_45_clk),
    .D(\game.scoring_button_1.next_good ),
    .RESET_B(net54),
    .Q(\game.hit_1 ));
 sky130_fd_sc_hd__dfrtp_2 _5908_ (.CLK(clknet_leaf_10_clk),
    .D(_0089_),
    .RESET_B(net57),
    .Q(\game.scoring_button_1.hit ));
 sky130_fd_sc_hd__dfrtp_1 _5909_ (.CLK(clknet_leaf_15_clk),
    .D(\game.scoring_button_1.next_count[0] ),
    .RESET_B(net62),
    .Q(\game.scoring_button_1.counts[0] ));
 sky130_fd_sc_hd__dfrtp_1 _5910_ (.CLK(clknet_leaf_16_clk),
    .D(\game.scoring_button_1.next_count[1] ),
    .RESET_B(net62),
    .Q(\game.scoring_button_1.counts[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5911_ (.CLK(clknet_leaf_16_clk),
    .D(\game.scoring_button_1.next_count[2] ),
    .RESET_B(net62),
    .Q(\game.scoring_button_1.counts[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5912_ (.CLK(clknet_leaf_16_clk),
    .D(\game.scoring_button_1.next_count[3] ),
    .RESET_B(net62),
    .Q(\game.scoring_button_1.counts[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5913_ (.CLK(clknet_leaf_15_clk),
    .D(\game.scoring_button_1.next_count[4] ),
    .RESET_B(net62),
    .Q(\game.scoring_button_1.counts[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5914_ (.CLK(clknet_leaf_15_clk),
    .D(\game.scoring_button_1.next_count[5] ),
    .RESET_B(net62),
    .Q(\game.scoring_button_1.counts[5] ));
 sky130_fd_sc_hd__dfrtp_1 _5915_ (.CLK(clknet_leaf_17_clk),
    .D(\game.scoring_button_1.next_count[6] ),
    .RESET_B(net62),
    .Q(\game.scoring_button_1.counts[6] ));
 sky130_fd_sc_hd__dfrtp_1 _5916_ (.CLK(clknet_leaf_14_clk),
    .D(\game.scoring_button_1.next_count[7] ),
    .RESET_B(net58),
    .Q(\game.scoring_button_1.counts[7] ));
 sky130_fd_sc_hd__dfrtp_1 _5917_ (.CLK(clknet_leaf_15_clk),
    .D(\game.scoring_button_1.next_count[8] ),
    .RESET_B(net58),
    .Q(\game.scoring_button_1.counts[8] ));
 sky130_fd_sc_hd__dfrtp_1 _5918_ (.CLK(clknet_leaf_15_clk),
    .D(\game.scoring_button_1.next_count[9] ),
    .RESET_B(net62),
    .Q(\game.scoring_button_1.counts[9] ));
 sky130_fd_sc_hd__dfrtp_1 _5919_ (.CLK(clknet_leaf_21_clk),
    .D(\game.scoring_button_1.next_count[10] ),
    .RESET_B(net60),
    .Q(\game.scoring_button_1.counts[10] ));
 sky130_fd_sc_hd__dfrtp_1 _5920_ (.CLK(clknet_leaf_9_clk),
    .D(\game.scoring_button_1.next_count[11] ),
    .RESET_B(net60),
    .Q(\game.scoring_button_1.counts[11] ));
 sky130_fd_sc_hd__dfrtp_1 _5921_ (.CLK(clknet_leaf_8_clk),
    .D(\game.scoring_button_1.next_count[12] ),
    .RESET_B(net60),
    .Q(\game.scoring_button_1.counts[12] ));
 sky130_fd_sc_hd__dfrtp_1 _5922_ (.CLK(clknet_leaf_8_clk),
    .D(\game.scoring_button_1.next_count[13] ),
    .RESET_B(net60),
    .Q(\game.scoring_button_1.counts[13] ));
 sky130_fd_sc_hd__dfrtp_1 _5923_ (.CLK(clknet_leaf_8_clk),
    .D(\game.scoring_button_1.next_count[14] ),
    .RESET_B(net60),
    .Q(\game.scoring_button_1.counts[14] ));
 sky130_fd_sc_hd__dfrtp_1 _5924_ (.CLK(clknet_leaf_13_clk),
    .D(\game.scoring_button_1.next_count[15] ),
    .RESET_B(net58),
    .Q(\game.scoring_button_1.counts[15] ));
 sky130_fd_sc_hd__dfrtp_1 _5925_ (.CLK(clknet_leaf_13_clk),
    .D(\game.scoring_button_1.next_count[16] ),
    .RESET_B(net58),
    .Q(\game.scoring_button_1.counts[16] ));
 sky130_fd_sc_hd__dfrtp_1 _5926_ (.CLK(clknet_leaf_13_clk),
    .D(\game.scoring_button_1.next_count[17] ),
    .RESET_B(net58),
    .Q(\game.scoring_button_1.counts[17] ));
 sky130_fd_sc_hd__dfrtp_1 _5927_ (.CLK(clknet_leaf_13_clk),
    .D(\game.scoring_button_1.next_count[18] ),
    .RESET_B(net58),
    .Q(\game.scoring_button_1.counts[18] ));
 sky130_fd_sc_hd__dfrtp_1 _5928_ (.CLK(clknet_leaf_12_clk),
    .D(\game.scoring_button_1.next_count[19] ),
    .RESET_B(net58),
    .Q(\game.scoring_button_1.counts[19] ));
 sky130_fd_sc_hd__dfrtp_1 _5929_ (.CLK(clknet_leaf_12_clk),
    .D(\game.scoring_button_1.next_count[20] ),
    .RESET_B(net58),
    .Q(\game.scoring_button_1.counts[20] ));
 sky130_fd_sc_hd__dfrtp_1 _5930_ (.CLK(clknet_leaf_13_clk),
    .D(\game.scoring_button_1.next_count[21] ),
    .RESET_B(net58),
    .Q(\game.scoring_button_1.counts[21] ));
 sky130_fd_sc_hd__dfrtp_1 _5931_ (.CLK(clknet_leaf_13_clk),
    .D(\game.scoring_button_1.next_count[22] ),
    .RESET_B(net58),
    .Q(\game.scoring_button_1.counts[22] ));
 sky130_fd_sc_hd__dfrtp_2 _5932_ (.CLK(clknet_leaf_61_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[0] ),
    .RESET_B(net53),
    .Q(\game.scoring_button_1.flash_counter_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _5933_ (.CLK(clknet_leaf_60_clk),
    .D(net112),
    .RESET_B(net51),
    .Q(\game.scoring_button_1.flash_counter_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5934_ (.CLK(clknet_leaf_60_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[2] ),
    .RESET_B(net51),
    .Q(\game.scoring_button_1.flash_counter_1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5935_ (.CLK(clknet_leaf_60_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[3] ),
    .RESET_B(net51),
    .Q(\game.scoring_button_1.flash_counter_1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5936_ (.CLK(clknet_leaf_56_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[4] ),
    .RESET_B(net51),
    .Q(\game.scoring_button_1.flash_counter_1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5937_ (.CLK(clknet_leaf_61_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[5] ),
    .RESET_B(net53),
    .Q(\game.scoring_button_1.flash_counter_1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _5938_ (.CLK(clknet_leaf_56_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[6] ),
    .RESET_B(net73),
    .Q(\game.scoring_button_1.flash_counter_1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _5939_ (.CLK(clknet_leaf_52_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[7] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_1.flash_counter_1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _5940_ (.CLK(clknet_leaf_46_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[8] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_1.flash_counter_1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _5941_ (.CLK(clknet_leaf_52_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[9] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_1.flash_counter_1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _5942_ (.CLK(clknet_leaf_46_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[10] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_1.flash_counter_1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _5943_ (.CLK(clknet_leaf_52_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[11] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_1.flash_counter_1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _5944_ (.CLK(clknet_leaf_46_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[12] ),
    .RESET_B(net55),
    .Q(\game.scoring_button_1.flash_counter_1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _5945_ (.CLK(clknet_leaf_47_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[13] ),
    .RESET_B(net56),
    .Q(\game.scoring_button_1.flash_counter_1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _5946_ (.CLK(clknet_leaf_45_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[14] ),
    .RESET_B(net53),
    .Q(\game.scoring_button_1.flash_counter_1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _5947_ (.CLK(clknet_leaf_45_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[15] ),
    .RESET_B(net54),
    .Q(\game.scoring_button_1.flash_counter_1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _5948_ (.CLK(clknet_leaf_45_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[16] ),
    .RESET_B(net54),
    .Q(\game.scoring_button_1.flash_counter_1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _5949_ (.CLK(clknet_leaf_45_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[17] ),
    .RESET_B(net53),
    .Q(\game.scoring_button_1.flash_counter_1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _5950_ (.CLK(clknet_leaf_61_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[18] ),
    .RESET_B(net53),
    .Q(\game.scoring_button_1.flash_counter_1[18] ));
 sky130_fd_sc_hd__dfrtp_1 _5951_ (.CLK(clknet_leaf_61_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[19] ),
    .RESET_B(net53),
    .Q(\game.scoring_button_1.flash_counter_1[19] ));
 sky130_fd_sc_hd__dfrtp_1 _5952_ (.CLK(clknet_leaf_45_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[20] ),
    .RESET_B(net53),
    .Q(\game.scoring_button_1.flash_counter_1[20] ));
 sky130_fd_sc_hd__dfrtp_1 _5953_ (.CLK(clknet_leaf_45_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[21] ),
    .RESET_B(net53),
    .Q(\game.scoring_button_1.flash_counter_1[21] ));
 sky130_fd_sc_hd__dfrtp_1 _5954_ (.CLK(clknet_leaf_61_clk),
    .D(\game.scoring_button_1.next_flash_counter_1[22] ),
    .RESET_B(net53),
    .Q(\game.scoring_button_1.flash_counter_1[22] ));
 sky130_fd_sc_hd__dfrtp_2 _5955_ (.CLK(clknet_leaf_33_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[0] ),
    .RESET_B(net71),
    .Q(\game.scoring_button_1.flash_counter_2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _5956_ (.CLK(clknet_leaf_34_clk),
    .D(net106),
    .RESET_B(net71),
    .Q(\game.scoring_button_1.flash_counter_2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5957_ (.CLK(clknet_leaf_34_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[2] ),
    .RESET_B(net72),
    .Q(\game.scoring_button_1.flash_counter_2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5958_ (.CLK(clknet_leaf_36_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[3] ),
    .RESET_B(net72),
    .Q(\game.scoring_button_1.flash_counter_2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5959_ (.CLK(clknet_leaf_36_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[4] ),
    .RESET_B(net72),
    .Q(\game.scoring_button_1.flash_counter_2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5960_ (.CLK(clknet_leaf_36_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[5] ),
    .RESET_B(net72),
    .Q(\game.scoring_button_1.flash_counter_2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _5961_ (.CLK(clknet_leaf_34_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[6] ),
    .RESET_B(net72),
    .Q(\game.scoring_button_1.flash_counter_2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _5962_ (.CLK(clknet_leaf_36_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[7] ),
    .RESET_B(net72),
    .Q(\game.scoring_button_1.flash_counter_2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _5963_ (.CLK(clknet_leaf_35_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[8] ),
    .RESET_B(net72),
    .Q(\game.scoring_button_1.flash_counter_2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _5964_ (.CLK(clknet_leaf_34_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[9] ),
    .RESET_B(net72),
    .Q(\game.scoring_button_1.flash_counter_2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _5965_ (.CLK(clknet_leaf_35_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[10] ),
    .RESET_B(net72),
    .Q(\game.scoring_button_1.flash_counter_2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _5966_ (.CLK(clknet_leaf_35_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[11] ),
    .RESET_B(net72),
    .Q(\game.scoring_button_1.flash_counter_2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _5967_ (.CLK(clknet_leaf_35_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[12] ),
    .RESET_B(net72),
    .Q(\game.scoring_button_1.flash_counter_2[12] ));
 sky130_fd_sc_hd__dfrtp_1 _5968_ (.CLK(clknet_leaf_31_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[13] ),
    .RESET_B(net69),
    .Q(\game.scoring_button_1.flash_counter_2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _5969_ (.CLK(clknet_leaf_31_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[14] ),
    .RESET_B(net69),
    .Q(\game.scoring_button_1.flash_counter_2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _5970_ (.CLK(clknet_leaf_31_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[15] ),
    .RESET_B(net70),
    .Q(\game.scoring_button_1.flash_counter_2[15] ));
 sky130_fd_sc_hd__dfrtp_1 _5971_ (.CLK(clknet_leaf_31_clk),
    .D(net195),
    .RESET_B(net70),
    .Q(\game.scoring_button_1.flash_counter_2[16] ));
 sky130_fd_sc_hd__dfrtp_1 _5972_ (.CLK(clknet_leaf_31_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[17] ),
    .RESET_B(net72),
    .Q(\game.scoring_button_1.flash_counter_2[17] ));
 sky130_fd_sc_hd__dfrtp_1 _5973_ (.CLK(clknet_leaf_31_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[18] ),
    .RESET_B(net70),
    .Q(\game.scoring_button_1.flash_counter_2[18] ));
 sky130_fd_sc_hd__dfrtp_1 _5974_ (.CLK(clknet_leaf_32_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[19] ),
    .RESET_B(net71),
    .Q(\game.scoring_button_1.flash_counter_2[19] ));
 sky130_fd_sc_hd__dfrtp_1 _5975_ (.CLK(clknet_leaf_34_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[20] ),
    .RESET_B(net72),
    .Q(\game.scoring_button_1.flash_counter_2[20] ));
 sky130_fd_sc_hd__dfrtp_1 _5976_ (.CLK(clknet_leaf_33_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[21] ),
    .RESET_B(net71),
    .Q(\game.scoring_button_1.flash_counter_2[21] ));
 sky130_fd_sc_hd__dfrtp_1 _5977_ (.CLK(clknet_leaf_34_clk),
    .D(\game.scoring_button_1.next_flash_counter_2[22] ),
    .RESET_B(net71),
    .Q(\game.scoring_button_1.flash_counter_2[22] ));
 sky130_fd_sc_hd__dfrtp_4 _5978_ (.CLK(clknet_leaf_10_clk),
    .D(\game.scoring_button_1.next_start_count ),
    .RESET_B(net57),
    .Q(\game.scoring_button_1.check_hit.in ));
 sky130_fd_sc_hd__dfrtp_1 _5979_ (.CLK(clknet_leaf_10_clk),
    .D(net81),
    .RESET_B(net61),
    .Q(\game.scoring_button_1.check_hit.edge_2 ));
 sky130_fd_sc_hd__dfrtp_1 _5980_ (.CLK(clknet_leaf_11_clk),
    .D(net95),
    .RESET_B(net61),
    .Q(\game.scoring_button_1.check_hit.edge_1 ));
 sky130_fd_sc_hd__dfrtp_1 _5981_ (.CLK(clknet_leaf_25_clk),
    .D(net98),
    .RESET_B(net64),
    .Q(\game.padded_notes1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _5982_ (.CLK(clknet_leaf_26_clk),
    .D(_0091_),
    .RESET_B(net68),
    .Q(\game.padded_notes1[1] ));
 sky130_fd_sc_hd__dfstp_1 _5983_ (.CLK(clknet_leaf_26_clk),
    .D(_0092_),
    .SET_B(net68),
    .Q(\game.padded_notes1[2] ));
 sky130_fd_sc_hd__dfstp_1 _5984_ (.CLK(clknet_leaf_33_clk),
    .D(_0093_),
    .SET_B(net68),
    .Q(\game.padded_notes1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5985_ (.CLK(clknet_leaf_32_clk),
    .D(_0094_),
    .RESET_B(net71),
    .Q(\game.padded_notes1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5986_ (.CLK(clknet_leaf_33_clk),
    .D(_0095_),
    .RESET_B(net71),
    .Q(\game.padded_notes1[5] ));
 sky130_fd_sc_hd__dfstp_1 _5987_ (.CLK(clknet_leaf_37_clk),
    .D(_0096_),
    .SET_B(net71),
    .Q(\game.padded_notes1[6] ));
 sky130_fd_sc_hd__dfstp_1 _5988_ (.CLK(clknet_leaf_33_clk),
    .D(_0097_),
    .SET_B(net71),
    .Q(\game.padded_notes1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _5989_ (.CLK(clknet_leaf_33_clk),
    .D(_0098_),
    .RESET_B(net71),
    .Q(\game.padded_notes1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _5990_ (.CLK(clknet_leaf_33_clk),
    .D(_0099_),
    .RESET_B(net71),
    .Q(\game.padded_notes1[9] ));
 sky130_fd_sc_hd__dfstp_1 _5991_ (.CLK(clknet_leaf_37_clk),
    .D(_0100_),
    .SET_B(net71),
    .Q(\game.padded_notes1[10] ));
 sky130_fd_sc_hd__dfstp_1 _5992_ (.CLK(clknet_leaf_37_clk),
    .D(_0101_),
    .SET_B(net71),
    .Q(\game.padded_notes1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _5993_ (.CLK(clknet_leaf_37_clk),
    .D(_0102_),
    .RESET_B(net71),
    .Q(\game.padded_notes1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _5994_ (.CLK(clknet_leaf_37_clk),
    .D(_0103_),
    .RESET_B(net71),
    .Q(\game.padded_notes1[13] ));
 sky130_fd_sc_hd__dfstp_1 _5995_ (.CLK(clknet_leaf_37_clk),
    .D(_0104_),
    .SET_B(net71),
    .Q(\game.padded_notes1[14] ));
 sky130_fd_sc_hd__dfstp_1 _5996_ (.CLK(clknet_leaf_38_clk),
    .D(_0105_),
    .SET_B(net66),
    .Q(\game.padded_notes1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _5997_ (.CLK(clknet_leaf_38_clk),
    .D(_0106_),
    .RESET_B(net66),
    .Q(\game.padded_notes1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _5998_ (.CLK(clknet_leaf_38_clk),
    .D(_0107_),
    .RESET_B(net66),
    .Q(\game.padded_notes1[17] ));
 sky130_fd_sc_hd__dfstp_1 _5999_ (.CLK(clknet_leaf_38_clk),
    .D(_0108_),
    .SET_B(net66),
    .Q(\game.padded_notes1[18] ));
 sky130_fd_sc_hd__dfstp_1 _6000_ (.CLK(clknet_leaf_38_clk),
    .D(_0109_),
    .SET_B(net66),
    .Q(\game.padded_notes1[19] ));
 sky130_fd_sc_hd__dfrtp_1 _6001_ (.CLK(clknet_leaf_38_clk),
    .D(_0110_),
    .RESET_B(net67),
    .Q(\game.padded_notes1[20] ));
 sky130_fd_sc_hd__dfrtp_1 _6002_ (.CLK(clknet_leaf_39_clk),
    .D(_0111_),
    .RESET_B(net67),
    .Q(\game.padded_notes1[21] ));
 sky130_fd_sc_hd__dfstp_1 _6003_ (.CLK(clknet_leaf_38_clk),
    .D(_0112_),
    .SET_B(net66),
    .Q(\game.padded_notes1[22] ));
 sky130_fd_sc_hd__dfstp_1 _6004_ (.CLK(clknet_leaf_39_clk),
    .D(_0113_),
    .SET_B(net66),
    .Q(\game.padded_notes1[23] ));
 sky130_fd_sc_hd__dfrtp_1 _6005_ (.CLK(clknet_leaf_39_clk),
    .D(_0114_),
    .RESET_B(net66),
    .Q(\game.padded_notes1[24] ));
 sky130_fd_sc_hd__dfrtp_1 _6006_ (.CLK(clknet_leaf_39_clk),
    .D(_0115_),
    .RESET_B(net66),
    .Q(\game.padded_notes1[25] ));
 sky130_fd_sc_hd__dfstp_1 _6007_ (.CLK(clknet_leaf_49_clk),
    .D(_0116_),
    .SET_B(net66),
    .Q(\game.padded_notes1[26] ));
 sky130_fd_sc_hd__dfstp_1 _6008_ (.CLK(clknet_leaf_49_clk),
    .D(_0117_),
    .SET_B(net56),
    .Q(\game.padded_notes1[27] ));
 sky130_fd_sc_hd__dfrtp_1 _6009_ (.CLK(clknet_leaf_49_clk),
    .D(_0118_),
    .RESET_B(net56),
    .Q(\game.padded_notes1[28] ));
 sky130_fd_sc_hd__dfrtp_1 _6010_ (.CLK(clknet_leaf_48_clk),
    .D(_0119_),
    .RESET_B(net56),
    .Q(\game.padded_notes1[29] ));
 sky130_fd_sc_hd__dfstp_1 _6011_ (.CLK(clknet_leaf_48_clk),
    .D(_0120_),
    .SET_B(net56),
    .Q(\game.padded_notes1[30] ));
 sky130_fd_sc_hd__dfstp_1 _6012_ (.CLK(clknet_leaf_43_clk),
    .D(_0121_),
    .SET_B(net65),
    .Q(\game.padded_notes1[31] ));
 sky130_fd_sc_hd__dfrtp_1 _6013_ (.CLK(clknet_leaf_22_clk),
    .D(net139),
    .RESET_B(net59),
    .Q(\game.out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6014_ (.CLK(clknet_leaf_22_clk),
    .D(net120),
    .RESET_B(net59),
    .Q(\game.out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6015_ (.CLK(clknet_leaf_6_clk),
    .D(_0124_),
    .RESET_B(net59),
    .Q(\game.out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6016_ (.CLK(clknet_leaf_5_clk),
    .D(net102),
    .RESET_B(net59),
    .Q(\game.out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6017_ (.CLK(clknet_leaf_5_clk),
    .D(net116),
    .RESET_B(net60),
    .Q(\game.out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6018_ (.CLK(clknet_leaf_5_clk),
    .D(_0127_),
    .RESET_B(net60),
    .Q(\game.out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6019_ (.CLK(clknet_leaf_5_clk),
    .D(net94),
    .RESET_B(net60),
    .Q(\game.out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6020_ (.CLK(clknet_leaf_59_clk),
    .D(_0129_),
    .RESET_B(net51),
    .Q(\game.flash_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6021_ (.CLK(clknet_leaf_59_clk),
    .D(_0130_),
    .RESET_B(net50),
    .Q(\game.flash_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6022_ (.CLK(clknet_leaf_59_clk),
    .D(_0131_),
    .RESET_B(net50),
    .Q(\game.flash_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6023_ (.CLK(clknet_leaf_64_clk),
    .D(_0132_),
    .RESET_B(net50),
    .Q(\game.flash_counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6024_ (.CLK(clknet_leaf_58_clk),
    .D(_0133_),
    .RESET_B(net50),
    .Q(\game.flash_counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6025_ (.CLK(clknet_leaf_58_clk),
    .D(_0134_),
    .RESET_B(net50),
    .Q(\game.flash_counter[5] ));
 sky130_fd_sc_hd__dfrtp_2 _6026_ (.CLK(clknet_leaf_58_clk),
    .D(_0135_),
    .RESET_B(net50),
    .Q(\game.flash_counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6027_ (.CLK(clknet_leaf_59_clk),
    .D(_0136_),
    .RESET_B(net50),
    .Q(\game.flash_counter[7] ));
 sky130_fd_sc_hd__dfrtp_2 _6028_ (.CLK(clknet_leaf_59_clk),
    .D(_0137_),
    .RESET_B(net51),
    .Q(\game.flash_counter[8] ));
 sky130_fd_sc_hd__dfrtp_2 _6029_ (.CLK(clknet_leaf_59_clk),
    .D(net130),
    .RESET_B(net51),
    .Q(\game.flash_counter[9] ));
 sky130_fd_sc_hd__dfrtp_2 _6030_ (.CLK(clknet_leaf_60_clk),
    .D(_0139_),
    .RESET_B(net51),
    .Q(\game.flash_counter[10] ));
 sky130_fd_sc_hd__dfrtp_2 _6031_ (.CLK(clknet_leaf_60_clk),
    .D(_0140_),
    .RESET_B(net51),
    .Q(\game.flash_counter[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6032_ (.CLK(clknet_leaf_60_clk),
    .D(_0141_),
    .RESET_B(net51),
    .Q(\game.flash_counter[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6033_ (.CLK(clknet_leaf_60_clk),
    .D(_0142_),
    .RESET_B(net51),
    .Q(\game.flash_counter[13] ));
 sky130_fd_sc_hd__dfrtp_2 _6034_ (.CLK(clknet_leaf_56_clk),
    .D(_0143_),
    .RESET_B(net51),
    .Q(\game.flash_counter[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6035_ (.CLK(clknet_leaf_57_clk),
    .D(_0144_),
    .RESET_B(net51),
    .Q(\game.flash_counter[15] ));
 sky130_fd_sc_hd__dfrtp_4 _6036_ (.CLK(clknet_leaf_58_clk),
    .D(_0145_),
    .RESET_B(net50),
    .Q(\game.flash_counter[16] ));
 sky130_fd_sc_hd__dfrtp_2 _6037_ (.CLK(clknet_leaf_58_clk),
    .D(_0146_),
    .RESET_B(net50),
    .Q(\game.flash_counter[17] ));
 sky130_fd_sc_hd__dfrtp_1 _6038_ (.CLK(clknet_leaf_57_clk),
    .D(_0147_),
    .RESET_B(net50),
    .Q(\game.flash_counter[18] ));
 sky130_fd_sc_hd__dfrtp_2 _6039_ (.CLK(clknet_leaf_57_clk),
    .D(_0148_),
    .RESET_B(net50),
    .Q(\game.flash_counter[19] ));
 sky130_fd_sc_hd__dfrtp_1 _6040_ (.CLK(clknet_leaf_57_clk),
    .D(_0149_),
    .RESET_B(net50),
    .Q(\game.flash_counter[20] ));
 sky130_fd_sc_hd__dfrtp_1 _6041_ (.CLK(clknet_leaf_57_clk),
    .D(_0150_),
    .RESET_B(net50),
    .Q(\game.flash_counter[21] ));
 sky130_fd_sc_hd__dfrtp_2 _6042_ (.CLK(clknet_leaf_58_clk),
    .D(_0151_),
    .RESET_B(net50),
    .Q(\game.flash_counter[22] ));
 sky130_fd_sc_hd__dfrtp_1 _6043_ (.CLK(clknet_leaf_58_clk),
    .D(_0152_),
    .RESET_B(net50),
    .Q(\game.flash_counter[23] ));
 sky130_fd_sc_hd__dfrtp_2 _6044_ (.CLK(clknet_leaf_13_clk),
    .D(_0009_),
    .RESET_B(net58),
    .Q(\game.counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6045_ (.CLK(clknet_leaf_16_clk),
    .D(_0020_),
    .RESET_B(net62),
    .Q(\game.counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6046_ (.CLK(clknet_leaf_16_clk),
    .D(_0024_),
    .RESET_B(net62),
    .Q(\game.counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6047_ (.CLK(clknet_leaf_16_clk),
    .D(_0025_),
    .RESET_B(net62),
    .Q(\game.counter[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6048_ (.CLK(clknet_leaf_15_clk),
    .D(_0026_),
    .RESET_B(net62),
    .Q(\game.counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6049_ (.CLK(clknet_leaf_15_clk),
    .D(_0027_),
    .RESET_B(net62),
    .Q(\game.counter[5] ));
 sky130_fd_sc_hd__dfrtp_2 _6050_ (.CLK(clknet_leaf_14_clk),
    .D(_0028_),
    .RESET_B(net58),
    .Q(\game.counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6051_ (.CLK(clknet_leaf_14_clk),
    .D(_0029_),
    .RESET_B(net58),
    .Q(\game.counter[7] ));
 sky130_fd_sc_hd__dfrtp_2 _6052_ (.CLK(clknet_leaf_14_clk),
    .D(_0030_),
    .RESET_B(net58),
    .Q(\game.counter[8] ));
 sky130_fd_sc_hd__dfrtp_4 _6053_ (.CLK(clknet_leaf_15_clk),
    .D(_0031_),
    .RESET_B(net63),
    .Q(\game.counter[9] ));
 sky130_fd_sc_hd__dfrtp_1 _6054_ (.CLK(clknet_leaf_8_clk),
    .D(_0010_),
    .RESET_B(net60),
    .Q(\game.counter[10] ));
 sky130_fd_sc_hd__dfrtp_2 _6055_ (.CLK(clknet_leaf_8_clk),
    .D(_0011_),
    .RESET_B(net60),
    .Q(\game.counter[11] ));
 sky130_fd_sc_hd__dfrtp_2 _6056_ (.CLK(clknet_leaf_8_clk),
    .D(_0012_),
    .RESET_B(net60),
    .Q(\game.counter[12] ));
 sky130_fd_sc_hd__dfrtp_1 _6057_ (.CLK(clknet_leaf_7_clk),
    .D(_0013_),
    .RESET_B(net59),
    .Q(\game.counter[13] ));
 sky130_fd_sc_hd__dfrtp_2 _6058_ (.CLK(clknet_leaf_9_clk),
    .D(_0014_),
    .RESET_B(net61),
    .Q(\game.counter[14] ));
 sky130_fd_sc_hd__dfrtp_2 _6059_ (.CLK(clknet_leaf_14_clk),
    .D(_0015_),
    .RESET_B(net61),
    .Q(\game.counter[15] ));
 sky130_fd_sc_hd__dfrtp_4 _6060_ (.CLK(clknet_leaf_12_clk),
    .D(_0016_),
    .RESET_B(net58),
    .Q(\game.counter[16] ));
 sky130_fd_sc_hd__dfrtp_2 _6061_ (.CLK(clknet_leaf_12_clk),
    .D(_0017_),
    .RESET_B(net58),
    .Q(\game.counter[17] ));
 sky130_fd_sc_hd__dfrtp_4 _6062_ (.CLK(clknet_leaf_12_clk),
    .D(_0018_),
    .RESET_B(net58),
    .Q(\game.counter[18] ));
 sky130_fd_sc_hd__dfrtp_1 _6063_ (.CLK(clknet_leaf_12_clk),
    .D(_0019_),
    .RESET_B(net58),
    .Q(\game.counter[19] ));
 sky130_fd_sc_hd__dfrtp_2 _6064_ (.CLK(clknet_leaf_12_clk),
    .D(_0021_),
    .RESET_B(net57),
    .Q(\game.counter[20] ));
 sky130_fd_sc_hd__dfrtp_4 _6065_ (.CLK(clknet_leaf_12_clk),
    .D(_0022_),
    .RESET_B(net57),
    .Q(\game.counter[21] ));
 sky130_fd_sc_hd__dfrtp_2 _6066_ (.CLK(clknet_leaf_12_clk),
    .D(_0023_),
    .RESET_B(net57),
    .Q(\game.counter[22] ));
 sky130_fd_sc_hd__dfrtp_2 _6067_ (.CLK(clknet_leaf_7_clk),
    .D(_0032_),
    .RESET_B(net59),
    .Q(\game.beat_clk ));
 sky130_fd_sc_hd__dfrtp_1 _6068_ (.CLK(clknet_leaf_25_clk),
    .D(_0153_),
    .RESET_B(net64),
    .Q(\disp_song.toggle_state ));
 sky130_fd_sc_hd__dfrtp_1 _6069_ (.CLK(clknet_leaf_62_clk),
    .D(\highest_score.nxt_mode[0] ),
    .RESET_B(net54),
    .Q(\highest_score.score_mode[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6070_ (.CLK(clknet_leaf_62_clk),
    .D(\highest_score.nxt_mode[1] ),
    .RESET_B(net53),
    .Q(\highest_score.score_mode[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6071_ (.CLK(clknet_leaf_10_clk),
    .D(_0154_),
    .RESET_B(net61),
    .Q(\game.scoring_button_1.acc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6072_ (.CLK(clknet_leaf_7_clk),
    .D(_0155_),
    .RESET_B(net59),
    .Q(\game.scoring_button_1.acc[2] ));
 sky130_fd_sc_hd__dfstp_4 _6073_ (.CLK(clknet_leaf_29_clk),
    .D(\disp_song.um.drum.next_idx2[0] ),
    .SET_B(net69),
    .Q(\disp_song.um.idx_note2[0] ));
 sky130_fd_sc_hd__dfstp_4 _6074_ (.CLK(clknet_leaf_28_clk),
    .D(\disp_song.um.drum.next_idx2[1] ),
    .SET_B(net68),
    .Q(\disp_song.um.idx_note2[1] ));
 sky130_fd_sc_hd__dfstp_2 _6075_ (.CLK(clknet_leaf_24_clk),
    .D(\disp_song.um.drum.next_idx2[2] ),
    .SET_B(net64),
    .Q(\disp_song.um.idx_note2[2] ));
 sky130_fd_sc_hd__dfstp_2 _6076_ (.CLK(clknet_leaf_21_clk),
    .D(\disp_song.um.drum.next_idx2[3] ),
    .SET_B(net60),
    .Q(\disp_song.um.idx_note2[3] ));
 sky130_fd_sc_hd__dfstp_2 _6077_ (.CLK(clknet_leaf_24_clk),
    .D(\disp_song.um.drum.next_idx2[4] ),
    .SET_B(net64),
    .Q(\disp_song.um.idx_note2[4] ));
 sky130_fd_sc_hd__dfstp_4 _6078_ (.CLK(clknet_leaf_40_clk),
    .D(\disp_song.um.drum.next_idx1[0] ),
    .SET_B(net66),
    .Q(\disp_song.um.idx_note1[0] ));
 sky130_fd_sc_hd__dfstp_1 _6079_ (.CLK(clknet_leaf_40_clk),
    .D(\disp_song.um.drum.next_idx1[1] ),
    .SET_B(net66),
    .Q(\disp_song.um.idx_note1[1] ));
 sky130_fd_sc_hd__dfstp_4 _6080_ (.CLK(clknet_leaf_43_clk),
    .D(\disp_song.um.drum.next_idx1[2] ),
    .SET_B(net64),
    .Q(\disp_song.um.idx_note1[2] ));
 sky130_fd_sc_hd__dfstp_2 _6081_ (.CLK(clknet_leaf_43_clk),
    .D(\disp_song.um.drum.next_idx1[3] ),
    .SET_B(net65),
    .Q(\disp_song.um.idx_note1[3] ));
 sky130_fd_sc_hd__dfstp_1 _6082_ (.CLK(clknet_leaf_42_clk),
    .D(\disp_song.um.drum.next_idx1[4] ),
    .SET_B(net64),
    .Q(\disp_song.um.idx_note1[4] ));
 sky130_fd_sc_hd__dfstp_1 _6083_ (.CLK(clknet_leaf_23_clk),
    .D(\disp_song.um.next_position[0] ),
    .SET_B(net64),
    .Q(\disp_song.mi6.in[0] ));
 sky130_fd_sc_hd__dfstp_1 _6084_ (.CLK(clknet_leaf_23_clk),
    .D(\disp_song.um.next_position[1] ),
    .SET_B(net65),
    .Q(\disp_song.mi6.in[1] ));
 sky130_fd_sc_hd__dfstp_2 _6085_ (.CLK(clknet_leaf_43_clk),
    .D(\disp_song.um.next_position[2] ),
    .SET_B(net65),
    .Q(\disp_song.mi6.in[2] ));
 sky130_fd_sc_hd__dfstp_4 _6086_ (.CLK(clknet_leaf_23_clk),
    .D(\disp_song.um.next_position[3] ),
    .SET_B(net65),
    .Q(\disp_song.mi6.in[3] ));
 sky130_fd_sc_hd__dfstp_1 _6087_ (.CLK(clknet_leaf_43_clk),
    .D(\disp_song.um.next_position[4] ),
    .SET_B(net65),
    .Q(\disp_song.mi6.in[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6088_ (.CLK(clknet_leaf_23_clk),
    .D(\disp_song.um.drum.next_note1[0] ),
    .RESET_B(net64),
    .Q(\disp_song.note1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6089_ (.CLK(clknet_leaf_43_clk),
    .D(\disp_song.um.drum.next_note1[1] ),
    .RESET_B(net64),
    .Q(\disp_song.note1[1] ));
 sky130_fd_sc_hd__dfstp_2 _6090_ (.CLK(clknet_leaf_42_clk),
    .D(\disp_song.um.drum.next_note1[2] ),
    .SET_B(net64),
    .Q(\disp_song.note1[2] ));
 sky130_fd_sc_hd__dfstp_1 _6091_ (.CLK(clknet_leaf_26_clk),
    .D(\disp_song.um.drum.next_note1[3] ),
    .SET_B(net64),
    .Q(\disp_song.note1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6092_ (.CLK(clknet_leaf_42_clk),
    .D(\disp_song.um.drum.next_note1[4] ),
    .RESET_B(net64),
    .Q(\disp_song.note1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6093_ (.CLK(clknet_leaf_25_clk),
    .D(\disp_song.um.drum.next_note1[5] ),
    .RESET_B(net65),
    .Q(\disp_song.note1[5] ));
 sky130_fd_sc_hd__dfstp_1 _6094_ (.CLK(clknet_leaf_37_clk),
    .D(\disp_song.um.drum.next_note1[6] ),
    .SET_B(net71),
    .Q(\disp_song.note1[6] ));
 sky130_fd_sc_hd__dfstp_1 _6095_ (.CLK(clknet_leaf_37_clk),
    .D(\disp_song.um.drum.next_note1[7] ),
    .SET_B(net71),
    .Q(\disp_song.note1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6096_ (.CLK(clknet_leaf_41_clk),
    .D(\disp_song.um.drum.next_note1[8] ),
    .RESET_B(net67),
    .Q(\disp_song.note1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _6097_ (.CLK(clknet_leaf_37_clk),
    .D(\disp_song.um.drum.next_note1[9] ),
    .RESET_B(net67),
    .Q(\disp_song.note1[9] ));
 sky130_fd_sc_hd__dfstp_1 _6098_ (.CLK(clknet_leaf_37_clk),
    .D(\disp_song.um.drum.next_note1[10] ),
    .SET_B(net71),
    .Q(\disp_song.note1[10] ));
 sky130_fd_sc_hd__dfstp_1 _6099_ (.CLK(clknet_leaf_37_clk),
    .D(\disp_song.um.drum.next_note1[11] ),
    .SET_B(net67),
    .Q(\disp_song.note1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6100_ (.CLK(clknet_leaf_37_clk),
    .D(\disp_song.um.drum.next_note1[12] ),
    .RESET_B(net67),
    .Q(\disp_song.note1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _6101_ (.CLK(clknet_leaf_37_clk),
    .D(\disp_song.um.drum.next_note1[13] ),
    .RESET_B(net71),
    .Q(\disp_song.note1[13] ));
 sky130_fd_sc_hd__dfstp_1 _6102_ (.CLK(clknet_leaf_37_clk),
    .D(\disp_song.um.drum.next_note1[14] ),
    .SET_B(net67),
    .Q(\disp_song.note1[14] ));
 sky130_fd_sc_hd__dfstp_1 _6103_ (.CLK(clknet_leaf_38_clk),
    .D(\disp_song.um.drum.next_note1[15] ),
    .SET_B(net67),
    .Q(\disp_song.note1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6104_ (.CLK(clknet_leaf_25_clk),
    .D(\disp_song.um.drum.next_note1[16] ),
    .RESET_B(net65),
    .Q(\disp_song.note1[16] ));
 sky130_fd_sc_hd__dfrtp_2 _6105_ (.CLK(clknet_leaf_42_clk),
    .D(\disp_song.um.drum.next_note1[17] ),
    .RESET_B(net67),
    .Q(\disp_song.note1[17] ));
 sky130_fd_sc_hd__dfstp_1 _6106_ (.CLK(clknet_leaf_38_clk),
    .D(\disp_song.um.drum.next_note1[18] ),
    .SET_B(net67),
    .Q(\disp_song.note1[18] ));
 sky130_fd_sc_hd__dfstp_1 _6107_ (.CLK(clknet_leaf_41_clk),
    .D(\disp_song.um.drum.next_note1[19] ),
    .SET_B(net67),
    .Q(\disp_song.note1[19] ));
 sky130_fd_sc_hd__dfrtp_1 _6108_ (.CLK(clknet_leaf_41_clk),
    .D(\disp_song.um.drum.next_note1[20] ),
    .RESET_B(net67),
    .Q(\disp_song.note1[20] ));
 sky130_fd_sc_hd__dfrtp_1 _6109_ (.CLK(clknet_leaf_38_clk),
    .D(\disp_song.um.drum.next_note1[21] ),
    .RESET_B(net67),
    .Q(\disp_song.note1[21] ));
 sky130_fd_sc_hd__dfstp_1 _6110_ (.CLK(clknet_leaf_38_clk),
    .D(\disp_song.um.drum.next_note1[22] ),
    .SET_B(net66),
    .Q(\disp_song.note1[22] ));
 sky130_fd_sc_hd__dfstp_1 _6111_ (.CLK(clknet_leaf_40_clk),
    .D(\disp_song.um.drum.next_note1[23] ),
    .SET_B(net66),
    .Q(\disp_song.note1[23] ));
 sky130_fd_sc_hd__dfrtp_1 _6112_ (.CLK(clknet_leaf_41_clk),
    .D(\disp_song.um.drum.next_note1[24] ),
    .RESET_B(net67),
    .Q(\disp_song.note1[24] ));
 sky130_fd_sc_hd__dfrtp_1 _6113_ (.CLK(clknet_leaf_40_clk),
    .D(\disp_song.um.drum.next_note1[25] ),
    .RESET_B(net66),
    .Q(\disp_song.note1[25] ));
 sky130_fd_sc_hd__dfstp_1 _6114_ (.CLK(clknet_leaf_39_clk),
    .D(\disp_song.um.drum.next_note1[26] ),
    .SET_B(net66),
    .Q(\disp_song.note1[26] ));
 sky130_fd_sc_hd__dfstp_1 _6115_ (.CLK(clknet_leaf_40_clk),
    .D(\disp_song.um.drum.next_note1[27] ),
    .SET_B(net66),
    .Q(\disp_song.note1[27] ));
 sky130_fd_sc_hd__dfrtp_1 _6116_ (.CLK(clknet_leaf_48_clk),
    .D(\disp_song.um.drum.next_note1[28] ),
    .RESET_B(net56),
    .Q(\disp_song.note1[28] ));
 sky130_fd_sc_hd__dfrtp_1 _6117_ (.CLK(clknet_leaf_40_clk),
    .D(\disp_song.um.drum.next_note1[29] ),
    .RESET_B(net66),
    .Q(\disp_song.note1[29] ));
 sky130_fd_sc_hd__dfstp_1 _6118_ (.CLK(clknet_leaf_48_clk),
    .D(\disp_song.um.drum.next_note1[30] ),
    .SET_B(net56),
    .Q(\disp_song.note1[30] ));
 sky130_fd_sc_hd__dfstp_1 _6119_ (.CLK(clknet_leaf_48_clk),
    .D(\disp_song.um.drum.next_note1[31] ),
    .SET_B(net56),
    .Q(\disp_song.note1[31] ));
 sky130_fd_sc_hd__dfrtp_1 _6120_ (.CLK(clknet_leaf_23_clk),
    .D(\disp_song.um.drum.next_note2[0] ),
    .RESET_B(net64),
    .Q(\disp_song.note2[0] ));
 sky130_fd_sc_hd__dfstp_1 _6121_ (.CLK(clknet_leaf_22_clk),
    .D(\disp_song.um.drum.next_note2[1] ),
    .SET_B(net60),
    .Q(\disp_song.note2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6122_ (.CLK(clknet_leaf_22_clk),
    .D(\disp_song.um.drum.next_note2[2] ),
    .RESET_B(net60),
    .Q(\disp_song.note2[2] ));
 sky130_fd_sc_hd__dfstp_1 _6123_ (.CLK(clknet_leaf_22_clk),
    .D(\disp_song.um.drum.next_note2[3] ),
    .SET_B(net60),
    .Q(\disp_song.note2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6124_ (.CLK(clknet_leaf_23_clk),
    .D(\disp_song.um.drum.next_note2[4] ),
    .RESET_B(net64),
    .Q(\disp_song.note2[4] ));
 sky130_fd_sc_hd__dfstp_1 _6125_ (.CLK(clknet_leaf_24_clk),
    .D(\disp_song.um.drum.next_note2[5] ),
    .SET_B(net64),
    .Q(\disp_song.note2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6126_ (.CLK(clknet_leaf_20_clk),
    .D(\disp_song.um.drum.next_note2[6] ),
    .RESET_B(net63),
    .Q(\disp_song.note2[6] ));
 sky130_fd_sc_hd__dfstp_1 _6127_ (.CLK(clknet_leaf_20_clk),
    .D(\disp_song.um.drum.next_note2[7] ),
    .SET_B(net63),
    .Q(\disp_song.note2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6128_ (.CLK(clknet_leaf_19_clk),
    .D(\disp_song.um.drum.next_note2[8] ),
    .RESET_B(net63),
    .Q(\disp_song.note2[8] ));
 sky130_fd_sc_hd__dfstp_1 _6129_ (.CLK(clknet_leaf_19_clk),
    .D(\disp_song.um.drum.next_note2[9] ),
    .SET_B(net63),
    .Q(\disp_song.note2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _6130_ (.CLK(clknet_leaf_19_clk),
    .D(\disp_song.um.drum.next_note2[10] ),
    .RESET_B(net63),
    .Q(\disp_song.note2[10] ));
 sky130_fd_sc_hd__dfstp_1 _6131_ (.CLK(clknet_leaf_19_clk),
    .D(\disp_song.um.drum.next_note2[11] ),
    .SET_B(net63),
    .Q(\disp_song.note2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6132_ (.CLK(clknet_leaf_20_clk),
    .D(\disp_song.um.drum.next_note2[12] ),
    .RESET_B(net63),
    .Q(\disp_song.note2[12] ));
 sky130_fd_sc_hd__dfstp_1 _6133_ (.CLK(clknet_leaf_19_clk),
    .D(\disp_song.um.drum.next_note2[13] ),
    .SET_B(net63),
    .Q(\disp_song.note2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6134_ (.CLK(clknet_leaf_20_clk),
    .D(\disp_song.um.drum.next_note2[14] ),
    .RESET_B(net63),
    .Q(\disp_song.note2[14] ));
 sky130_fd_sc_hd__dfstp_1 _6135_ (.CLK(clknet_leaf_29_clk),
    .D(\disp_song.um.drum.next_note2[15] ),
    .SET_B(net69),
    .Q(\disp_song.note2[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6136_ (.CLK(clknet_leaf_25_clk),
    .D(\disp_song.um.drum.next_note2[16] ),
    .RESET_B(net64),
    .Q(\disp_song.note2[16] ));
 sky130_fd_sc_hd__dfstp_1 _6137_ (.CLK(clknet_leaf_28_clk),
    .D(\disp_song.um.drum.next_note2[17] ),
    .SET_B(net68),
    .Q(\disp_song.note2[17] ));
 sky130_fd_sc_hd__dfrtp_1 _6138_ (.CLK(clknet_leaf_29_clk),
    .D(\disp_song.um.drum.next_note2[18] ),
    .RESET_B(net69),
    .Q(\disp_song.note2[18] ));
 sky130_fd_sc_hd__dfstp_1 _6139_ (.CLK(clknet_leaf_28_clk),
    .D(\disp_song.um.drum.next_note2[19] ),
    .SET_B(net68),
    .Q(\disp_song.note2[19] ));
 sky130_fd_sc_hd__dfrtp_1 _6140_ (.CLK(clknet_leaf_28_clk),
    .D(\disp_song.um.drum.next_note2[20] ),
    .RESET_B(net68),
    .Q(\disp_song.note2[20] ));
 sky130_fd_sc_hd__dfstp_1 _6141_ (.CLK(clknet_leaf_30_clk),
    .D(\disp_song.um.drum.next_note2[21] ),
    .SET_B(net69),
    .Q(\disp_song.note2[21] ));
 sky130_fd_sc_hd__dfrtp_1 _6142_ (.CLK(clknet_leaf_30_clk),
    .D(\disp_song.um.drum.next_note2[22] ),
    .RESET_B(net70),
    .Q(\disp_song.note2[22] ));
 sky130_fd_sc_hd__dfstp_1 _6143_ (.CLK(clknet_leaf_30_clk),
    .D(\disp_song.um.drum.next_note2[23] ),
    .SET_B(net69),
    .Q(\disp_song.note2[23] ));
 sky130_fd_sc_hd__dfrtp_1 _6144_ (.CLK(clknet_leaf_28_clk),
    .D(\disp_song.um.drum.next_note2[24] ),
    .RESET_B(net68),
    .Q(\disp_song.note2[24] ));
 sky130_fd_sc_hd__dfstp_1 _6145_ (.CLK(clknet_leaf_27_clk),
    .D(\disp_song.um.drum.next_note2[25] ),
    .SET_B(net68),
    .Q(\disp_song.note2[25] ));
 sky130_fd_sc_hd__dfrtp_1 _6146_ (.CLK(clknet_leaf_26_clk),
    .D(net149),
    .RESET_B(net68),
    .Q(\disp_song.note2[26] ));
 sky130_fd_sc_hd__dfstp_1 _6147_ (.CLK(clknet_leaf_26_clk),
    .D(\disp_song.um.drum.next_note2[27] ),
    .SET_B(net68),
    .Q(\disp_song.note2[27] ));
 sky130_fd_sc_hd__dfrtp_1 _6148_ (.CLK(clknet_leaf_27_clk),
    .D(\disp_song.um.drum.next_note2[28] ),
    .RESET_B(net68),
    .Q(\disp_song.note2[28] ));
 sky130_fd_sc_hd__dfstp_1 _6149_ (.CLK(clknet_leaf_28_clk),
    .D(\disp_song.um.drum.next_note2[29] ),
    .SET_B(net68),
    .Q(\disp_song.note2[29] ));
 sky130_fd_sc_hd__dfrtp_1 _6150_ (.CLK(clknet_leaf_32_clk),
    .D(\disp_song.um.drum.next_note2[30] ),
    .RESET_B(net70),
    .Q(\disp_song.note2[30] ));
 sky130_fd_sc_hd__dfstp_1 _6151_ (.CLK(clknet_leaf_29_clk),
    .D(\disp_song.um.drum.next_note2[31] ),
    .SET_B(net69),
    .Q(\disp_song.note2[31] ));
 sky130_fd_sc_hd__dfrtp_1 _6152_ (.CLK(clknet_leaf_31_clk),
    .D(net1),
    .RESET_B(net70),
    .Q(\disp_song.um.boton0e.sync_b ));
 sky130_fd_sc_hd__dfrtp_1 _6153_ (.CLK(clknet_leaf_26_clk),
    .D(net83),
    .RESET_B(net70),
    .Q(\disp_song.um.boton0e.edge_2 ));
 sky130_fd_sc_hd__dfrtp_1 _6154_ (.CLK(clknet_leaf_31_clk),
    .D(net79),
    .RESET_B(net70),
    .Q(\disp_song.um.boton0e.edge_1 ));
 sky130_fd_sc_hd__dfrtp_1 _6155_ (.CLK(clknet_leaf_13_clk),
    .D(net2),
    .RESET_B(net58),
    .Q(\disp_song.um.boton1e.sync_b ));
 sky130_fd_sc_hd__dfrtp_1 _6156_ (.CLK(clknet_3_5__leaf_clk),
    .D(\disp_song.um.boton1e.edge_1 ),
    .RESET_B(net63),
    .Q(\disp_song.um.boton1e.edge_2 ));
 sky130_fd_sc_hd__dfrtp_2 _6157_ (.CLK(clknet_leaf_13_clk),
    .D(net76),
    .RESET_B(net58),
    .Q(\disp_song.um.boton1e.edge_1 ));
 sky130_fd_sc_hd__dfrtp_1 _6158_ (.CLK(clknet_leaf_30_clk),
    .D(net4),
    .RESET_B(net70),
    .Q(\disp_song.um.boton2e.sync_b ));
 sky130_fd_sc_hd__dfrtp_1 _6159_ (.CLK(clknet_leaf_31_clk),
    .D(net78),
    .RESET_B(net70),
    .Q(\disp_song.um.boton2e.edge_2 ));
 sky130_fd_sc_hd__dfrtp_1 _6160_ (.CLK(clknet_leaf_30_clk),
    .D(net74),
    .RESET_B(net70),
    .Q(\disp_song.um.boton2e.edge_1 ));
 sky130_fd_sc_hd__dfrtp_1 _6161_ (.CLK(clknet_leaf_8_clk),
    .D(\disp_song.um.drum.next_d2[0] ),
    .RESET_B(net60),
    .Q(\disp_song.display_note2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6162_ (.CLK(clknet_leaf_8_clk),
    .D(\disp_song.um.drum.next_d2[1] ),
    .RESET_B(net60),
    .Q(\disp_song.display_note2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6163_ (.CLK(clknet_leaf_21_clk),
    .D(\disp_song.um.drum.next_d2[2] ),
    .RESET_B(net61),
    .Q(\disp_song.display_note2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6164_ (.CLK(clknet_leaf_22_clk),
    .D(\disp_song.um.drum.next_d2[3] ),
    .RESET_B(net61),
    .Q(\disp_song.display_note2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6165_ (.CLK(clknet_leaf_8_clk),
    .D(\disp_song.um.drum.next_d2[4] ),
    .RESET_B(net61),
    .Q(\disp_song.display_note2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6166_ (.CLK(clknet_leaf_22_clk),
    .D(\disp_song.um.drum.next_d2[5] ),
    .RESET_B(net61),
    .Q(\disp_song.display_note2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6167_ (.CLK(clknet_leaf_5_clk),
    .D(\disp_song.um.drum.next_d2[6] ),
    .RESET_B(net60),
    .Q(\disp_song.display_note2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6168_ (.CLK(clknet_leaf_44_clk),
    .D(\disp_song.um.drum.next_d1[0] ),
    .RESET_B(net54),
    .Q(\disp_song.display_note1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6169_ (.CLK(clknet_leaf_45_clk),
    .D(\disp_song.um.drum.next_d1[1] ),
    .RESET_B(net54),
    .Q(\disp_song.display_note1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6170_ (.CLK(clknet_leaf_44_clk),
    .D(\disp_song.um.drum.next_d1[2] ),
    .RESET_B(net65),
    .Q(\disp_song.display_note1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6171_ (.CLK(clknet_leaf_43_clk),
    .D(\disp_song.um.drum.next_d1[3] ),
    .RESET_B(net65),
    .Q(\disp_song.display_note1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6172_ (.CLK(clknet_leaf_43_clk),
    .D(\disp_song.um.drum.next_d1[4] ),
    .RESET_B(net65),
    .Q(\disp_song.display_note1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6173_ (.CLK(clknet_leaf_45_clk),
    .D(\disp_song.um.drum.next_d1[5] ),
    .RESET_B(net54),
    .Q(\disp_song.display_note1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6174_ (.CLK(clknet_leaf_45_clk),
    .D(\disp_song.um.drum.next_d1[6] ),
    .RESET_B(net54),
    .Q(\disp_song.display_note1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6175_ (.CLK(clknet_leaf_24_clk),
    .D(\disp_song.next_red ),
    .RESET_B(net65),
    .Q(\disp_song.toggle_red ));
 sky130_fd_sc_hd__dfrtp_1 _6176_ (.CLK(clknet_leaf_44_clk),
    .D(\disp_song.next_green ),
    .RESET_B(net54),
    .Q(\disp_song.toggle_green ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__buf_8 fanout46 (.A(net73),
    .X(net46));
 sky130_fd_sc_hd__buf_4 fanout47 (.A(net73),
    .X(net47));
 sky130_fd_sc_hd__buf_8 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__buf_8 fanout49 (.A(net73),
    .X(net49));
 sky130_fd_sc_hd__buf_8 fanout50 (.A(net52),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_8 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__buf_8 fanout52 (.A(net73),
    .X(net52));
 sky130_fd_sc_hd__buf_8 fanout53 (.A(net73),
    .X(net53));
 sky130_fd_sc_hd__buf_4 fanout54 (.A(net73),
    .X(net54));
 sky130_fd_sc_hd__buf_6 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__buf_6 fanout56 (.A(net73),
    .X(net56));
 sky130_fd_sc_hd__buf_6 fanout57 (.A(net61),
    .X(net57));
 sky130_fd_sc_hd__buf_6 fanout58 (.A(net61),
    .X(net58));
 sky130_fd_sc_hd__buf_6 fanout59 (.A(net60),
    .X(net59));
 sky130_fd_sc_hd__buf_8 fanout60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_8 fanout61 (.A(net73),
    .X(net61));
 sky130_fd_sc_hd__buf_6 fanout62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__buf_8 fanout63 (.A(net73),
    .X(net63));
 sky130_fd_sc_hd__buf_6 fanout64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__buf_6 fanout65 (.A(net73),
    .X(net65));
 sky130_fd_sc_hd__buf_6 fanout66 (.A(net73),
    .X(net66));
 sky130_fd_sc_hd__buf_4 fanout67 (.A(net73),
    .X(net67));
 sky130_fd_sc_hd__buf_6 fanout68 (.A(net70),
    .X(net68));
 sky130_fd_sc_hd__buf_8 fanout69 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_8 fanout70 (.A(net73),
    .X(net70));
 sky130_fd_sc_hd__buf_6 fanout71 (.A(net73),
    .X(net71));
 sky130_fd_sc_hd__buf_4 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__buf_12 fanout73 (.A(net6),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\disp_song.um.boton2e.sync_b ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\disp_song.um.boton0e.edge_1 ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\game.scoring_button_2.flash_counter_1[13] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\game.scoring_button_2.flash_counter_1[16] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\game.flash_counter[21] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\game.scoring_button_2.flash_counter_1[4] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\game.scoring_button_1.flash_counter_2[4] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\game.addhits.add1.b[3] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\pulseout.fin_pulse[0] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\game.scoring_button_1.flash_counter_1[16] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\game.scoring_button_1.flash_counter_2[19] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\game.addhits.add4.b[0] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\game.scoring_button_2.check_hit.edge_1 ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\disp_song.note1[12] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\game.scoring_button_1.flash_counter_2[13] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\game.scoring_button_2.flash_counter_2[16] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\game.scoring_button_2.next_flash_counter_2[16] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\game.flash_counter[8] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\game.addhits.add2.b[0] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\game.addhits.a[12] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\game.addhits.add4.b[1] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\disp_song.note2[22] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\game.scoring_button_2.flash_counter_1[7] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\game.scoring_button_1.flash_counter_1[22] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\game.scoring_button_2.next_flash_counter_1[7] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\game.scoring_button_1.flash_counter_2[16] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\game.scoring_button_1.next_flash_counter_2[16] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\game.addhits.a[10] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\disp_song.note1[30] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\game.addhits.add3.b[2] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\game.counter[2] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\disp_song.note2[30] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\game.scoring_button_2.flash_counter_2[4] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\game.addhits.a[3] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\game.scoring_button_1.flash_counter_2[22] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\game.scoring_button_1.acc[1] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\disp_song.note1[23] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\disp_song.note1[22] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\game.addhits.a[14] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\game.scoring_button_1.flash_counter_1[4] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\game.addhits.a[2] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\game.padded_notes2[8] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\game.padded_notes1[24] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\game.padded_notes2[22] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\game.padded_notes1[28] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\game.scoring_button_2.flash_counter_2[22] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\game.addhits.add4.b[2] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\game.padded_notes1[9] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\game.addhits.a[13] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\game.addhits.a[8] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\game.padded_notes1[25] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\game.padded_notes1[4] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\game.addhits.add3.b[3] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\game.addhits.a[7] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\game.padded_notes2[24] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\game.padded_notes1[20] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\game.scoring_button_2.next_flash_counter_2[22] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\game.padded_notes1[29] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\game.padded_notes1[8] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\game.padded_notes1[21] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\game.padded_notes1[16] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\game.padded_notes2[6] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\game.addhits.a[11] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\game.padded_notes2[10] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\game.padded_notes2[18] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\game.padded_notes2[14] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\game.padded_notes1[1] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\game.scoring_button_2.flash_counter_1[22] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\game.padded_notes2[28] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\game.padded_notes2[30] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\game.padded_notes2[12] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\disp_song.note2[23] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\disp_song.note1[15] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\game.padded_notes1[17] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\game.padded_notes2[26] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\disp_song.note1[18] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\game.padded_notes1[12] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\game.padded_notes2[2] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\game.scoring_button_2.check_hit.in ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\game.padded_notes1[13] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\disp_song.note2[29] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\disp_song.note1[21] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\disp_song.note1[13] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\disp_song.note1[8] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\game.addmisses.a[12] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\game.addhits.add3.b[0] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\disp_song.note1[14] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\game.padded_notes2[20] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\game.scoring_button_2.acc[1] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\game.padded_notes2[0] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\game.addhits.add2.b[2] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\game.padded_notes2[4] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\disp_song.note2[31] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\game.padded_notes1[5] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\game.addhits.a[6] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\game.addhits.add3.b[1] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\disp_song.note1[24] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\game.addhits.a[9] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\game.padded_notes2[16] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\disp_song.note1[6] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0050_),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\game.flash_counter[18] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_2635_),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\pulseout.fin_pulse[5] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\disp_song.um.idx_note2[2] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\game.addhits.a[4] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\disp_song.note1[7] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\game.out[12] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\modetrans.mode[4] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\modetrans.u2.sync_pb ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\game.out[6] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0128_),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\game.scoring_button_1.check_hit.in ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\game.flash_counter[4] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\disp_song.note1[0] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_0090_),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\game.flash_counter[1] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_2596_),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\game.out[2] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_0125_),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\disp_song.um.boton1e.sync_b ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\game.scoring_button_2.flash_counter_1[1] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\game.scoring_button_2.next_flash_counter_1[1] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\game.scoring_button_1.flash_counter_2[1] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\game.scoring_button_1.next_flash_counter_2[1] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\game.scoring_button_2.flash_counter_2[1] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\game.scoring_button_2.next_flash_counter_2[1] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\game.counter[0] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\game.out[13] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\game.scoring_button_1.flash_counter_1[1] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\game.scoring_button_1.next_flash_counter_1[1] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\modetrans.u3.sync_pb ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\game.flash_counter[2] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\modetrans.u2.Q2 ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\game.out[4] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_0126_),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\game.out[11] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_0086_),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\game.out[1] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_0123_),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\game.flash_counter[14] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\disp_song.note1[28] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\disp_song.um.boton2e.edge_1 ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\game.beat_clk ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\game.flash_counter[0] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\game.flash_counter[22] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\game.flash_counter[11] ),
    .X(net126));
 sky130_fd_sc_hd__buf_1 hold54 (.A(\game.out[5] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\pulseout.fin_pulse[2] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\game.flash_counter[9] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_0138_),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\game.scoring_button_2.hit ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0049_),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\disp_song.um.boton0e.sync_b ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\game.out[7] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_0082_),
    .X(net134));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold62 (.A(\game.out[12] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0087_),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\game.flash_counter[17] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\game.out[0] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0122_),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\game.out[9] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0084_),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\game.flash_counter[6] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\modetrans.u3.Q1 ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\game.out[8] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\game.counter[12] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\game.out[10] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\game.flash_counter[5] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\pulseout.fin_pulse[4] ),
    .X(net147));
 sky130_fd_sc_hd__buf_1 hold75 (.A(\disp_song.um.boton1e.edge_2 ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\disp_song.um.drum.next_note2[26] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\disp_song.note1[25] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\game.scoring_button_2.flash_counter_2[7] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\highest_score.highest_score[7] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\game.scoring_button_1.check_hit.edge_1 ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\game.addhits.add2.b[3] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\disp_song.note1[26] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\game.scoring_button_1.flash_counter_1[13] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\game.scoring_button_2.flash_counter_1[10] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\game.scoring_button_1.flash_counter_1[10] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\game.scoring_button_1.flash_counter_2[10] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\game.scoring_button_2.flash_counter_2[13] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\disp_song.note1[31] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\game.scoring_button_1.flash_counter_2[7] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\game.scoring_button_1.flash_counter_1[7] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\modetrans.u2.Q1 ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\disp_song.note1[20] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\modetrans.mode[4] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\disp_song.note1[29] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\game.scoring_button_2.flash_counter_2[10] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\game.addhits.add1.b[2] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\game.counter[4] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\game.scoring_button_2.flash_counter_2[19] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\game.scoring_button_1.hit ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\game.scoring_button_2.flash_counter_1[19] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\game.scoring_button_1.flash_counter_1[19] ),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(button[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(button[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(button[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(button[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(chip_select),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(n_rst),
    .X(net6));
 sky130_fd_sc_hd__buf_1 max_cap37 (.A(_2610_),
    .X(net37));
 sky130_fd_sc_hd__buf_2 max_cap42 (.A(_0842_),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 max_cap43 (.A(_0811_),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 max_cap44 (.A(_0885_),
    .X(net44));
 sky130_fd_sc_hd__buf_2 max_cap45 (.A(_1313_),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 output10 (.A(net10),
    .X(bottom_row[3]));
 sky130_fd_sc_hd__clkbuf_4 output11 (.A(net11),
    .X(bottom_row[4]));
 sky130_fd_sc_hd__clkbuf_4 output12 (.A(net12),
    .X(bottom_row[5]));
 sky130_fd_sc_hd__clkbuf_4 output13 (.A(net13),
    .X(bottom_row[6]));
 sky130_fd_sc_hd__clkbuf_4 output14 (.A(net14),
    .X(green_disp));
 sky130_fd_sc_hd__clkbuf_4 output15 (.A(net15),
    .X(red_disp));
 sky130_fd_sc_hd__clkbuf_4 output16 (.A(net16),
    .X(ss0[0]));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(ss0[1]));
 sky130_fd_sc_hd__clkbuf_4 output18 (.A(net18),
    .X(ss0[2]));
 sky130_fd_sc_hd__clkbuf_4 output19 (.A(net19),
    .X(ss0[3]));
 sky130_fd_sc_hd__clkbuf_4 output20 (.A(net20),
    .X(ss0[4]));
 sky130_fd_sc_hd__clkbuf_4 output21 (.A(net21),
    .X(ss0[5]));
 sky130_fd_sc_hd__clkbuf_4 output22 (.A(net22),
    .X(ss0[6]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(ss1[0]));
 sky130_fd_sc_hd__clkbuf_4 output24 (.A(net24),
    .X(ss1[1]));
 sky130_fd_sc_hd__clkbuf_4 output25 (.A(net25),
    .X(ss1[2]));
 sky130_fd_sc_hd__clkbuf_4 output26 (.A(net26),
    .X(ss1[3]));
 sky130_fd_sc_hd__clkbuf_4 output27 (.A(net27),
    .X(ss1[4]));
 sky130_fd_sc_hd__clkbuf_4 output28 (.A(net28),
    .X(ss1[5]));
 sky130_fd_sc_hd__clkbuf_4 output29 (.A(net29),
    .X(ss1[6]));
 sky130_fd_sc_hd__clkbuf_4 output30 (.A(net30),
    .X(top_row[0]));
 sky130_fd_sc_hd__clkbuf_4 output31 (.A(net31),
    .X(top_row[1]));
 sky130_fd_sc_hd__clkbuf_4 output32 (.A(net32),
    .X(top_row[2]));
 sky130_fd_sc_hd__clkbuf_4 output33 (.A(net33),
    .X(top_row[3]));
 sky130_fd_sc_hd__clkbuf_4 output34 (.A(net34),
    .X(top_row[4]));
 sky130_fd_sc_hd__clkbuf_4 output35 (.A(net35),
    .X(top_row[5]));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net36),
    .X(top_row[6]));
 sky130_fd_sc_hd__clkbuf_4 output7 (.A(net7),
    .X(bottom_row[0]));
 sky130_fd_sc_hd__clkbuf_4 output8 (.A(net8),
    .X(bottom_row[1]));
 sky130_fd_sc_hd__clkbuf_4 output9 (.A(net9),
    .X(bottom_row[2]));
 sky130_fd_sc_hd__buf_2 wire38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__buf_2 wire39 (.A(_0878_),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 wire40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 wire41 (.A(_0852_),
    .X(net41));
endmodule

